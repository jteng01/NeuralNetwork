module mlp_neural_net #(
    parameter int INPUTS           = 784,
    parameter int OUTPUTS          = 10,
    parameter int OUTPUT_IDX_BITS  = 4
) (
    input  logic signed [31:0] data_inputs  [0:INPUTS-1],
    output logic signed [31:0] data_outputs [0:OUTPUTS-1],
    output logic [OUTPUT_IDX_BITS-1:0] predicted_class
);


    //Layer 0: 784 inputs, 128 neurons
    localparam logic signed [31:0] layer0_weights [0:127][0:783] = '{
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd750501, 32'sd1197721, 32'sd1313312, 32'sd1514653, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd327160, 32'sd447521, 32'sd2020916, 32'sd662856, 32'sd1248200, 32'sd2063605, 32'sd1863258, 32'sd2600131, 32'sd728646, 32'sd141799, 32'sd279471, 32'sd461735, 32'sd1379954, 32'sd14443, 32'sd873770, -32'sd542380, -32'sd160523, -32'sd11474, 32'sd602004, 32'sd593453, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1114274, 32'sd464871, -32'sd638918, -32'sd800600, 32'sd1672851, 32'sd206363, 32'sd655611, -32'sd748958, 32'sd1974611, 32'sd869311, -32'sd927711, -32'sd41482, 32'sd367647, 32'sd1346340, 32'sd1195030, 32'sd2897798, 32'sd3591810, 32'sd2994325, 32'sd380459, 32'sd1830042, 32'sd623538, 32'sd766499, 32'sd1584409, 32'sd500890, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1445449, 32'sd104232, 32'sd85107, 32'sd612265, -32'sd663523, 32'sd225410, -32'sd470220, -32'sd514560, 32'sd1022063, 32'sd1173082, 32'sd284125, -32'sd773759, -32'sd277231, -32'sd1225094, -32'sd583147, 32'sd1495672, 32'sd561007, -32'sd2101128, 32'sd1494208, 32'sd911829, 32'sd129107, 32'sd557933, 32'sd1548751, 32'sd133, 32'sd488338, 32'sd0, 32'sd0, 32'sd116655, 32'sd542403, -32'sd290347, -32'sd970661, 32'sd1517160, -32'sd2012514, -32'sd1972628, -32'sd1291879, -32'sd2872801, -32'sd775804, -32'sd981948, -32'sd3540352, -32'sd2275671, -32'sd2244788, 32'sd1375305, -32'sd1296127, 32'sd761854, 32'sd1621725, 32'sd1885679, 32'sd1415387, 32'sd880337, 32'sd17632, 32'sd1406190, -32'sd252221, 32'sd1161032, 32'sd216401, 32'sd1324920, 32'sd0, 32'sd748047, 32'sd141222, -32'sd822591, -32'sd1287441, -32'sd1286653, -32'sd407551, -32'sd2426067, -32'sd1601477, -32'sd1792220, -32'sd800604, -32'sd1216377, -32'sd3815991, -32'sd754782, -32'sd1011685, 32'sd260978, -32'sd1746137, 32'sd609138, -32'sd1363494, 32'sd1097256, 32'sd2389714, 32'sd137041, 32'sd675737, 32'sd10635, 32'sd304894, -32'sd731224, -32'sd1278338, 32'sd189605, 32'sd0, 32'sd694681, -32'sd994063, -32'sd53748, -32'sd626244, 32'sd1137062, -32'sd371150, -32'sd211593, -32'sd2926264, -32'sd2681455, -32'sd1616643, -32'sd2470746, 32'sd1412260, -32'sd185080, -32'sd114577, 32'sd407001, -32'sd2831964, -32'sd659921, 32'sd288612, 32'sd2090602, 32'sd2069310, 32'sd392891, 32'sd1692138, -32'sd1629244, 32'sd1056305, 32'sd91207, 32'sd589519, -32'sd68154, 32'sd405775, -32'sd40991, -32'sd687738, 32'sd552025, -32'sd206106, -32'sd712521, -32'sd1550693, -32'sd557517, -32'sd2213003, -32'sd1576974, -32'sd645147, 32'sd622355, 32'sd95659, 32'sd2580402, -32'sd713698, -32'sd2414923, 32'sd30794, 32'sd457126, 32'sd2995867, 32'sd1831785, 32'sd572459, 32'sd971947, 32'sd3407158, 32'sd1470599, 32'sd869260, -32'sd14142, -32'sd657197, -32'sd57611, 32'sd398417, 32'sd767951, 32'sd152939, -32'sd118149, 32'sd1167721, 32'sd171300, -32'sd423135, -32'sd603177, -32'sd1530403, -32'sd942498, -32'sd2430463, -32'sd1368946, 32'sd3105176, 32'sd1934607, 32'sd1215670, 32'sd616014, 32'sd1844159, 32'sd642590, 32'sd1576588, -32'sd37603, 32'sd2449376, 32'sd546751, 32'sd2181592, 32'sd1973215, 32'sd2983549, 32'sd1894133, 32'sd404434, 32'sd961618, 32'sd522172, 32'sd771781, 32'sd1444620, 32'sd215638, 32'sd1887952, 32'sd1500660, 32'sd1367518, -32'sd798863, -32'sd2251011, -32'sd2819696, -32'sd267227, 32'sd1199743, 32'sd2639814, 32'sd1383041, 32'sd3378062, 32'sd1592967, -32'sd144414, 32'sd241447, 32'sd1292105, 32'sd373116, 32'sd1806178, -32'sd42, -32'sd185911, 32'sd965149, 32'sd1873998, 32'sd1197734, 32'sd25537, -32'sd1321076, -32'sd1049424, -32'sd492294, -32'sd179495, -32'sd295296, 32'sd778234, 32'sd2514416, 32'sd1132635, -32'sd1740719, -32'sd1398104, 32'sd201833, 32'sd193710, 32'sd362787, 32'sd1089431, 32'sd2267897, 32'sd2093207, 32'sd1484096, -32'sd69612, -32'sd334494, -32'sd345240, -32'sd423183, 32'sd1004770, 32'sd1190641, 32'sd1626264, 32'sd928745, -32'sd884781, 32'sd626282, 32'sd1195436, 32'sd647821, 32'sd680851, -32'sd941803, -32'sd1627092, -32'sd1184436, 32'sd2697739, -32'sd714928, 32'sd1477215, 32'sd1724358, 32'sd2560467, -32'sd96719, -32'sd984286, 32'sd2223008, 32'sd1610315, 32'sd913806, 32'sd62293, -32'sd1028350, -32'sd2871288, -32'sd4071654, -32'sd2408635, -32'sd1005948, 32'sd3799, -32'sd2655057, -32'sd2736131, -32'sd1314971, -32'sd764775, -32'sd1231535, -32'sd246881, -32'sd320048, 32'sd15549, -32'sd951328, -32'sd532004, 32'sd1496464, 32'sd619512, 32'sd22333, 32'sd666528, 32'sd1614714, 32'sd2105247, 32'sd1475934, -32'sd1364525, 32'sd978164, 32'sd194500, 32'sd854319, -32'sd1576816, -32'sd1538614, -32'sd4508727, -32'sd5244016, -32'sd2650904, -32'sd1396339, -32'sd1494691, -32'sd1170588, -32'sd1624400, -32'sd1465390, 32'sd1341547, 32'sd889876, -32'sd1584121, 32'sd199865, 32'sd138404, 32'sd195042, -32'sd167010, 32'sd347012, -32'sd1299003, 32'sd173678, 32'sd1793342, 32'sd1646246, -32'sd1479242, -32'sd359534, 32'sd639697, -32'sd705395, 32'sd1103099, -32'sd971862, -32'sd249516, -32'sd414294, -32'sd3933440, -32'sd2228809, -32'sd1357401, -32'sd2160607, -32'sd2786434, -32'sd2380059, 32'sd1376233, 32'sd1497695, 32'sd459315, -32'sd560121, -32'sd1922662, 32'sd1349320, -32'sd351033, 32'sd674469, 32'sd771684, -32'sd514507, 32'sd17448, 32'sd495135, -32'sd1239591, 32'sd458089, -32'sd1816370, -32'sd391650, 32'sd898703, -32'sd975406, -32'sd323856, -32'sd2840785, -32'sd2507312, -32'sd1074244, -32'sd3565506, 32'sd1467263, -32'sd729572, 32'sd213670, 32'sd12885, 32'sd659160, 32'sd491326, 32'sd1078025, -32'sd595316, -32'sd716347, -32'sd363215, 32'sd1153919, -32'sd308287, -32'sd1172802, -32'sd1066424, -32'sd617386, 32'sd1178969, 32'sd1086535, -32'sd1593363, 32'sd598471, -32'sd634440, -32'sd886189, -32'sd845309, 32'sd142688, 32'sd601357, 32'sd372383, -32'sd914116, -32'sd390766, -32'sd1091699, 32'sd3690851, 32'sd2164450, -32'sd192960, -32'sd1618219, 32'sd1822789, 32'sd111349, 32'sd776903, 32'sd1878566, -32'sd474411, 32'sd1992443, 32'sd416676, 32'sd451824, -32'sd201552, -32'sd993049, -32'sd1258705, -32'sd261162, -32'sd238611, -32'sd508228, 32'sd1291296, 32'sd1833760, 32'sd1099156, -32'sd344854, -32'sd94395, 32'sd3166213, -32'sd940624, 32'sd1514768, -32'sd218942, 32'sd186692, 32'sd2487615, 32'sd1905466, -32'sd68856, -32'sd3639890, 32'sd585650, 32'sd522882, 32'sd142129, 32'sd1535913, 32'sd1752801, 32'sd1452390, 32'sd1096738, 32'sd0, -32'sd276553, 32'sd701802, 32'sd558978, -32'sd1001839, -32'sd1077302, -32'sd82692, 32'sd1402581, 32'sd1409030, 32'sd987904, 32'sd196714, -32'sd648860, -32'sd1342960, -32'sd1689515, 32'sd243079, 32'sd2734051, 32'sd828203, 32'sd1094898, 32'sd107426, -32'sd747040, -32'sd1636786, -32'sd55691, 32'sd1476693, 32'sd2344878, 32'sd974644, 32'sd404567, 32'sd518709, -32'sd160762, 32'sd886247, 32'sd414513, 32'sd644028, 32'sd1237305, -32'sd979303, 32'sd875663, 32'sd715367, 32'sd3105706, 32'sd2035297, -32'sd754600, -32'sd1778072, -32'sd3679298, -32'sd995882, -32'sd2725193, 32'sd441585, 32'sd1658770, 32'sd3588867, 32'sd1117306, 32'sd432325, -32'sd2101709, -32'sd2282476, -32'sd1681173, 32'sd383623, 32'sd1116986, -32'sd139756, -32'sd1539001, -32'sd234845, 32'sd153553, 32'sd61239, 32'sd249421, 32'sd1860808, -32'sd1296572, -32'sd1012916, 32'sd691179, 32'sd1992474, 32'sd906552, 32'sd1787234, -32'sd1090235, -32'sd1661259, -32'sd1589316, 32'sd312170, -32'sd412506, -32'sd475338, 32'sd2068051, 32'sd2182756, -32'sd529969, -32'sd721578, -32'sd3950100, -32'sd2372879, -32'sd602473, 32'sd2839177, 32'sd686267, -32'sd628877, -32'sd1701956, -32'sd1488545, -32'sd569220, 32'sd0, 32'sd148430, 32'sd952323, 32'sd109162, -32'sd430183, 32'sd1675616, 32'sd1997134, 32'sd1660997, 32'sd3087988, 32'sd1001383, 32'sd1514680, 32'sd1506309, 32'sd1419701, 32'sd1311518, -32'sd1730534, -32'sd199742, -32'sd1053690, -32'sd1144272, -32'sd1318429, -32'sd767801, -32'sd2150322, -32'sd877411, 32'sd1191164, -32'sd446877, -32'sd120812, -32'sd2159048, -32'sd1032320, 32'sd501293, -32'sd183302, 32'sd192026, 32'sd245930, 32'sd1391998, 32'sd1704377, 32'sd317492, -32'sd358547, 32'sd1291820, 32'sd103879, 32'sd1147430, 32'sd346927, 32'sd79882, 32'sd1512659, 32'sd2251792, -32'sd1019651, -32'sd836293, -32'sd834961, 32'sd967648, -32'sd3302057, -32'sd1120834, -32'sd1297972, -32'sd1301868, 32'sd155468, -32'sd896962, -32'sd2193450, -32'sd107796, -32'sd762622, 32'sd838688, 32'sd624097, 32'sd63587, 32'sd138257, 32'sd2071451, -32'sd200899, -32'sd1267976, 32'sd1814681, 32'sd89182, -32'sd679525, -32'sd560469, 32'sd2484124, -32'sd125135, 32'sd892089, 32'sd788309, 32'sd185911, -32'sd760726, 32'sd14961, 32'sd1315275, -32'sd1227719, 32'sd11282, 32'sd217290, -32'sd949965, 32'sd1810871, 32'sd772707, -32'sd1392752, -32'sd1655042, -32'sd345200, 32'sd732819, 32'sd0, 32'sd759274, -32'sd74100, 32'sd62008, 32'sd1609379, -32'sd1164283, 32'sd3310385, 32'sd2724872, 32'sd1804158, 32'sd380016, 32'sd739972, 32'sd932461, 32'sd2224956, 32'sd1422139, 32'sd995339, -32'sd624971, -32'sd1166895, -32'sd2562867, -32'sd1365333, -32'sd1522493, 32'sd728153, -32'sd184754, 32'sd1604235, -32'sd114287, -32'sd1974609, 32'sd713062, -32'sd1271215, 32'sd0, 32'sd0, 32'sd0, 32'sd385012, -32'sd912528, -32'sd209121, 32'sd201746, 32'sd1016748, 32'sd2650096, 32'sd672999, -32'sd310843, 32'sd57635, 32'sd1151036, 32'sd235338, -32'sd798981, -32'sd2194605, 32'sd252296, 32'sd1115157, 32'sd963477, -32'sd506077, 32'sd1235027, -32'sd256707, -32'sd730260, -32'sd1648992, 32'sd1074742, -32'sd2231471, 32'sd195469, 32'sd52370, 32'sd0, 32'sd0, 32'sd0, 32'sd268502, 32'sd309935, 32'sd24130, -32'sd398572, -32'sd213580, -32'sd66223, -32'sd2697746, 32'sd1252737, 32'sd2021522, 32'sd2745619, 32'sd851293, 32'sd167586, -32'sd1370325, 32'sd521029, 32'sd362088, 32'sd2124582, 32'sd1679947, 32'sd2785333, 32'sd2155552, 32'sd1597994, 32'sd27496, 32'sd543262, 32'sd256088, 32'sd138476, 32'sd45050, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1143509, -32'sd917694, 32'sd36539, -32'sd2031677, 32'sd994089, -32'sd1135248, 32'sd324550, -32'sd10678, 32'sd2376021, 32'sd3578327, 32'sd2436787, -32'sd835124, 32'sd1664498, -32'sd91864, -32'sd2030333, -32'sd1054676, -32'sd2052450, -32'sd618787, 32'sd550392, -32'sd471966, 32'sd996536, 32'sd120175, 32'sd539354, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1460230, 32'sd1233075, 32'sd286822, -32'sd229457, 32'sd196255, 32'sd1505214, -32'sd948458, 32'sd1224689, 32'sd2028054, 32'sd475991, 32'sd2127859, -32'sd256640, -32'sd1234094, -32'sd663089, 32'sd724357, -32'sd47733, 32'sd1245092, 32'sd307126, -32'sd789690, 32'sd318434, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd740667, 32'sd362289, 32'sd1002445, 32'sd1056804, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd192193, -32'sd647478, -32'sd705342, -32'sd960735, -32'sd1013810, 32'sd223338, 32'sd639129, 32'sd28830, -32'sd160741, -32'sd119570, 32'sd41559, -32'sd342744, -32'sd1150450, -32'sd2027071, -32'sd582260, 32'sd657052, 32'sd142577, -32'sd711022, -32'sd1028060, -32'sd1064479, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd143240, -32'sd792910, -32'sd1456331, 32'sd837349, -32'sd1014685, -32'sd51920, -32'sd652918, 32'sd1190347, 32'sd1444654, 32'sd1430745, 32'sd486145, 32'sd323558, 32'sd1043034, -32'sd1328082, -32'sd1178064, -32'sd616393, 32'sd246168, -32'sd3082959, -32'sd1894646, -32'sd1622722, -32'sd821889, -32'sd169514, -32'sd321798, -32'sd30169, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd158984, -32'sd1403471, -32'sd844945, -32'sd145670, 32'sd365099, -32'sd7589, 32'sd1646557, 32'sd1427512, 32'sd390152, -32'sd404158, -32'sd323004, 32'sd624990, -32'sd106564, 32'sd871072, -32'sd839245, -32'sd1413947, 32'sd1879433, 32'sd1159136, -32'sd340618, -32'sd1298433, 32'sd481886, 32'sd623522, 32'sd794648, -32'sd96201, 32'sd190192, 32'sd0, 32'sd0, -32'sd666480, -32'sd1239218, -32'sd746517, 32'sd676457, -32'sd821969, -32'sd761343, -32'sd673903, -32'sd911425, 32'sd388167, 32'sd167975, 32'sd828118, 32'sd190775, -32'sd480148, 32'sd184643, 32'sd1461186, 32'sd679764, 32'sd973891, 32'sd1720416, 32'sd1723453, 32'sd498367, -32'sd1151563, 32'sd565895, 32'sd525966, -32'sd578521, 32'sd1461720, -32'sd447349, -32'sd41192, 32'sd0, -32'sd47098, -32'sd1698289, -32'sd20674, 32'sd88867, -32'sd1100453, -32'sd779389, -32'sd2824533, 32'sd288019, -32'sd151543, -32'sd769809, -32'sd639507, -32'sd1474359, 32'sd158483, -32'sd958628, 32'sd807878, 32'sd1664451, 32'sd579847, 32'sd1098227, 32'sd1459029, 32'sd2306567, 32'sd2367203, 32'sd329133, -32'sd509790, 32'sd46192, 32'sd533650, -32'sd37908, -32'sd328683, 32'sd0, 32'sd419455, -32'sd1957092, 32'sd482716, 32'sd807910, -32'sd624796, -32'sd239179, -32'sd471137, -32'sd2175464, -32'sd2878222, -32'sd1698076, -32'sd1347320, -32'sd1629136, -32'sd1091376, -32'sd888545, 32'sd2231576, 32'sd4299749, 32'sd2065062, 32'sd3146282, 32'sd491816, -32'sd95801, 32'sd834147, 32'sd397611, -32'sd283070, -32'sd2983481, 32'sd566692, 32'sd560971, 32'sd25191, -32'sd160626, 32'sd503083, -32'sd1283412, 32'sd428472, -32'sd166016, -32'sd2224566, -32'sd847847, -32'sd3288585, -32'sd1821958, -32'sd4713256, -32'sd4222816, -32'sd835334, 32'sd865644, 32'sd1546454, 32'sd807072, 32'sd2563792, 32'sd1194819, 32'sd2487712, -32'sd324957, -32'sd19736, -32'sd3095356, 32'sd970752, 32'sd1612073, 32'sd1008583, -32'sd2397969, -32'sd1636790, 32'sd690359, -32'sd685689, -32'sd1251847, -32'sd1915347, -32'sd515418, -32'sd108562, -32'sd162354, -32'sd403479, -32'sd1315218, -32'sd1676876, -32'sd2480223, -32'sd1865461, -32'sd445521, -32'sd308691, 32'sd689516, -32'sd186571, 32'sd616853, -32'sd899990, -32'sd184945, -32'sd1282094, 32'sd137208, 32'sd878968, -32'sd404574, -32'sd1844177, 32'sd867632, 32'sd986122, -32'sd1374439, 32'sd1041128, 32'sd1011726, 32'sd332615, -32'sd1430827, 32'sd1410059, -32'sd1878220, -32'sd2348750, -32'sd1494354, -32'sd3514034, -32'sd1315619, 32'sd840468, -32'sd242850, 32'sd477617, 32'sd1444463, 32'sd2106582, 32'sd705737, 32'sd44610, -32'sd1071879, -32'sd1182409, -32'sd2444020, -32'sd2432578, 32'sd1463946, 32'sd1429470, 32'sd2063611, 32'sd1425257, -32'sd571489, 32'sd165669, -32'sd1532379, 32'sd2269012, 32'sd15452, -32'sd1362434, -32'sd1093830, 32'sd809671, -32'sd75439, 32'sd551745, -32'sd563763, -32'sd798023, 32'sd1245183, -32'sd513458, 32'sd318569, 32'sd375582, 32'sd939360, 32'sd1899699, 32'sd48631, -32'sd1604610, -32'sd2758561, -32'sd2072499, -32'sd2268710, -32'sd2066647, 32'sd1449185, 32'sd758927, 32'sd1101504, -32'sd156580, 32'sd1662504, 32'sd1835133, 32'sd788511, -32'sd285402, -32'sd418912, 32'sd769171, -32'sd1373960, -32'sd1325304, 32'sd70800, -32'sd1050764, -32'sd410683, 32'sd1273740, 32'sd2598945, 32'sd3332839, -32'sd1550865, -32'sd937412, -32'sd684349, 32'sd536807, -32'sd3041571, -32'sd4505772, -32'sd2413525, -32'sd1069873, -32'sd688519, -32'sd2063633, 32'sd1446802, 32'sd2479965, -32'sd120198, 32'sd863627, 32'sd834140, 32'sd782765, -32'sd139360, 32'sd127779, 32'sd26909, -32'sd1618236, -32'sd1434059, -32'sd2039315, -32'sd1250661, 32'sd1341314, 32'sd2289050, 32'sd2028496, 32'sd3003831, 32'sd363154, -32'sd630256, -32'sd478666, -32'sd1732692, -32'sd3385884, -32'sd3681990, -32'sd2861949, 32'sd1832931, -32'sd929813, -32'sd768329, 32'sd395898, -32'sd601030, -32'sd394137, -32'sd1230999, 32'sd1824116, -32'sd110107, 32'sd2178624, 32'sd1514203, -32'sd458801, -32'sd1993815, 32'sd181909, -32'sd581898, -32'sd1967735, 32'sd49932, 32'sd2979814, 32'sd904644, -32'sd1717001, -32'sd95845, -32'sd1531476, -32'sd1019919, 32'sd466391, -32'sd2220229, -32'sd3369726, -32'sd4171615, -32'sd1183198, 32'sd2135749, -32'sd244483, -32'sd934747, -32'sd639212, -32'sd1159843, -32'sd1462153, -32'sd580686, -32'sd282304, 32'sd292828, 32'sd130508, -32'sd1021830, -32'sd2255240, -32'sd2220412, -32'sd1368582, -32'sd861023, -32'sd2262874, -32'sd440390, 32'sd972709, -32'sd2872910, -32'sd2194709, -32'sd2620075, -32'sd4570470, -32'sd4272107, -32'sd2816773, -32'sd2965186, -32'sd1781424, -32'sd630535, 32'sd370954, 32'sd2866153, 32'sd1862377, -32'sd60960, -32'sd2592468, -32'sd944390, -32'sd977109, -32'sd3833780, -32'sd1875832, -32'sd1365128, -32'sd1640280, -32'sd1543700, 32'sd259617, 32'sd1155754, -32'sd1082141, 32'sd167822, -32'sd224776, 32'sd291326, -32'sd1347879, -32'sd2231086, -32'sd3404208, -32'sd3090484, -32'sd1876091, -32'sd918712, -32'sd2087702, -32'sd711332, -32'sd624552, -32'sd852967, 32'sd1905264, 32'sd3328525, 32'sd100462, -32'sd879464, -32'sd1633950, -32'sd420439, -32'sd1108308, -32'sd2405594, -32'sd3519746, -32'sd514534, -32'sd1166132, -32'sd2234772, -32'sd1164719, -32'sd380308, 32'sd682893, 32'sd424430, -32'sd1046699, -32'sd1155331, 32'sd348907, -32'sd1275598, -32'sd2637525, -32'sd1803398, -32'sd189972, 32'sd571091, 32'sd1126751, 32'sd1264381, 32'sd1479331, 32'sd559916, 32'sd832276, 32'sd2617291, -32'sd1238258, -32'sd1454899, -32'sd2082346, -32'sd3137169, -32'sd2192178, -32'sd1186877, -32'sd509845, -32'sd787138, 32'sd514117, -32'sd230993, -32'sd1031193, -32'sd1815680, 32'sd162472, 32'sd0, -32'sd867482, -32'sd1636220, -32'sd137893, -32'sd240891, -32'sd378440, -32'sd438545, 32'sd1001450, 32'sd959965, 32'sd1677021, 32'sd2050157, 32'sd1791070, 32'sd1838227, -32'sd227298, -32'sd728629, 32'sd1499890, -32'sd980495, -32'sd776261, -32'sd2475831, -32'sd1373493, -32'sd1891332, -32'sd2589355, -32'sd538715, -32'sd1567368, -32'sd1463482, 32'sd784854, -32'sd456567, -32'sd206973, -32'sd585592, -32'sd1263714, -32'sd816810, -32'sd67799, 32'sd701841, 32'sd1555529, 32'sd1981072, 32'sd2894457, 32'sd637476, 32'sd66026, 32'sd617407, -32'sd969610, -32'sd1878768, -32'sd1913401, 32'sd1046026, 32'sd922291, 32'sd1674396, -32'sd169478, -32'sd1042787, -32'sd2544729, -32'sd754386, -32'sd996807, -32'sd1527813, -32'sd2578439, -32'sd812209, -32'sd117196, 32'sd880949, 32'sd795430, -32'sd740279, -32'sd1323484, -32'sd2464143, -32'sd2038528, 32'sd812877, 32'sd60587, 32'sd854466, 32'sd984722, 32'sd230530, 32'sd382210, -32'sd1865413, -32'sd2445455, -32'sd1115655, -32'sd1343767, 32'sd631431, 32'sd1686397, 32'sd1355989, 32'sd474769, 32'sd434509, -32'sd1125660, 32'sd1200942, 32'sd897531, -32'sd1199534, -32'sd555965, 32'sd1327860, -32'sd1148301, -32'sd159181, -32'sd1388630, 32'sd0, -32'sd1916800, -32'sd1691657, -32'sd208041, 32'sd117874, 32'sd1655108, 32'sd214735, 32'sd3377729, 32'sd3393804, 32'sd2617084, -32'sd691371, -32'sd2398969, 32'sd34036, -32'sd1529520, 32'sd484239, 32'sd1674270, 32'sd1171061, 32'sd3350437, 32'sd2784407, 32'sd406333, 32'sd1965687, 32'sd891765, -32'sd574210, 32'sd69935, -32'sd329125, 32'sd605394, 32'sd162315, -32'sd658295, 32'sd12608, -32'sd1284813, -32'sd1719668, -32'sd648306, 32'sd1418020, 32'sd1465566, 32'sd736510, 32'sd2340596, 32'sd2573556, -32'sd29639, -32'sd721575, -32'sd128658, -32'sd1236184, 32'sd1850692, 32'sd1736635, 32'sd2012709, 32'sd847772, 32'sd2218825, 32'sd2697994, 32'sd3513440, 32'sd27893, 32'sd786634, 32'sd172541, 32'sd306074, -32'sd126139, 32'sd229861, 32'sd15415, 32'sd263298, -32'sd26288, 32'sd32823, -32'sd298985, 32'sd1642285, 32'sd1998321, 32'sd171803, 32'sd2159317, 32'sd1226331, 32'sd147417, -32'sd17313, -32'sd145535, 32'sd1526293, 32'sd2540297, 32'sd1787347, 32'sd2203361, 32'sd102851, 32'sd577465, 32'sd1022913, 32'sd1204091, 32'sd1667839, 32'sd81950, 32'sd742054, 32'sd920297, 32'sd607828, 32'sd236091, 32'sd613065, -32'sd451443, 32'sd241488, 32'sd0, -32'sd907244, 32'sd335363, 32'sd165652, -32'sd197847, 32'sd956480, -32'sd12632, -32'sd501465, 32'sd361356, -32'sd484037, 32'sd2246128, 32'sd2902011, 32'sd1517249, 32'sd1449848, 32'sd94454, -32'sd893372, 32'sd2076666, -32'sd367500, 32'sd56857, -32'sd334497, -32'sd237160, 32'sd2312112, 32'sd1363969, 32'sd1342484, -32'sd280096, -32'sd1570753, -32'sd1639636, 32'sd0, 32'sd0, 32'sd0, -32'sd413535, 32'sd259568, 32'sd929069, -32'sd1681754, -32'sd860927, -32'sd1180565, -32'sd708294, -32'sd1541278, -32'sd275729, 32'sd1287150, -32'sd384488, -32'sd653211, -32'sd2493899, -32'sd23722, -32'sd1400746, 32'sd490367, 32'sd1109772, -32'sd656907, -32'sd388225, 32'sd684867, -32'sd1388592, 32'sd398459, -32'sd184313, -32'sd616708, -32'sd75276, 32'sd0, 32'sd0, 32'sd0, -32'sd1005724, 32'sd282194, -32'sd2108228, -32'sd1196752, -32'sd499416, -32'sd2044264, 32'sd233727, -32'sd1126078, -32'sd1584480, -32'sd708092, -32'sd2327121, 32'sd389681, 32'sd1012109, -32'sd866014, -32'sd988223, -32'sd1389416, -32'sd1712832, -32'sd2400147, 32'sd61542, -32'sd523272, -32'sd698126, -32'sd1691742, -32'sd1555716, 32'sd302116, -32'sd261038, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd210132, -32'sd405523, -32'sd1005958, -32'sd594044, -32'sd1251545, 32'sd978624, 32'sd992818, 32'sd433, 32'sd275477, -32'sd631351, -32'sd79905, -32'sd1454924, -32'sd2018065, -32'sd145032, -32'sd2177920, -32'sd2208173, -32'sd1799380, -32'sd2226275, -32'sd1363320, -32'sd1225968, -32'sd1741418, -32'sd1202106, -32'sd267454, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd55423, -32'sd422393, -32'sd1415731, -32'sd548344, -32'sd1627785, 32'sd500572, 32'sd492285, -32'sd774063, -32'sd1143373, 32'sd684548, -32'sd437815, 32'sd569921, 32'sd652612, -32'sd1424759, -32'sd637232, -32'sd1312151, -32'sd1358374, -32'sd1814060, -32'sd229375, -32'sd54832, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd419850, -32'sd644834, 32'sd874385, 32'sd595174, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1940465, -32'sd1003282, 32'sd1082246, 32'sd342891, 32'sd1323320, 32'sd866883, 32'sd148961, 32'sd1051049, 32'sd1160906, 32'sd1164142, 32'sd446985, 32'sd2560875, 32'sd1276213, 32'sd1319938, 32'sd1670287, 32'sd275655, 32'sd557643, 32'sd1222994, 32'sd265706, 32'sd517196, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1280246, -32'sd22262, 32'sd1683328, -32'sd390925, 32'sd143661, -32'sd646512, 32'sd1430815, 32'sd716249, -32'sd1151342, 32'sd1258192, -32'sd2090225, 32'sd891364, -32'sd1172001, 32'sd933587, 32'sd2403255, 32'sd2118054, 32'sd2345848, 32'sd496535, 32'sd636161, 32'sd1720376, 32'sd415642, 32'sd1178595, 32'sd884375, 32'sd900973, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1118628, 32'sd773020, -32'sd528701, 32'sd1169175, 32'sd766021, 32'sd1582000, 32'sd1091607, 32'sd539305, -32'sd46919, -32'sd1436464, 32'sd18679, 32'sd385994, 32'sd438007, -32'sd1575252, -32'sd301453, 32'sd722542, 32'sd1015564, -32'sd471567, 32'sd1288517, 32'sd1017772, 32'sd533217, 32'sd449186, -32'sd618304, 32'sd665650, 32'sd1888226, 32'sd0, 32'sd0, 32'sd411881, 32'sd245520, -32'sd609621, -32'sd88754, 32'sd2757282, 32'sd707471, 32'sd1288288, -32'sd200289, -32'sd1040885, -32'sd599946, -32'sd1409743, 32'sd1598978, 32'sd2091292, 32'sd1436517, 32'sd728481, -32'sd293260, 32'sd891621, -32'sd675876, 32'sd167464, 32'sd749892, 32'sd357073, 32'sd680576, -32'sd120182, 32'sd849315, 32'sd671455, -32'sd966004, 32'sd194563, 32'sd0, 32'sd873289, 32'sd1475203, 32'sd1187164, 32'sd1425155, 32'sd909459, 32'sd62123, 32'sd652730, 32'sd1172271, 32'sd273863, -32'sd1504891, -32'sd160245, 32'sd559612, 32'sd542412, -32'sd738085, -32'sd916581, 32'sd973976, 32'sd1055984, 32'sd1168832, 32'sd2232222, 32'sd1028141, -32'sd200741, 32'sd586427, -32'sd207982, 32'sd210198, 32'sd635948, 32'sd952193, 32'sd978310, 32'sd0, -32'sd242771, -32'sd186552, 32'sd929401, -32'sd359920, -32'sd892448, -32'sd127806, 32'sd308111, -32'sd619229, 32'sd87294, -32'sd790546, 32'sd1406826, 32'sd1067436, 32'sd144686, -32'sd2457732, -32'sd522845, -32'sd1205843, 32'sd2622815, 32'sd468228, 32'sd581830, 32'sd349893, 32'sd588416, 32'sd339554, 32'sd197935, -32'sd1234355, 32'sd2114468, 32'sd1312469, 32'sd285531, 32'sd1906677, -32'sd17701, 32'sd163319, -32'sd840362, -32'sd509606, 32'sd657024, 32'sd45643, -32'sd462954, 32'sd605118, 32'sd458708, 32'sd1182994, 32'sd1314553, 32'sd1630567, -32'sd1358720, -32'sd205548, 32'sd401425, -32'sd1807319, -32'sd97693, -32'sd2425383, -32'sd2897954, -32'sd211782, 32'sd122161, 32'sd706408, -32'sd30850, 32'sd1481166, 32'sd99123, -32'sd263420, 32'sd97467, 32'sd1299246, 32'sd1026902, 32'sd526967, -32'sd964902, 32'sd690799, -32'sd1106930, -32'sd1622359, 32'sd6987, 32'sd375916, -32'sd1267891, 32'sd672161, 32'sd1320468, -32'sd361656, -32'sd791177, -32'sd1921008, -32'sd328069, 32'sd459335, -32'sd1250364, -32'sd1720884, -32'sd3506834, -32'sd1615434, -32'sd1177445, -32'sd858356, 32'sd1595432, -32'sd1037819, -32'sd1883393, 32'sd295756, 32'sd72541, 32'sd972811, -32'sd232547, 32'sd221951, -32'sd1009324, 32'sd1614787, 32'sd818987, -32'sd243235, 32'sd653419, 32'sd2102050, -32'sd83838, 32'sd1769418, 32'sd406824, -32'sd1476958, -32'sd1265981, 32'sd411817, -32'sd1162809, -32'sd2845992, -32'sd846133, -32'sd2407302, -32'sd2641097, -32'sd2574370, -32'sd2133551, 32'sd144668, 32'sd513163, -32'sd2303587, 32'sd133770, 32'sd1719907, -32'sd267905, 32'sd506441, -32'sd1099309, 32'sd135951, -32'sd808930, 32'sd365509, 32'sd1501015, 32'sd1038902, 32'sd222600, -32'sd325384, 32'sd94934, -32'sd259732, -32'sd335888, -32'sd1204926, -32'sd2405003, -32'sd1343212, -32'sd3336424, -32'sd2787256, -32'sd3879176, -32'sd3463583, -32'sd4403583, -32'sd1068042, -32'sd1583522, -32'sd670868, -32'sd1572644, -32'sd1209496, 32'sd418454, 32'sd738817, 32'sd249207, -32'sd955542, 32'sd729912, -32'sd1487890, 32'sd572473, -32'sd931321, -32'sd1104344, -32'sd1812251, -32'sd860310, -32'sd489301, -32'sd1233604, 32'sd214649, -32'sd2469937, -32'sd1498454, -32'sd1940187, -32'sd849510, -32'sd3208868, -32'sd2693577, -32'sd1776340, -32'sd3578486, -32'sd1784364, -32'sd1448694, -32'sd1941752, 32'sd211894, -32'sd249017, -32'sd419094, 32'sd167416, 32'sd552352, -32'sd121280, 32'sd1194705, 32'sd1015905, 32'sd1167430, 32'sd964531, -32'sd212270, 32'sd395575, -32'sd1773833, -32'sd1648569, 32'sd642937, -32'sd1345842, -32'sd1574156, -32'sd6209, -32'sd768957, -32'sd2095422, -32'sd261941, -32'sd1443059, -32'sd3231937, -32'sd2035383, 32'sd67189, -32'sd1694750, -32'sd2462489, -32'sd3186894, -32'sd2068536, 32'sd944955, 32'sd447504, -32'sd2174397, 32'sd704349, 32'sd298637, 32'sd1600159, 32'sd1021737, 32'sd849567, -32'sd1110744, -32'sd596141, -32'sd5883, 32'sd1060792, 32'sd329976, -32'sd2038477, -32'sd1722066, 32'sd168552, 32'sd1433270, 32'sd10476, 32'sd75644, -32'sd284692, -32'sd1192715, -32'sd659912, 32'sd44300, 32'sd892254, -32'sd1346082, -32'sd2543238, -32'sd635431, -32'sd1399022, 32'sd523152, 32'sd1759516, 32'sd1266020, 32'sd1375608, 32'sd1640118, 32'sd589747, 32'sd597720, 32'sd809174, -32'sd1104328, 32'sd293969, 32'sd809970, -32'sd263893, -32'sd1239333, 32'sd272636, -32'sd409699, 32'sd1745886, 32'sd1265245, 32'sd1163050, 32'sd1115209, 32'sd862259, 32'sd1023479, 32'sd1485476, -32'sd1014132, 32'sd786777, -32'sd1779318, -32'sd84221, 32'sd928113, 32'sd138268, 32'sd703707, -32'sd87391, -32'sd485101, 32'sd2220981, 32'sd233848, 32'sd303468, 32'sd1229878, -32'sd1181833, 32'sd735690, -32'sd564603, 32'sd1625081, 32'sd1806688, -32'sd534249, 32'sd541957, -32'sd1762834, 32'sd106076, -32'sd396232, 32'sd168447, 32'sd1511083, 32'sd997146, 32'sd2610368, 32'sd1966883, 32'sd1355277, 32'sd2017055, -32'sd527533, 32'sd684908, 32'sd642778, -32'sd1437538, -32'sd118544, 32'sd295750, 32'sd957385, 32'sd536574, -32'sd537547, 32'sd1507791, 32'sd200246, -32'sd374033, -32'sd763873, 32'sd487342, 32'sd527686, 32'sd261130, -32'sd158166, -32'sd1411186, -32'sd1614589, -32'sd685426, -32'sd309649, -32'sd1562647, -32'sd241923, 32'sd3009839, 32'sd2261088, 32'sd1998664, 32'sd335070, 32'sd261358, -32'sd1663872, 32'sd2130811, 32'sd486170, -32'sd670376, -32'sd438077, 32'sd379527, 32'sd269379, -32'sd634034, 32'sd621665, 32'sd0, 32'sd459688, 32'sd218455, 32'sd1762728, 32'sd431682, -32'sd777668, 32'sd2063013, 32'sd1253694, 32'sd1178617, -32'sd2386543, -32'sd1527217, -32'sd338137, -32'sd396031, 32'sd1434299, 32'sd3098244, 32'sd804624, 32'sd978114, 32'sd1421280, -32'sd864606, 32'sd382580, 32'sd884471, -32'sd59851, -32'sd798878, 32'sd1205253, 32'sd523708, -32'sd839399, -32'sd2131982, -32'sd982612, 32'sd1427432, 32'sd420628, -32'sd153688, 32'sd148198, 32'sd840681, -32'sd724947, -32'sd66942, -32'sd307600, 32'sd771576, -32'sd750087, -32'sd672209, -32'sd805734, 32'sd370654, 32'sd585779, 32'sd1145963, 32'sd1291912, 32'sd2324842, 32'sd2246800, 32'sd942017, 32'sd653453, -32'sd576066, 32'sd256598, -32'sd1006740, 32'sd698152, 32'sd234662, 32'sd2380936, 32'sd427568, -32'sd391250, 32'sd541745, 32'sd384438, 32'sd1286414, -32'sd1010017, 32'sd997889, -32'sd1060201, -32'sd395103, 32'sd951088, 32'sd2153069, -32'sd946564, -32'sd446007, -32'sd493567, 32'sd1145091, 32'sd1032675, 32'sd1539981, 32'sd984105, 32'sd2418031, 32'sd1835663, 32'sd481216, 32'sd766564, 32'sd704187, -32'sd592729, -32'sd36160, 32'sd1648772, -32'sd1917639, 32'sd1487362, 32'sd1166929, 32'sd420267, 32'sd0, 32'sd420214, 32'sd1228787, 32'sd264114, -32'sd579148, 32'sd850891, -32'sd411711, 32'sd1346204, 32'sd1235053, 32'sd797672, 32'sd824179, 32'sd2162728, 32'sd1044015, 32'sd807889, 32'sd1754420, 32'sd715046, 32'sd965539, -32'sd1075248, 32'sd1741647, 32'sd1777397, 32'sd1624328, 32'sd465673, -32'sd287815, -32'sd132707, 32'sd1659951, -32'sd1409738, -32'sd594206, 32'sd1969937, 32'sd1118515, 32'sd742634, -32'sd53888, -32'sd1020929, 32'sd25919, 32'sd1931600, 32'sd1111218, 32'sd1170839, -32'sd145515, 32'sd2123219, -32'sd366060, -32'sd331695, -32'sd152824, 32'sd909740, 32'sd721610, 32'sd242688, -32'sd248638, 32'sd1228759, 32'sd2106529, 32'sd1156538, 32'sd448474, -32'sd70095, 32'sd340504, -32'sd410942, 32'sd1726577, -32'sd1270377, 32'sd212777, 32'sd225033, 32'sd783420, -32'sd1460915, -32'sd437811, -32'sd8508, 32'sd1903537, 32'sd1397061, -32'sd1523947, 32'sd982600, 32'sd1252943, 32'sd1575137, -32'sd1622488, 32'sd210354, 32'sd630036, -32'sd1601145, -32'sd862222, -32'sd1261557, -32'sd334157, -32'sd406203, -32'sd1347484, -32'sd472616, 32'sd1626617, -32'sd189579, 32'sd269384, -32'sd50216, -32'sd623714, -32'sd198749, 32'sd400907, 32'sd1134073, 32'sd0, -32'sd748296, -32'sd464500, 32'sd225456, 32'sd1018995, -32'sd1213258, 32'sd515060, -32'sd504749, 32'sd58370, 32'sd1221600, -32'sd1594189, 32'sd591149, 32'sd768420, -32'sd756260, -32'sd1974250, -32'sd1461218, -32'sd602095, -32'sd1731764, -32'sd1115733, -32'sd1450155, -32'sd6482, 32'sd210997, 32'sd1206754, 32'sd373988, -32'sd244588, 32'sd760777, -32'sd280950, 32'sd0, 32'sd0, 32'sd0, 32'sd1159477, 32'sd64917, 32'sd1800575, -32'sd32839, -32'sd1164648, -32'sd502865, 32'sd871268, 32'sd14688, -32'sd583807, -32'sd648645, 32'sd107191, -32'sd2388711, -32'sd4864278, -32'sd3410117, -32'sd876839, 32'sd260355, 32'sd139624, -32'sd475678, 32'sd297829, 32'sd163583, 32'sd216061, 32'sd400919, -32'sd678085, 32'sd167713, -32'sd216665, 32'sd0, 32'sd0, 32'sd0, -32'sd1135881, -32'sd487331, 32'sd1465580, 32'sd607522, 32'sd1861933, 32'sd1143134, -32'sd307729, 32'sd1042128, 32'sd1279112, -32'sd763895, -32'sd386375, -32'sd531032, 32'sd88186, -32'sd920809, 32'sd809085, 32'sd1327817, 32'sd941566, -32'sd2448922, -32'sd1293131, 32'sd1518420, 32'sd1659580, -32'sd417979, 32'sd298513, 32'sd1207015, 32'sd1193630, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1182401, -32'sd207736, 32'sd1014656, 32'sd251752, -32'sd1078591, -32'sd296283, 32'sd1249563, 32'sd939466, -32'sd715254, 32'sd1057724, 32'sd1043576, 32'sd1807467, 32'sd2229125, -32'sd895827, 32'sd23008, 32'sd803600, 32'sd572957, -32'sd1238398, -32'sd92153, 32'sd856883, -32'sd104396, 32'sd277092, 32'sd1097435, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1584050, 32'sd1670312, 32'sd957181, 32'sd1473607, 32'sd101715, 32'sd1072175, 32'sd1724835, 32'sd2135884, 32'sd3191853, 32'sd2545411, 32'sd2090724, 32'sd1474921, 32'sd1838522, -32'sd17956, -32'sd126268, -32'sd49726, -32'sd65849, 32'sd64147, 32'sd1793497, 32'sd223509, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1013366, 32'sd792018, -32'sd1027925, -32'sd410350, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1817813, 32'sd1009072, -32'sd796237, -32'sd588679, -32'sd461308, 32'sd826802, 32'sd927637, -32'sd486850, 32'sd1019702, -32'sd535119, 32'sd194202, 32'sd147062, 32'sd767113, 32'sd672147, 32'sd1161123, -32'sd302695, 32'sd654168, -32'sd144175, -32'sd852387, 32'sd93118, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd168267, -32'sd796809, 32'sd669960, -32'sd267200, -32'sd848266, 32'sd1346401, -32'sd139716, 32'sd285540, 32'sd382457, -32'sd644126, 32'sd719469, -32'sd1340392, -32'sd561473, -32'sd238273, -32'sd930771, -32'sd295425, -32'sd1450538, 32'sd1383140, 32'sd1133494, 32'sd513097, -32'sd666573, 32'sd666043, -32'sd167690, 32'sd273792, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd336860, -32'sd1311552, 32'sd2268202, -32'sd877755, 32'sd164880, -32'sd197298, -32'sd16328, -32'sd117018, 32'sd1128347, -32'sd430993, -32'sd2651694, -32'sd682254, 32'sd791410, 32'sd503035, 32'sd796483, -32'sd127660, 32'sd2155347, 32'sd1617955, 32'sd298265, 32'sd527639, 32'sd21115, 32'sd102262, 32'sd876978, -32'sd1178300, -32'sd926446, 32'sd0, 32'sd0, 32'sd781282, 32'sd1177663, 32'sd529947, 32'sd413899, -32'sd263154, -32'sd161527, -32'sd485714, -32'sd2599908, -32'sd998553, 32'sd85577, 32'sd462059, 32'sd1628156, 32'sd125187, 32'sd902506, -32'sd374343, 32'sd1647636, -32'sd1302352, 32'sd498001, 32'sd1130275, 32'sd976338, -32'sd2937, 32'sd169780, -32'sd1141915, -32'sd1348147, 32'sd78120, 32'sd111822, 32'sd1449, 32'sd0, -32'sd74548, -32'sd1345061, -32'sd872952, -32'sd1668413, -32'sd1444105, 32'sd55117, -32'sd598883, -32'sd604873, 32'sd627358, 32'sd653219, 32'sd667023, 32'sd25396, 32'sd200196, -32'sd1343277, -32'sd1427688, -32'sd973709, 32'sd1749400, 32'sd270103, 32'sd748978, -32'sd1415015, 32'sd1043795, 32'sd1637509, -32'sd695360, 32'sd1202297, -32'sd1301880, 32'sd540140, -32'sd957909, 32'sd0, -32'sd528862, 32'sd40895, -32'sd508974, 32'sd173026, 32'sd873470, -32'sd2369583, -32'sd551426, -32'sd689969, 32'sd92851, 32'sd713783, 32'sd2621504, 32'sd339180, 32'sd589430, -32'sd782587, -32'sd2514404, -32'sd2943622, 32'sd482892, 32'sd881235, 32'sd1173473, 32'sd1264586, -32'sd2215330, 32'sd425019, 32'sd1106190, -32'sd830060, 32'sd124006, 32'sd510177, 32'sd1699253, 32'sd195452, 32'sd915245, 32'sd340425, -32'sd2811389, -32'sd787281, -32'sd700702, -32'sd2392025, 32'sd295599, 32'sd1460435, 32'sd1834795, 32'sd379498, 32'sd815780, -32'sd1672508, -32'sd736050, 32'sd783472, -32'sd236094, -32'sd2661634, -32'sd1359893, 32'sd1825174, 32'sd1214554, 32'sd884462, 32'sd1911151, 32'sd1518510, 32'sd100633, -32'sd1441535, -32'sd640863, 32'sd151824, -32'sd294272, -32'sd366394, 32'sd263615, 32'sd1164256, -32'sd1273913, -32'sd668276, -32'sd1879706, 32'sd453967, 32'sd937762, 32'sd964911, 32'sd1889554, -32'sd706255, -32'sd1052871, -32'sd963262, 32'sd208266, -32'sd371872, 32'sd1528850, -32'sd702582, 32'sd369628, 32'sd834747, -32'sd762642, -32'sd636796, 32'sd1092443, 32'sd996713, 32'sd362089, 32'sd739866, 32'sd566576, -32'sd686275, -32'sd795243, -32'sd925039, -32'sd993139, 32'sd1563164, 32'sd635050, -32'sd971181, -32'sd2295627, -32'sd2196517, 32'sd1123997, 32'sd2352468, -32'sd146283, 32'sd940643, 32'sd1684766, -32'sd1988472, -32'sd3033566, -32'sd50390, -32'sd2116027, 32'sd196624, -32'sd1462924, -32'sd2507466, -32'sd2531162, -32'sd3050516, -32'sd728843, -32'sd796153, -32'sd1128078, -32'sd2520909, -32'sd3298053, -32'sd215298, -32'sd943323, -32'sd633999, -32'sd930743, 32'sd494052, -32'sd159333, -32'sd656765, -32'sd1610123, -32'sd1104306, 32'sd1922688, 32'sd2291321, 32'sd2657231, 32'sd2105802, 32'sd1829909, 32'sd187480, -32'sd3612127, -32'sd4655502, -32'sd2331223, 32'sd1441370, -32'sd825938, -32'sd615758, -32'sd78566, -32'sd748398, -32'sd1953393, -32'sd1580909, -32'sd1263148, -32'sd360373, -32'sd2184922, -32'sd14427, 32'sd576794, 32'sd1034347, 32'sd2390162, -32'sd26215, 32'sd282492, 32'sd172199, -32'sd1623267, -32'sd1323453, 32'sd2039335, 32'sd2415105, 32'sd3407793, 32'sd3295951, 32'sd897960, -32'sd1582503, -32'sd2143716, -32'sd733700, 32'sd830124, 32'sd1496326, 32'sd1105503, 32'sd1182637, -32'sd330215, -32'sd1410543, -32'sd1106156, -32'sd1677773, -32'sd2161210, 32'sd481670, -32'sd2456419, -32'sd1305232, -32'sd120103, 32'sd33066, -32'sd1200643, -32'sd1571151, 32'sd628788, -32'sd270408, -32'sd1627730, -32'sd1544810, -32'sd390665, 32'sd2612136, 32'sd4492731, 32'sd763164, 32'sd813683, -32'sd560738, -32'sd2634490, -32'sd1363319, 32'sd2341214, 32'sd1536926, 32'sd1109646, 32'sd468810, 32'sd912074, 32'sd240108, 32'sd757431, 32'sd181525, -32'sd1637617, 32'sd207655, 32'sd763988, -32'sd2391245, -32'sd386106, -32'sd251236, -32'sd463096, 32'sd665, -32'sd326153, 32'sd408807, -32'sd945187, -32'sd907517, 32'sd1401470, 32'sd721172, 32'sd4215277, 32'sd2103225, -32'sd1112306, -32'sd1269694, -32'sd1507343, 32'sd306955, 32'sd2905161, -32'sd928993, -32'sd2027413, 32'sd805865, 32'sd844791, 32'sd2428215, -32'sd870729, 32'sd1036971, 32'sd1509820, 32'sd872958, 32'sd1993602, -32'sd852707, 32'sd259172, 32'sd566949, -32'sd587379, 32'sd292356, -32'sd1866146, -32'sd920017, 32'sd622522, -32'sd622918, 32'sd1105604, 32'sd2348298, 32'sd2042844, 32'sd3142793, 32'sd1559853, -32'sd517890, -32'sd422762, 32'sd725278, -32'sd1906119, 32'sd271469, 32'sd1561605, 32'sd1113045, -32'sd87813, 32'sd1693211, 32'sd600004, 32'sd1987116, 32'sd2020974, 32'sd647577, 32'sd713667, -32'sd1119020, -32'sd974509, -32'sd1218397, -32'sd477036, -32'sd1558238, -32'sd571006, -32'sd630431, 32'sd337453, -32'sd2486698, -32'sd682744, 32'sd2033479, 32'sd2888561, 32'sd3411390, 32'sd2171031, 32'sd3207807, 32'sd397610, -32'sd1099284, -32'sd1925834, -32'sd1609402, 32'sd60097, 32'sd249965, -32'sd463542, 32'sd2605599, 32'sd1282610, -32'sd1649969, 32'sd1009408, 32'sd710982, 32'sd434190, 32'sd245012, -32'sd1188036, 32'sd414833, 32'sd179418, -32'sd968617, -32'sd771504, 32'sd1366924, -32'sd2023769, -32'sd3012537, -32'sd2536397, 32'sd2621186, 32'sd202454, 32'sd1440917, 32'sd2580075, 32'sd1617340, -32'sd1001766, -32'sd2910152, -32'sd515867, 32'sd138495, 32'sd129265, -32'sd957222, 32'sd2149959, -32'sd318197, -32'sd48405, -32'sd1725128, 32'sd300528, -32'sd1700239, 32'sd921617, -32'sd1727570, 32'sd958921, 32'sd0, 32'sd55450, 32'sd520347, 32'sd52239, 32'sd195392, -32'sd2259336, -32'sd1525965, -32'sd2686620, 32'sd609121, -32'sd671185, 32'sd2148184, 32'sd3278094, 32'sd3715896, 32'sd1456320, -32'sd1502400, -32'sd2845412, -32'sd2106378, -32'sd1358503, 32'sd43329, 32'sd1538790, -32'sd878865, -32'sd877768, -32'sd516977, -32'sd31467, 32'sd929901, 32'sd15743, 32'sd896537, 32'sd360103, -32'sd461191, -32'sd384899, 32'sd681242, 32'sd209271, -32'sd495918, -32'sd3056874, -32'sd2530952, -32'sd1691486, -32'sd1161729, 32'sd2275578, 32'sd1018653, -32'sd1237255, 32'sd1392713, -32'sd78672, -32'sd1668850, -32'sd1288055, -32'sd2250863, 32'sd446132, 32'sd320709, 32'sd1363484, 32'sd158081, -32'sd546531, -32'sd228007, 32'sd191344, -32'sd497357, 32'sd183744, 32'sd1006220, -32'sd317928, -32'sd613577, -32'sd951504, -32'sd871043, -32'sd1238248, -32'sd1206619, -32'sd180226, -32'sd539234, -32'sd1148885, -32'sd1438373, -32'sd604528, -32'sd1279737, -32'sd307618, 32'sd321997, 32'sd1726381, 32'sd58505, -32'sd2407183, -32'sd3060235, 32'sd182836, 32'sd2262326, 32'sd426294, -32'sd246271, -32'sd2679928, 32'sd958474, 32'sd1050587, 32'sd840798, -32'sd468967, -32'sd564526, -32'sd1954976, 32'sd0, -32'sd461524, -32'sd866467, -32'sd765057, -32'sd414709, -32'sd1202786, -32'sd750773, -32'sd3375840, -32'sd958132, -32'sd1889483, -32'sd2134201, 32'sd767756, 32'sd738020, 32'sd734143, -32'sd744733, -32'sd1215977, 32'sd762359, 32'sd1972117, 32'sd2356030, 32'sd426784, -32'sd857385, -32'sd723416, 32'sd362703, -32'sd392977, -32'sd624704, -32'sd358392, -32'sd1438823, 32'sd646863, -32'sd663608, -32'sd472441, 32'sd332535, -32'sd1621769, -32'sd169276, 32'sd1354532, -32'sd1919257, -32'sd3174850, -32'sd1628661, -32'sd44567, -32'sd1833357, -32'sd1058215, 32'sd2564823, -32'sd78938, 32'sd450975, -32'sd1663146, -32'sd971425, 32'sd1206527, 32'sd2235244, 32'sd101849, 32'sd1466164, -32'sd511374, 32'sd1358286, 32'sd183118, -32'sd1109002, -32'sd373181, 32'sd770978, -32'sd1204344, -32'sd687489, 32'sd1432382, 32'sd847059, 32'sd134682, -32'sd820848, 32'sd289904, -32'sd2736994, -32'sd3124263, -32'sd2354189, -32'sd1204405, 32'sd879101, 32'sd24687, 32'sd246088, -32'sd1039994, -32'sd53060, 32'sd1237594, 32'sd2430247, 32'sd1091544, 32'sd1205973, 32'sd1087336, -32'sd551186, 32'sd183572, -32'sd2062007, -32'sd1153597, -32'sd1395010, 32'sd721876, -32'sd506693, 32'sd738459, 32'sd0, 32'sd197651, -32'sd1147328, 32'sd1250909, -32'sd917171, 32'sd1385417, -32'sd682850, -32'sd812667, -32'sd1013804, 32'sd57988, 32'sd539796, -32'sd537976, 32'sd1024679, 32'sd285556, 32'sd915346, 32'sd1934376, 32'sd2719182, 32'sd1346933, -32'sd616801, -32'sd1867724, -32'sd1773048, 32'sd109448, -32'sd2752830, 32'sd280299, 32'sd532460, 32'sd840489, 32'sd641273, 32'sd0, 32'sd0, 32'sd0, 32'sd244450, -32'sd150052, -32'sd1006800, -32'sd1014418, -32'sd1472493, 32'sd454303, 32'sd98191, -32'sd334992, -32'sd726203, 32'sd879574, -32'sd1121170, 32'sd364965, -32'sd388350, -32'sd283270, -32'sd380047, -32'sd1716669, -32'sd2443292, -32'sd469794, 32'sd189633, 32'sd410119, -32'sd347777, -32'sd309597, -32'sd412376, -32'sd1529566, -32'sd437596, 32'sd0, 32'sd0, 32'sd0, 32'sd295709, 32'sd628835, -32'sd194588, -32'sd714544, 32'sd701470, 32'sd108669, 32'sd232152, 32'sd2789203, -32'sd147518, -32'sd1408882, -32'sd2432355, -32'sd2112171, -32'sd191909, -32'sd1349670, -32'sd220695, 32'sd1666934, 32'sd1961344, -32'sd292, -32'sd595403, -32'sd486113, 32'sd1075550, 32'sd702701, -32'sd957009, -32'sd880426, 32'sd430830, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd151518, -32'sd450644, -32'sd146729, 32'sd832249, 32'sd627725, 32'sd1199370, 32'sd328714, 32'sd597066, 32'sd1091673, -32'sd83845, 32'sd674353, -32'sd414011, -32'sd2591285, -32'sd1781607, -32'sd386613, -32'sd33774, -32'sd68994, -32'sd1013464, 32'sd416206, 32'sd870351, 32'sd1241788, -32'sd485010, -32'sd443824, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd723040, -32'sd447259, 32'sd1633990, 32'sd464646, 32'sd59714, -32'sd673324, -32'sd235748, 32'sd1171625, 32'sd1560767, 32'sd1563519, -32'sd66593, -32'sd672881, -32'sd1042346, -32'sd236749, -32'sd1299653, -32'sd802443, 32'sd114599, -32'sd1107980, -32'sd1315007, 32'sd345097, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1518077, 32'sd153931, -32'sd435805, -32'sd39125, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd748264, 32'sd771716, -32'sd325719, -32'sd948170, -32'sd1918692, -32'sd540882, 32'sd1731541, 32'sd1270695, 32'sd1646805, 32'sd1462391, 32'sd2078348, 32'sd1713487, 32'sd131473, 32'sd736475, 32'sd1563712, 32'sd308393, 32'sd614676, 32'sd24443, -32'sd41831, 32'sd385606, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1238365, -32'sd257785, 32'sd1210564, -32'sd281415, 32'sd428356, 32'sd56854, 32'sd790773, -32'sd254644, -32'sd341777, -32'sd487555, -32'sd1716663, 32'sd273061, 32'sd2302663, 32'sd1163293, 32'sd415045, 32'sd791008, -32'sd748090, 32'sd16878, 32'sd696639, 32'sd1021222, 32'sd829477, 32'sd1001155, 32'sd942666, 32'sd42318, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd499635, 32'sd495119, -32'sd745483, -32'sd107757, -32'sd1423306, -32'sd731844, -32'sd484157, 32'sd121764, 32'sd1131000, 32'sd430197, -32'sd1106364, 32'sd1801002, 32'sd1374905, 32'sd14097, 32'sd776353, 32'sd1752032, 32'sd1299854, -32'sd173711, 32'sd1566008, 32'sd597043, 32'sd798680, -32'sd776710, 32'sd672177, -32'sd880092, 32'sd83735, 32'sd0, 32'sd0, 32'sd1208429, 32'sd569589, -32'sd386247, -32'sd2307983, -32'sd184592, 32'sd1014669, 32'sd639942, -32'sd574376, 32'sd2251966, 32'sd1221635, 32'sd109001, -32'sd474306, 32'sd176911, -32'sd263649, -32'sd1306985, 32'sd502307, -32'sd1328794, 32'sd224780, 32'sd1178510, 32'sd2384319, -32'sd302622, 32'sd573569, 32'sd1724011, -32'sd460482, 32'sd274508, 32'sd189117, 32'sd828818, 32'sd0, 32'sd368434, 32'sd1329285, 32'sd1113286, -32'sd168732, -32'sd1913345, -32'sd479343, -32'sd2036918, 32'sd1075370, -32'sd32379, 32'sd1262208, -32'sd169395, -32'sd425915, -32'sd330204, -32'sd265685, -32'sd180888, -32'sd2892539, -32'sd2075483, -32'sd1183414, -32'sd184688, -32'sd2132520, -32'sd1987365, -32'sd167733, 32'sd1122491, 32'sd191842, 32'sd839831, 32'sd940276, 32'sd177546, 32'sd0, 32'sd853904, 32'sd651567, 32'sd728084, 32'sd1460152, 32'sd671592, 32'sd1346137, 32'sd1458598, -32'sd559988, -32'sd921605, -32'sd639474, 32'sd450917, -32'sd1318473, -32'sd191596, -32'sd1451146, -32'sd558553, 32'sd763419, -32'sd784761, -32'sd212211, -32'sd1373447, -32'sd529612, 32'sd36382, -32'sd519029, 32'sd692671, -32'sd142999, 32'sd723304, 32'sd782246, -32'sd1041249, 32'sd950977, 32'sd3511, -32'sd612247, -32'sd1399406, 32'sd1103159, 32'sd1503212, 32'sd350749, 32'sd1038946, 32'sd75589, 32'sd74020, -32'sd766157, -32'sd1311706, -32'sd77103, -32'sd2361308, -32'sd2391148, 32'sd486282, 32'sd1343203, 32'sd901386, 32'sd292209, -32'sd367567, -32'sd453160, 32'sd266977, 32'sd304402, 32'sd435730, 32'sd1904191, -32'sd1031367, 32'sd602659, -32'sd169640, 32'sd169403, 32'sd747765, 32'sd257050, 32'sd853100, 32'sd1315858, 32'sd655700, -32'sd4467, 32'sd2130526, 32'sd2234192, 32'sd1737981, 32'sd1152743, 32'sd782230, -32'sd829272, -32'sd2948400, 32'sd301750, 32'sd1920005, 32'sd3903970, 32'sd710532, 32'sd157527, 32'sd223885, -32'sd355188, 32'sd277121, -32'sd234786, -32'sd416988, 32'sd1877260, -32'sd1669086, -32'sd1197826, 32'sd101829, 32'sd1876709, 32'sd1537926, -32'sd61985, 32'sd97725, 32'sd1085721, 32'sd1000952, -32'sd722974, 32'sd496934, 32'sd2238024, 32'sd457748, 32'sd1856047, -32'sd1063153, -32'sd3669314, -32'sd1348016, 32'sd954093, 32'sd520401, 32'sd1860396, -32'sd1060845, 32'sd956951, 32'sd2402795, 32'sd3194411, 32'sd463527, 32'sd664747, 32'sd1238983, -32'sd112830, 32'sd1227358, -32'sd629472, -32'sd32038, 32'sd1691594, -32'sd130354, 32'sd1531464, -32'sd1169106, 32'sd2252599, 32'sd1124090, -32'sd521491, -32'sd493288, 32'sd917092, 32'sd1140637, 32'sd2104178, 32'sd2235090, -32'sd1532173, -32'sd1638943, -32'sd2360919, -32'sd379453, 32'sd1176181, 32'sd27347, 32'sd2082240, 32'sd1617643, 32'sd1849162, 32'sd1088126, 32'sd1424466, 32'sd388057, 32'sd533202, -32'sd544908, -32'sd769261, -32'sd1541542, 32'sd135589, 32'sd30595, -32'sd608648, -32'sd188055, 32'sd629929, 32'sd55569, 32'sd78186, -32'sd454525, 32'sd1620171, 32'sd3259756, 32'sd1713610, 32'sd2452158, -32'sd1383290, -32'sd3493823, -32'sd1358944, -32'sd1677085, -32'sd180621, 32'sd2108725, -32'sd177469, 32'sd359512, 32'sd1713985, -32'sd515377, 32'sd871019, -32'sd289844, 32'sd738151, 32'sd302098, -32'sd50857, 32'sd305126, 32'sd607164, 32'sd791739, 32'sd1271829, -32'sd473937, -32'sd611874, 32'sd1331940, 32'sd903168, 32'sd2265522, 32'sd697754, 32'sd3056053, 32'sd4081642, 32'sd762318, -32'sd355704, -32'sd4072293, -32'sd6176098, -32'sd2037769, 32'sd2221735, -32'sd94538, 32'sd1073030, -32'sd1329036, 32'sd126148, 32'sd209858, 32'sd360865, 32'sd1700739, 32'sd922848, 32'sd173888, 32'sd2307228, 32'sd1533210, 32'sd988061, 32'sd481741, 32'sd381293, 32'sd630903, 32'sd201753, 32'sd1406233, 32'sd2115744, 32'sd2527565, 32'sd4132459, 32'sd2181138, 32'sd4336053, 32'sd1851890, -32'sd3405568, -32'sd4934356, -32'sd5987179, -32'sd1247784, -32'sd214833, -32'sd431921, 32'sd251880, -32'sd321206, 32'sd662384, 32'sd1875441, 32'sd1198766, 32'sd2345316, 32'sd277567, 32'sd1003112, 32'sd1956397, -32'sd1800752, 32'sd388674, 32'sd1394707, 32'sd1408965, 32'sd606159, 32'sd456373, 32'sd2039323, 32'sd1990716, 32'sd2935480, 32'sd1616572, 32'sd3597185, 32'sd2624167, 32'sd34455, -32'sd1371832, -32'sd4527540, -32'sd3268208, -32'sd2081556, 32'sd603472, -32'sd563256, 32'sd686284, -32'sd1377865, 32'sd115927, 32'sd339655, 32'sd1492552, 32'sd1227766, -32'sd41212, 32'sd865351, -32'sd757727, 32'sd305170, 32'sd1450172, -32'sd921158, 32'sd473799, -32'sd1059861, -32'sd1657361, 32'sd558171, 32'sd1726888, 32'sd1897160, 32'sd460061, 32'sd2110299, -32'sd851173, -32'sd2382742, -32'sd4146554, -32'sd4462685, -32'sd3692155, -32'sd2133242, -32'sd1919209, -32'sd2738495, -32'sd1084292, 32'sd364665, -32'sd406724, 32'sd515903, 32'sd880164, 32'sd996638, -32'sd1382936, 32'sd1376919, -32'sd115424, 32'sd457874, 32'sd523527, 32'sd721117, 32'sd229085, 32'sd791065, -32'sd391959, -32'sd214007, 32'sd2379523, 32'sd1782230, 32'sd2290090, -32'sd1620349, -32'sd1687164, -32'sd3969803, -32'sd5608488, -32'sd4447509, -32'sd1750747, 32'sd370339, -32'sd2273108, -32'sd1538873, -32'sd750228, -32'sd550511, 32'sd899456, 32'sd1537037, 32'sd1044777, -32'sd1306076, -32'sd1009278, 32'sd2369214, -32'sd139473, 32'sd718253, 32'sd0, -32'sd671216, 32'sd1073744, 32'sd1149432, 32'sd2044828, 32'sd1723592, 32'sd1168587, 32'sd773734, 32'sd70752, 32'sd788882, -32'sd2895233, -32'sd4285206, -32'sd3656972, -32'sd2844140, -32'sd624108, -32'sd804231, 32'sd1038926, -32'sd1164065, 32'sd1194622, 32'sd1216455, 32'sd143305, 32'sd675704, -32'sd1100683, 32'sd89001, 32'sd886504, 32'sd1183338, -32'sd164386, -32'sd767772, 32'sd717755, -32'sd1050674, 32'sd117755, 32'sd132844, 32'sd435104, -32'sd142479, -32'sd197066, 32'sd146077, 32'sd1005819, 32'sd627884, 32'sd462379, -32'sd2822569, -32'sd4074760, -32'sd1117372, -32'sd438214, -32'sd1119869, -32'sd391612, -32'sd124345, 32'sd1676744, 32'sd152121, 32'sd1240780, 32'sd90775, -32'sd434854, -32'sd1110682, 32'sd1893978, 32'sd854972, -32'sd1463379, 32'sd750130, 32'sd456328, 32'sd1041221, 32'sd452651, 32'sd1010649, 32'sd471188, 32'sd426, -32'sd130855, -32'sd173543, -32'sd438501, 32'sd24742, -32'sd12042, -32'sd2582246, -32'sd447208, 32'sd18767, 32'sd1646795, -32'sd1157496, -32'sd1975488, -32'sd2175296, 32'sd1842267, -32'sd1106284, -32'sd936510, -32'sd1261436, -32'sd1281405, -32'sd468180, 32'sd1147683, 32'sd31409, -32'sd1183021, -32'sd211657, 32'sd0, 32'sd1577999, 32'sd309479, 32'sd1230167, -32'sd1032863, 32'sd322380, 32'sd14959, 32'sd1223324, -32'sd287626, -32'sd615984, 32'sd747990, -32'sd1665416, -32'sd568335, 32'sd281903, -32'sd1539735, -32'sd297822, 32'sd462153, 32'sd888435, 32'sd1460300, 32'sd1033221, -32'sd7065, -32'sd217721, -32'sd485826, -32'sd3698291, -32'sd1442718, 32'sd242552, 32'sd1277773, -32'sd302360, 32'sd731267, 32'sd1200394, 32'sd542892, 32'sd484292, -32'sd45202, 32'sd131018, -32'sd1488791, 32'sd614388, 32'sd743079, -32'sd386459, 32'sd242112, 32'sd2157306, 32'sd706205, -32'sd566754, -32'sd1623579, -32'sd563930, 32'sd362365, -32'sd929721, 32'sd810096, -32'sd134929, -32'sd1095120, -32'sd16764, 32'sd512242, -32'sd1369313, 32'sd632302, 32'sd1248387, 32'sd651730, 32'sd437497, -32'sd345957, 32'sd855527, 32'sd988974, -32'sd1437652, 32'sd297137, 32'sd432912, -32'sd130756, -32'sd865347, 32'sd1126073, -32'sd934970, 32'sd761233, 32'sd43150, -32'sd224850, 32'sd1406158, 32'sd11754, -32'sd915725, 32'sd66468, 32'sd429621, -32'sd1150092, -32'sd1500770, -32'sd326729, 32'sd474798, -32'sd879564, -32'sd248668, -32'sd1215691, 32'sd1835873, 32'sd615945, 32'sd514359, 32'sd0, 32'sd697125, -32'sd1079784, -32'sd612824, 32'sd1197630, 32'sd640039, 32'sd1412590, 32'sd211323, 32'sd1662618, 32'sd1109702, -32'sd21418, -32'sd1098274, 32'sd548474, 32'sd550134, 32'sd113726, -32'sd510026, -32'sd374242, 32'sd393983, -32'sd371933, -32'sd685218, 32'sd1123701, 32'sd451256, 32'sd775440, 32'sd440420, 32'sd88657, 32'sd1133879, 32'sd658283, 32'sd0, 32'sd0, 32'sd0, 32'sd569765, 32'sd1034147, 32'sd1305613, 32'sd2164685, 32'sd894997, -32'sd536007, 32'sd67434, 32'sd767486, -32'sd1419147, -32'sd468909, 32'sd1182563, -32'sd560619, -32'sd1338168, 32'sd136402, -32'sd501354, 32'sd513666, 32'sd154038, -32'sd924903, -32'sd1241086, 32'sd1515873, -32'sd989160, -32'sd1661579, 32'sd1100668, 32'sd1022124, 32'sd977627, 32'sd0, 32'sd0, 32'sd0, -32'sd346708, 32'sd6837, 32'sd1158151, 32'sd600132, 32'sd841280, -32'sd1098417, 32'sd1642013, 32'sd466855, -32'sd219116, 32'sd808661, 32'sd1909737, 32'sd681896, 32'sd310030, -32'sd118393, 32'sd2996198, 32'sd387426, 32'sd348341, -32'sd1806865, -32'sd1120922, 32'sd270740, 32'sd831091, 32'sd1165418, -32'sd590612, -32'sd49788, 32'sd374085, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd95682, -32'sd869915, 32'sd1405795, 32'sd133778, 32'sd132540, 32'sd1064674, -32'sd887327, -32'sd1317665, -32'sd749448, 32'sd826378, 32'sd921678, -32'sd718277, -32'sd784467, 32'sd545620, 32'sd1214821, -32'sd673040, 32'sd1397196, 32'sd1573467, -32'sd117900, 32'sd849524, -32'sd514677, 32'sd1892599, 32'sd1483955, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1770179, 32'sd926368, -32'sd29773, 32'sd623578, -32'sd189635, 32'sd28735, 32'sd1041623, 32'sd680932, 32'sd1537857, 32'sd303174, -32'sd17267, 32'sd191451, 32'sd3795, 32'sd186925, -32'sd809007, 32'sd31115, -32'sd1930355, -32'sd547250, 32'sd565675, 32'sd655577, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd356646, -32'sd173567, 32'sd460439, -32'sd801581, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd755367, 32'sd751001, -32'sd452426, -32'sd641153, -32'sd664101, 32'sd115395, 32'sd545367, -32'sd158555, 32'sd735150, 32'sd14530, 32'sd1882792, 32'sd103123, -32'sd417528, 32'sd835719, -32'sd68888, -32'sd1255601, -32'sd80775, -32'sd1124252, -32'sd1357709, 32'sd679092, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd106943, -32'sd564175, 32'sd577781, -32'sd923639, -32'sd959490, 32'sd751054, 32'sd564926, -32'sd273515, 32'sd1114901, 32'sd1211146, -32'sd858527, 32'sd1074810, 32'sd294944, -32'sd458388, -32'sd1528348, -32'sd862958, -32'sd1689345, -32'sd1868846, -32'sd2197728, -32'sd408535, -32'sd162008, -32'sd474696, -32'sd923803, -32'sd837049, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd350821, 32'sd857681, 32'sd457852, -32'sd1463617, -32'sd735134, -32'sd1649947, -32'sd159506, 32'sd973431, -32'sd216804, -32'sd3259510, -32'sd793228, -32'sd253255, -32'sd1119907, 32'sd552845, 32'sd1060521, 32'sd597316, 32'sd439268, -32'sd6019, -32'sd795503, -32'sd417451, 32'sd381791, -32'sd128460, -32'sd1621821, -32'sd67516, -32'sd116028, 32'sd0, 32'sd0, -32'sd745344, -32'sd563057, -32'sd959872, -32'sd456451, 32'sd217429, 32'sd474886, -32'sd321558, -32'sd1090939, -32'sd720589, -32'sd755314, 32'sd204233, 32'sd1050213, 32'sd820188, 32'sd1925989, -32'sd163460, 32'sd915942, 32'sd102925, 32'sd1867332, 32'sd1916145, 32'sd1594434, -32'sd953903, -32'sd419391, -32'sd456638, -32'sd1117255, -32'sd1304000, -32'sd86625, 32'sd360137, 32'sd0, 32'sd65361, 32'sd182008, -32'sd1251850, -32'sd933135, 32'sd1580577, 32'sd892310, -32'sd2338441, -32'sd730095, 32'sd700272, -32'sd492567, 32'sd1823108, 32'sd285664, 32'sd956357, 32'sd1822234, 32'sd1214681, 32'sd639427, 32'sd2134490, 32'sd1111371, -32'sd781239, 32'sd1302803, 32'sd487401, 32'sd313562, -32'sd509858, -32'sd1500199, 32'sd1290774, 32'sd1750498, -32'sd37184, 32'sd0, -32'sd40334, -32'sd683866, 32'sd890865, 32'sd545824, -32'sd1193563, -32'sd648291, 32'sd351297, -32'sd1340087, -32'sd516313, 32'sd206649, 32'sd1856025, 32'sd1729553, 32'sd336270, -32'sd949529, 32'sd1424843, 32'sd2486877, 32'sd3338188, 32'sd662252, 32'sd2399679, 32'sd887310, 32'sd1168176, 32'sd760715, 32'sd441476, -32'sd1128615, -32'sd904023, -32'sd412731, -32'sd460576, -32'sd338450, -32'sd4466, 32'sd684513, -32'sd75775, 32'sd436238, -32'sd365225, -32'sd725177, -32'sd1338303, -32'sd2930562, -32'sd735800, 32'sd1239627, 32'sd808409, 32'sd355788, -32'sd222307, -32'sd1076264, -32'sd451911, 32'sd278444, 32'sd1452757, 32'sd1420306, 32'sd1109082, 32'sd1378285, 32'sd1585319, -32'sd281149, 32'sd495901, -32'sd739422, 32'sd425201, -32'sd489416, -32'sd431597, 32'sd672816, -32'sd436323, 32'sd1218302, -32'sd700369, -32'sd567454, -32'sd1227226, -32'sd1165866, -32'sd337461, 32'sd587866, 32'sd2016203, 32'sd1399616, 32'sd1023081, 32'sd38400, -32'sd57038, -32'sd85744, 32'sd236878, 32'sd220857, 32'sd1290384, 32'sd1475969, 32'sd2214136, 32'sd2247896, -32'sd13757, 32'sd70261, 32'sd1267665, -32'sd658723, -32'sd506113, -32'sd1438474, 32'sd736198, -32'sd347701, -32'sd806782, 32'sd1656732, 32'sd2630973, 32'sd469178, 32'sd1680545, 32'sd2145526, 32'sd1025768, 32'sd2290867, 32'sd1956507, 32'sd1139365, -32'sd2294662, -32'sd3121960, -32'sd1781806, -32'sd1601938, -32'sd368489, 32'sd230590, -32'sd1890725, 32'sd1242677, 32'sd757599, 32'sd905233, -32'sd73508, -32'sd22349, -32'sd67835, 32'sd903650, 32'sd167694, 32'sd524547, -32'sd524966, -32'sd861833, 32'sd685397, 32'sd1259603, 32'sd1206735, 32'sd1125884, 32'sd3030664, -32'sd92831, 32'sd2362525, 32'sd2275630, -32'sd583128, -32'sd419044, -32'sd1073158, -32'sd1262541, -32'sd2911712, -32'sd1237826, 32'sd599866, -32'sd740719, 32'sd414084, 32'sd1670402, -32'sd843477, 32'sd619229, -32'sd139441, 32'sd1898379, 32'sd1219316, -32'sd284822, 32'sd773500, 32'sd685044, 32'sd795461, 32'sd68014, -32'sd1638601, -32'sd1544, 32'sd1541332, -32'sd969082, 32'sd1495206, 32'sd885345, 32'sd2086705, 32'sd265340, -32'sd76638, -32'sd220995, 32'sd1499833, 32'sd658696, 32'sd730451, -32'sd2172059, -32'sd1556812, -32'sd725990, -32'sd1952595, -32'sd2478300, 32'sd40995, 32'sd1043889, 32'sd2595988, 32'sd2265194, 32'sd2145558, -32'sd385982, -32'sd357979, 32'sd218649, 32'sd1707363, -32'sd8045, -32'sd807704, -32'sd384109, 32'sd1877272, -32'sd1427283, -32'sd810962, 32'sd2389603, 32'sd1210477, -32'sd1665478, 32'sd179060, 32'sd1104417, 32'sd1889330, 32'sd1194046, -32'sd1763417, -32'sd1989586, -32'sd3247539, -32'sd2493790, 32'sd199410, -32'sd2026487, -32'sd720759, 32'sd2172019, 32'sd914885, 32'sd1572831, 32'sd1364202, 32'sd469414, 32'sd464232, -32'sd1462292, 32'sd1177621, 32'sd392972, 32'sd119850, 32'sd530502, 32'sd2264239, -32'sd594710, -32'sd703360, 32'sd341396, -32'sd1608221, 32'sd891003, -32'sd256282, -32'sd543164, -32'sd147197, -32'sd887039, 32'sd213444, -32'sd938476, -32'sd841262, 32'sd293508, -32'sd1151923, -32'sd1280504, 32'sd420687, 32'sd1781227, 32'sd3154686, 32'sd1382598, 32'sd163720, -32'sd1882032, -32'sd1295731, -32'sd1574791, 32'sd1524488, 32'sd207416, -32'sd208165, -32'sd1571417, -32'sd714268, 32'sd1422291, -32'sd59054, -32'sd1489508, 32'sd322855, -32'sd2970171, -32'sd2954060, -32'sd1400547, -32'sd1393818, -32'sd1422343, 32'sd1555431, -32'sd30378, 32'sd891446, 32'sd1038637, -32'sd1012565, -32'sd1864492, -32'sd913332, -32'sd409855, 32'sd1081257, 32'sd69548, -32'sd955203, -32'sd2265878, 32'sd1292325, 32'sd2243181, -32'sd46367, -32'sd165795, -32'sd634210, -32'sd275506, 32'sd1100018, 32'sd147037, 32'sd244050, -32'sd161952, -32'sd490143, -32'sd967673, 32'sd952728, -32'sd643287, 32'sd556746, 32'sd732294, 32'sd504734, -32'sd1045856, -32'sd247408, -32'sd653237, -32'sd1451786, -32'sd1493158, -32'sd1226931, 32'sd729002, 32'sd1557715, 32'sd83386, -32'sd2396439, -32'sd241570, -32'sd2138217, 32'sd204604, 32'sd361797, 32'sd436166, 32'sd818383, -32'sd930904, 32'sd1790729, 32'sd616524, -32'sd1494154, 32'sd1096349, -32'sd1372909, 32'sd1582479, -32'sd269174, 32'sd717242, 32'sd1192101, 32'sd2849231, 32'sd2686279, -32'sd1888843, 32'sd203527, 32'sd642474, -32'sd1830133, -32'sd1635323, 32'sd142458, -32'sd1420876, 32'sd155706, -32'sd543959, -32'sd239417, 32'sd920503, 32'sd853693, -32'sd869721, 32'sd20318, 32'sd0, 32'sd605601, 32'sd665117, 32'sd1516287, 32'sd1609852, -32'sd461451, 32'sd1362977, 32'sd125089, 32'sd591240, 32'sd97585, 32'sd1027688, 32'sd3765591, 32'sd3276793, 32'sd2349632, -32'sd613411, -32'sd3744225, -32'sd3393874, -32'sd2612005, -32'sd3058381, -32'sd1598109, -32'sd355896, -32'sd2618507, -32'sd1312444, 32'sd800683, -32'sd707041, 32'sd566150, 32'sd1130627, -32'sd13422, -32'sd695728, 32'sd274343, 32'sd450278, -32'sd148926, 32'sd262937, -32'sd314290, 32'sd935800, -32'sd223045, 32'sd137142, 32'sd2059952, 32'sd2178589, 32'sd4122835, 32'sd1760352, -32'sd961807, -32'sd3397608, -32'sd5442987, -32'sd3332978, -32'sd472125, -32'sd158443, -32'sd2961315, -32'sd1730636, -32'sd1910135, 32'sd465604, -32'sd367853, 32'sd1446222, -32'sd816566, 32'sd427586, -32'sd1132478, -32'sd673574, -32'sd568691, -32'sd716147, -32'sd1602451, 32'sd673859, -32'sd1756287, 32'sd454252, -32'sd51743, 32'sd881715, 32'sd2152300, 32'sd2858389, 32'sd2831003, 32'sd1292135, 32'sd818163, -32'sd5015799, -32'sd3431996, -32'sd995004, 32'sd558012, -32'sd1379705, -32'sd2911493, -32'sd616450, -32'sd641357, 32'sd735990, 32'sd1173835, 32'sd129671, 32'sd126645, 32'sd196723, 32'sd153764, 32'sd0, -32'sd1402024, 32'sd1697315, 32'sd1381968, 32'sd272384, -32'sd26590, 32'sd1394085, 32'sd1980060, 32'sd3894192, 32'sd2438573, 32'sd2228263, 32'sd2802945, 32'sd981061, -32'sd1253832, -32'sd5568046, -32'sd876694, 32'sd890668, 32'sd481238, 32'sd557690, 32'sd208063, -32'sd1183405, 32'sd535946, -32'sd1642240, 32'sd28479, 32'sd1648202, 32'sd889876, 32'sd998436, 32'sd885594, -32'sd712944, -32'sd728371, 32'sd527248, -32'sd22428, 32'sd698944, 32'sd781837, 32'sd1522836, 32'sd744299, 32'sd978833, 32'sd2054439, 32'sd2182278, 32'sd1370403, -32'sd368731, -32'sd4280824, -32'sd2558202, -32'sd1177595, 32'sd581521, 32'sd1650257, 32'sd616699, -32'sd228119, -32'sd722901, 32'sd1060306, -32'sd173661, -32'sd2144368, 32'sd616320, 32'sd244148, 32'sd1630783, -32'sd117289, -32'sd488653, 32'sd385807, -32'sd587109, -32'sd1443608, -32'sd587371, 32'sd731916, 32'sd2547557, 32'sd1524199, 32'sd1511176, 32'sd2404018, 32'sd2121670, -32'sd784646, -32'sd1547686, -32'sd2711529, -32'sd791862, -32'sd486073, -32'sd1899924, 32'sd1444688, 32'sd2116406, 32'sd329259, 32'sd1917094, 32'sd65382, 32'sd583255, -32'sd2267472, -32'sd1639215, -32'sd65822, 32'sd829290, 32'sd1464528, 32'sd0, -32'sd215425, -32'sd1234695, -32'sd2236664, -32'sd83213, 32'sd309060, 32'sd712423, 32'sd1918296, 32'sd2413620, 32'sd1968278, 32'sd702420, 32'sd1094857, -32'sd755772, -32'sd909518, -32'sd1507580, -32'sd1077321, -32'sd1393751, -32'sd1573312, -32'sd471129, 32'sd1340145, -32'sd1329623, -32'sd282067, 32'sd241156, -32'sd1891917, -32'sd733338, -32'sd144481, 32'sd395283, 32'sd0, 32'sd0, 32'sd0, -32'sd374680, -32'sd748275, -32'sd801603, 32'sd615158, 32'sd279696, 32'sd1291508, 32'sd1760902, 32'sd998050, 32'sd1095223, 32'sd836356, 32'sd2388782, 32'sd644951, -32'sd629579, -32'sd2268767, -32'sd3560301, -32'sd1923063, 32'sd576460, 32'sd1677826, -32'sd660873, 32'sd256823, 32'sd706600, -32'sd636646, 32'sd217355, 32'sd1707720, -32'sd493368, 32'sd0, 32'sd0, 32'sd0, -32'sd123309, 32'sd422719, 32'sd180849, -32'sd609509, 32'sd926674, 32'sd1153306, 32'sd639744, 32'sd2753612, 32'sd1026765, -32'sd1381649, 32'sd121526, -32'sd492056, 32'sd593117, -32'sd2299283, -32'sd3068629, -32'sd1931366, -32'sd939588, 32'sd366141, 32'sd195184, 32'sd1588722, -32'sd208837, 32'sd1118375, 32'sd730588, -32'sd1076838, 32'sd904819, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd559684, 32'sd1301310, 32'sd914754, 32'sd369479, 32'sd589307, 32'sd646727, -32'sd417533, -32'sd216652, -32'sd2573125, -32'sd1127128, 32'sd40262, 32'sd389647, 32'sd93487, -32'sd947708, -32'sd25907, 32'sd187227, 32'sd1076091, 32'sd953151, 32'sd500141, 32'sd208493, -32'sd343999, 32'sd152907, -32'sd765354, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd333649, -32'sd639826, -32'sd172358, -32'sd479485, -32'sd1371170, -32'sd897502, 32'sd441846, -32'sd511318, 32'sd736947, 32'sd84476, 32'sd1119153, -32'sd559477, 32'sd469036, -32'sd1324788, -32'sd696777, 32'sd530050, -32'sd1437897, 32'sd279580, 32'sd1268462, 32'sd1350093, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd341873, -32'sd204485, 32'sd1295518, 32'sd1866507, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1169352, 32'sd226813, 32'sd1575041, 32'sd24179, 32'sd373368, -32'sd396043, -32'sd467167, 32'sd1828742, 32'sd962928, 32'sd955614, -32'sd1731885, -32'sd189467, 32'sd1313906, -32'sd352333, -32'sd1393161, -32'sd840205, -32'sd715821, -32'sd509436, 32'sd151422, -32'sd96325, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd123086, -32'sd267778, 32'sd42582, 32'sd1809749, -32'sd399056, 32'sd23311, 32'sd109101, -32'sd525804, 32'sd464386, 32'sd2492897, 32'sd1453653, 32'sd454215, -32'sd203356, -32'sd1883175, -32'sd409356, -32'sd223559, -32'sd1069248, -32'sd1837706, -32'sd2513877, -32'sd1559514, -32'sd171700, -32'sd416028, -32'sd687309, 32'sd270362, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd795643, 32'sd1089308, -32'sd570459, 32'sd763610, 32'sd137779, -32'sd417350, 32'sd2248080, 32'sd1907771, 32'sd464103, 32'sd2084764, 32'sd2929218, -32'sd1002565, 32'sd866488, 32'sd1307008, -32'sd462693, 32'sd461706, 32'sd1237840, -32'sd694118, 32'sd1344635, -32'sd1274687, -32'sd1091298, -32'sd1945802, 32'sd441533, 32'sd453674, -32'sd338940, 32'sd0, 32'sd0, -32'sd377206, 32'sd843598, -32'sd595931, 32'sd578739, 32'sd293840, 32'sd1132159, 32'sd1145250, 32'sd936688, 32'sd1047053, 32'sd344723, 32'sd2413322, 32'sd1969415, 32'sd749508, 32'sd92924, 32'sd1291146, -32'sd579168, 32'sd806593, 32'sd1426532, 32'sd1083451, 32'sd588062, -32'sd1784728, -32'sd1551030, -32'sd1537415, -32'sd1275846, -32'sd761449, -32'sd1065703, -32'sd535027, 32'sd0, -32'sd874255, 32'sd871402, 32'sd1429265, 32'sd1578351, -32'sd347945, -32'sd568904, -32'sd815157, 32'sd745615, 32'sd114558, 32'sd778576, -32'sd2778869, -32'sd3149171, -32'sd544793, -32'sd21443, 32'sd1276335, -32'sd900803, -32'sd1613166, -32'sd430103, 32'sd2038955, 32'sd1336889, -32'sd433156, 32'sd1874751, 32'sd2994247, -32'sd1152700, -32'sd2286024, 32'sd270323, 32'sd381997, 32'sd0, 32'sd129552, 32'sd686204, 32'sd175136, 32'sd626548, 32'sd484120, 32'sd1565575, 32'sd1463213, 32'sd486487, 32'sd1204088, -32'sd52931, -32'sd1234862, -32'sd513830, 32'sd461235, 32'sd894506, -32'sd950669, -32'sd1021240, -32'sd2118513, -32'sd810072, -32'sd1563549, 32'sd46570, -32'sd901363, 32'sd1729351, 32'sd2363596, -32'sd83868, 32'sd1269771, 32'sd269443, -32'sd1646251, -32'sd174435, -32'sd368846, -32'sd2672902, -32'sd962399, 32'sd1086455, 32'sd1580002, 32'sd3322990, 32'sd2428712, 32'sd274658, -32'sd2348614, -32'sd443840, 32'sd536844, 32'sd958006, -32'sd240326, -32'sd512472, -32'sd433575, -32'sd1079056, -32'sd487663, -32'sd1580342, -32'sd360079, -32'sd860451, 32'sd429425, 32'sd446575, 32'sd418, 32'sd277993, -32'sd593094, 32'sd2004224, 32'sd26157, -32'sd241999, -32'sd322638, -32'sd874290, -32'sd2728472, -32'sd803261, 32'sd1084465, -32'sd882211, -32'sd3184806, -32'sd2231040, -32'sd5406617, -32'sd1347332, 32'sd107190, -32'sd1046553, -32'sd2422776, -32'sd1158265, -32'sd1224817, -32'sd141884, 32'sd609185, 32'sd1670583, 32'sd1005054, 32'sd306740, 32'sd1008155, 32'sd448480, 32'sd1027214, -32'sd1034590, 32'sd854091, 32'sd1867705, -32'sd1391213, 32'sd73414, -32'sd1554487, 32'sd723161, 32'sd1006231, -32'sd405451, 32'sd171717, -32'sd3400611, -32'sd6383314, -32'sd4240891, -32'sd4263800, -32'sd2431992, 32'sd214893, 32'sd412910, -32'sd1009899, -32'sd1697254, -32'sd1577259, 32'sd575007, 32'sd819317, 32'sd2784503, 32'sd2047365, 32'sd614773, -32'sd281815, -32'sd197929, -32'sd346803, 32'sd286511, -32'sd1884179, 32'sd1299083, 32'sd369766, -32'sd180028, -32'sd154784, 32'sd312566, 32'sd1956013, -32'sd1246668, -32'sd2540256, -32'sd1805628, -32'sd3160973, -32'sd3332357, 32'sd21369, -32'sd560930, -32'sd1051013, 32'sd1151477, 32'sd1283059, -32'sd2180099, -32'sd693634, 32'sd2036396, 32'sd326761, 32'sd1666094, 32'sd2418217, 32'sd683354, 32'sd1608866, -32'sd969740, 32'sd545188, 32'sd272546, -32'sd1546421, 32'sd1709502, -32'sd368054, -32'sd1415734, -32'sd914416, -32'sd316767, -32'sd1454722, 32'sd1813040, -32'sd1219699, 32'sd779598, -32'sd555538, -32'sd978198, -32'sd532192, -32'sd316687, -32'sd71623, 32'sd1835838, 32'sd450024, -32'sd614444, 32'sd600297, 32'sd377656, 32'sd969444, 32'sd372037, 32'sd1037014, -32'sd573511, -32'sd1311922, -32'sd1917683, -32'sd709034, -32'sd1544819, -32'sd1959362, -32'sd1709760, -32'sd151072, 32'sd486711, -32'sd101607, -32'sd1182877, -32'sd340707, 32'sd786899, 32'sd577717, 32'sd173600, 32'sd254535, -32'sd160066, -32'sd1976707, -32'sd1302619, -32'sd563386, 32'sd559483, -32'sd2685417, -32'sd832573, -32'sd230592, 32'sd752422, -32'sd95558, 32'sd661168, 32'sd489502, -32'sd1765957, -32'sd2958372, -32'sd721530, -32'sd1035517, -32'sd2344537, -32'sd554491, -32'sd2067788, 32'sd1368509, 32'sd617212, -32'sd470553, 32'sd1067610, 32'sd1909482, 32'sd323283, 32'sd71024, 32'sd120191, 32'sd107262, -32'sd690657, 32'sd1065983, -32'sd33459, -32'sd1588181, -32'sd1848765, -32'sd1512183, 32'sd1596954, -32'sd1180374, 32'sd1757369, 32'sd1382778, -32'sd282741, 32'sd860231, 32'sd339767, 32'sd468686, -32'sd1434432, -32'sd50252, -32'sd921291, -32'sd501216, -32'sd873761, -32'sd196327, 32'sd218674, -32'sd341803, -32'sd111239, -32'sd168970, -32'sd42027, 32'sd48968, -32'sd170231, -32'sd1972357, -32'sd2045122, -32'sd1102420, -32'sd673878, -32'sd2214086, -32'sd2676371, 32'sd493578, 32'sd946225, 32'sd235408, 32'sd760014, -32'sd379403, 32'sd751754, 32'sd1147552, -32'sd232717, 32'sd1083393, -32'sd1939236, 32'sd595440, -32'sd1481931, -32'sd856195, -32'sd1138807, 32'sd838005, -32'sd1195367, -32'sd9538, -32'sd240379, -32'sd895615, 32'sd1628410, -32'sd595176, -32'sd835017, -32'sd2846421, -32'sd1198010, -32'sd3700014, -32'sd1911897, -32'sd2298956, 32'sd801113, 32'sd257005, 32'sd1035748, 32'sd1663715, 32'sd316273, -32'sd1604836, -32'sd767167, 32'sd1330438, 32'sd1470322, -32'sd1268899, 32'sd209322, -32'sd405861, 32'sd48111, -32'sd173776, -32'sd741837, 32'sd405148, 32'sd741490, -32'sd1233749, 32'sd1509184, -32'sd163404, 32'sd1723577, 32'sd1317110, 32'sd241948, -32'sd579506, -32'sd1144411, -32'sd1443055, -32'sd1426343, -32'sd2046177, 32'sd1018578, 32'sd1533264, 32'sd2281007, 32'sd1184315, 32'sd359694, -32'sd1735980, 32'sd162111, -32'sd221307, 32'sd278085, 32'sd1102376, 32'sd2383369, 32'sd2331076, 32'sd444747, -32'sd1236309, 32'sd1302304, 32'sd932386, 32'sd0, 32'sd654222, 32'sd506508, -32'sd416420, 32'sd1223988, 32'sd1802757, 32'sd663717, 32'sd642218, 32'sd1055852, -32'sd992435, 32'sd1378121, 32'sd205452, 32'sd161214, 32'sd2426628, 32'sd3109787, -32'sd16759, -32'sd2646920, -32'sd1853856, -32'sd543386, 32'sd1558850, 32'sd789368, 32'sd1014990, 32'sd415811, 32'sd1397821, 32'sd2136975, 32'sd1657456, -32'sd90533, -32'sd7115, -32'sd526434, 32'sd369625, 32'sd2122276, 32'sd116899, 32'sd74763, 32'sd727671, 32'sd997190, 32'sd194635, -32'sd31743, 32'sd2231987, 32'sd3055210, 32'sd2630796, -32'sd140490, 32'sd404016, 32'sd790418, -32'sd1209766, -32'sd150412, -32'sd1233840, -32'sd1233059, 32'sd930779, -32'sd418630, -32'sd1077702, 32'sd437261, -32'sd7954, 32'sd1279772, 32'sd1446000, 32'sd1115316, 32'sd790941, 32'sd764283, 32'sd297583, -32'sd682081, 32'sd1626861, -32'sd1312872, -32'sd199247, 32'sd2433084, 32'sd2027351, 32'sd1944248, 32'sd2549143, 32'sd3320855, 32'sd3335025, 32'sd1813453, 32'sd2313353, 32'sd1128296, -32'sd552952, -32'sd1002750, -32'sd1022174, -32'sd930716, -32'sd431238, -32'sd323969, -32'sd76296, 32'sd672092, 32'sd567706, 32'sd589267, -32'sd487476, 32'sd261793, 32'sd301107, 32'sd0, 32'sd646335, -32'sd1799502, 32'sd49716, -32'sd433464, 32'sd1127928, 32'sd2474588, 32'sd2057983, 32'sd3480224, 32'sd3142446, 32'sd1212078, 32'sd363088, -32'sd54125, 32'sd1728739, 32'sd3438686, -32'sd554200, -32'sd70545, -32'sd374593, -32'sd1575167, -32'sd1791777, -32'sd228001, -32'sd249155, -32'sd2447542, 32'sd892292, 32'sd1658954, 32'sd173919, 32'sd621992, -32'sd115408, 32'sd120472, 32'sd1702578, -32'sd480793, -32'sd1224120, 32'sd247988, 32'sd1583, -32'sd512958, 32'sd139786, 32'sd914024, 32'sd1222563, -32'sd176179, 32'sd690718, 32'sd58288, 32'sd1559686, -32'sd416500, -32'sd1638704, -32'sd368837, -32'sd199224, 32'sd2533005, 32'sd2069469, -32'sd344435, -32'sd699645, 32'sd390056, -32'sd1475312, -32'sd552252, 32'sd2023801, 32'sd476599, 32'sd973911, -32'sd369683, -32'sd338719, 32'sd1042065, -32'sd1880930, -32'sd276177, -32'sd431530, -32'sd466252, -32'sd726830, 32'sd1174667, 32'sd1332067, 32'sd1360443, 32'sd1213974, -32'sd1221320, -32'sd1284679, -32'sd872356, 32'sd1045909, 32'sd918267, 32'sd1006700, 32'sd2944219, 32'sd724065, -32'sd954136, -32'sd1020371, -32'sd1292591, -32'sd712022, -32'sd1297291, -32'sd1164089, 32'sd630020, 32'sd492878, 32'sd0, 32'sd1000248, -32'sd299127, 32'sd1023041, -32'sd217553, -32'sd49904, -32'sd649362, -32'sd2383024, -32'sd1838687, 32'sd399294, 32'sd1106628, 32'sd570552, -32'sd1645455, 32'sd99162, 32'sd1938539, 32'sd2069203, 32'sd2122373, 32'sd2722856, 32'sd2448731, 32'sd83204, -32'sd2503351, -32'sd298890, 32'sd753726, -32'sd887175, 32'sd936592, -32'sd1107823, -32'sd790996, 32'sd0, 32'sd0, 32'sd0, -32'sd688489, 32'sd381783, 32'sd1067896, -32'sd882856, -32'sd2838588, -32'sd1346786, -32'sd3838059, -32'sd1951592, -32'sd2531055, -32'sd128965, -32'sd1039862, 32'sd156831, 32'sd1126472, 32'sd3101228, 32'sd2734044, 32'sd2722335, 32'sd1259343, 32'sd436450, -32'sd187962, 32'sd1853248, 32'sd323924, -32'sd1808403, 32'sd856413, 32'sd1245946, 32'sd1082101, 32'sd0, 32'sd0, 32'sd0, 32'sd175314, 32'sd363502, -32'sd432716, -32'sd1090905, -32'sd2315906, -32'sd1740330, -32'sd480232, -32'sd871890, -32'sd2717642, -32'sd1654047, 32'sd456591, 32'sd509754, -32'sd447616, 32'sd1411910, 32'sd3328990, 32'sd1667540, 32'sd2794212, 32'sd3009860, 32'sd1790037, 32'sd1572073, 32'sd190811, 32'sd180737, -32'sd988757, 32'sd817641, 32'sd742930, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd416047, -32'sd622339, -32'sd1276284, -32'sd330275, -32'sd606088, -32'sd220854, -32'sd898884, -32'sd2073246, -32'sd1244342, -32'sd1247598, 32'sd382973, -32'sd2323167, -32'sd1342224, -32'sd1262901, -32'sd1015584, -32'sd297298, 32'sd595490, 32'sd1311467, 32'sd1792055, -32'sd149653, 32'sd1975174, -32'sd240159, -32'sd52711, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd337267, -32'sd55589, -32'sd341648, 32'sd135216, 32'sd609522, -32'sd49045, 32'sd867899, -32'sd1339686, -32'sd937084, -32'sd1230121, 32'sd162567, -32'sd1330714, -32'sd1479771, -32'sd300256, -32'sd596281, -32'sd1742610, 32'sd24678, -32'sd1839739, -32'sd1064777, 32'sd617177, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd181599, 32'sd1447079, 32'sd1100991, 32'sd658081, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd362603, 32'sd274249, 32'sd642032, 32'sd75951, 32'sd339181, 32'sd76351, 32'sd1141336, 32'sd155988, 32'sd498849, -32'sd1870221, 32'sd878768, -32'sd661951, 32'sd462369, 32'sd635471, -32'sd271499, -32'sd529330, -32'sd774862, 32'sd898925, 32'sd80292, 32'sd19047, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd162952, 32'sd164086, 32'sd345652, 32'sd1624216, 32'sd1374987, -32'sd1136305, -32'sd515781, 32'sd499204, 32'sd1636279, -32'sd1240762, -32'sd193944, -32'sd25458, 32'sd1696251, -32'sd1306253, -32'sd941660, 32'sd632066, 32'sd84575, -32'sd2196661, -32'sd2827548, -32'sd375856, 32'sd746526, -32'sd659945, 32'sd51101, 32'sd1759667, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd246382, -32'sd111062, -32'sd274448, 32'sd561280, 32'sd626624, -32'sd412298, 32'sd526311, 32'sd947184, 32'sd1951752, 32'sd1284813, -32'sd482561, -32'sd1547523, -32'sd660893, -32'sd818076, 32'sd194557, -32'sd515123, -32'sd1704788, -32'sd2282074, -32'sd2394511, -32'sd2558273, -32'sd2458071, -32'sd1113289, 32'sd783002, -32'sd696359, 32'sd940326, 32'sd0, 32'sd0, 32'sd470413, 32'sd1068294, 32'sd38339, 32'sd1482856, 32'sd528436, -32'sd875202, -32'sd939376, -32'sd1676149, -32'sd1302883, 32'sd316300, -32'sd306778, 32'sd280012, 32'sd2055153, 32'sd1204095, 32'sd803744, 32'sd322866, -32'sd266535, -32'sd1464000, -32'sd2127230, -32'sd653395, 32'sd19813, -32'sd574220, -32'sd2690919, -32'sd2487149, -32'sd618838, -32'sd735040, 32'sd318182, 32'sd0, 32'sd749088, 32'sd166378, -32'sd169899, 32'sd924692, -32'sd1116670, -32'sd2344878, -32'sd2263678, -32'sd1897562, -32'sd2927679, -32'sd2372296, -32'sd1005680, 32'sd5686, -32'sd779245, 32'sd2333660, 32'sd2029484, 32'sd3285262, 32'sd3606511, 32'sd1956874, 32'sd2031350, -32'sd270795, -32'sd398490, -32'sd2682834, -32'sd3923495, -32'sd1844512, 32'sd227090, -32'sd950015, 32'sd889515, 32'sd0, 32'sd212251, -32'sd601426, 32'sd634738, 32'sd1146910, -32'sd1038715, -32'sd410376, -32'sd55428, -32'sd359057, -32'sd507572, 32'sd921966, -32'sd1415143, -32'sd900550, -32'sd2660869, -32'sd1836422, 32'sd1837340, 32'sd1591828, 32'sd2497323, 32'sd2538949, 32'sd1217719, 32'sd796068, -32'sd2109338, -32'sd1945541, -32'sd1141687, -32'sd1091238, 32'sd1328762, -32'sd694510, -32'sd321772, 32'sd1292054, -32'sd245745, -32'sd2288231, 32'sd2522510, 32'sd1781926, 32'sd77683, 32'sd660089, -32'sd873130, -32'sd273581, 32'sd363306, 32'sd1305299, -32'sd571350, -32'sd772238, -32'sd2971586, -32'sd2839090, -32'sd223837, 32'sd171353, 32'sd2820888, 32'sd1548945, 32'sd1195520, 32'sd272888, -32'sd2180824, 32'sd322262, -32'sd3607451, -32'sd173845, 32'sd1261325, -32'sd589522, 32'sd646589, -32'sd13975, -32'sd255169, -32'sd138174, -32'sd628993, -32'sd1745187, -32'sd868963, -32'sd333798, -32'sd1012952, -32'sd1550956, -32'sd1599471, 32'sd545741, -32'sd1905327, -32'sd2223788, -32'sd1617928, -32'sd228390, -32'sd519549, 32'sd2168782, 32'sd857341, 32'sd2231407, 32'sd1703940, 32'sd237870, -32'sd387551, -32'sd1273376, 32'sd988746, -32'sd1328749, -32'sd2586791, -32'sd1348618, 32'sd603414, 32'sd803265, -32'sd1428676, 32'sd1010326, -32'sd1294831, -32'sd81038, -32'sd2668544, -32'sd2208067, -32'sd1939847, -32'sd2086240, -32'sd1391562, -32'sd1017079, -32'sd24728, 32'sd41355, 32'sd145835, -32'sd755776, 32'sd2303269, 32'sd1808396, 32'sd790885, 32'sd1580919, 32'sd1243549, -32'sd37349, -32'sd1332200, 32'sd405907, 32'sd1074395, 32'sd855370, -32'sd1435306, -32'sd546641, -32'sd314517, -32'sd367439, 32'sd276641, -32'sd1679518, -32'sd627066, 32'sd1017727, -32'sd1385541, -32'sd785319, -32'sd537227, -32'sd421137, -32'sd2794368, -32'sd1404865, -32'sd520253, -32'sd397369, -32'sd605009, -32'sd1031329, 32'sd918819, 32'sd2551540, 32'sd135580, 32'sd1356249, 32'sd2292335, -32'sd771480, -32'sd878072, -32'sd145039, -32'sd885065, 32'sd400752, -32'sd2939693, -32'sd640812, 32'sd714027, -32'sd226301, -32'sd2770539, 32'sd580053, 32'sd195967, 32'sd750787, -32'sd587585, -32'sd1592260, -32'sd2973164, -32'sd2478600, -32'sd1572071, -32'sd493374, -32'sd740527, 32'sd984203, -32'sd378964, 32'sd228402, -32'sd667253, 32'sd1241764, -32'sd2209555, 32'sd602790, 32'sd1098167, -32'sd1008909, -32'sd1297649, -32'sd1432296, -32'sd469369, 32'sd80212, -32'sd226162, -32'sd401343, -32'sd2378000, 32'sd1366155, 32'sd103050, 32'sd851308, 32'sd1032961, -32'sd389657, -32'sd981250, -32'sd554085, -32'sd2008477, -32'sd1321543, -32'sd1097797, 32'sd1503775, -32'sd1471642, -32'sd5214, 32'sd199832, -32'sd2343296, -32'sd555467, 32'sd137544, -32'sd580894, -32'sd3019752, -32'sd309991, -32'sd1322836, -32'sd2536999, -32'sd2286017, -32'sd172440, -32'sd616003, 32'sd567441, 32'sd633656, -32'sd507723, 32'sd585986, 32'sd159090, 32'sd2481, 32'sd1500510, 32'sd936980, -32'sd1212474, 32'sd419515, -32'sd1208723, 32'sd435869, 32'sd1506929, 32'sd105990, 32'sd629354, 32'sd1635755, -32'sd117610, -32'sd2032750, -32'sd1280635, -32'sd1112733, -32'sd176447, -32'sd380196, -32'sd2432338, -32'sd234945, -32'sd1015518, -32'sd453735, -32'sd1395089, -32'sd773631, 32'sd1064210, 32'sd250579, -32'sd354178, -32'sd178236, -32'sd1669790, -32'sd1333647, -32'sd431944, -32'sd1458781, -32'sd1791204, -32'sd285184, 32'sd2560556, 32'sd903122, 32'sd420042, 32'sd349407, 32'sd1245387, 32'sd519533, -32'sd157176, -32'sd534234, -32'sd1659265, -32'sd455257, 32'sd1027939, -32'sd2632100, -32'sd1199651, -32'sd718781, 32'sd990645, -32'sd2144636, -32'sd539253, 32'sd561769, 32'sd37596, 32'sd879495, 32'sd210934, 32'sd45344, 32'sd10111, -32'sd306748, 32'sd103151, -32'sd1096010, 32'sd1782261, 32'sd2598241, 32'sd3564835, 32'sd3153689, 32'sd2751247, 32'sd206556, -32'sd193804, 32'sd1153969, 32'sd434446, -32'sd275039, 32'sd675446, 32'sd488126, -32'sd289686, -32'sd1343864, 32'sd559442, -32'sd632811, -32'sd1358009, 32'sd1433861, 32'sd1046001, 32'sd1004125, 32'sd2215003, -32'sd467269, -32'sd1236997, 32'sd848069, -32'sd560529, -32'sd1548710, 32'sd846190, -32'sd619941, 32'sd957321, 32'sd1063037, 32'sd2375035, 32'sd2608472, 32'sd2542054, -32'sd2034205, -32'sd2395418, -32'sd1203794, -32'sd249313, -32'sd1796813, -32'sd62586, 32'sd1971254, 32'sd2273286, -32'sd1668460, -32'sd1903907, -32'sd1431852, 32'sd1050610, 32'sd2462429, 32'sd1101479, -32'sd991952, 32'sd290037, 32'sd1803259, 32'sd81658, 32'sd0, 32'sd984267, 32'sd534094, -32'sd872582, 32'sd653694, 32'sd1848019, 32'sd1275855, 32'sd1219636, 32'sd1872269, 32'sd1275182, 32'sd563966, -32'sd809132, 32'sd482691, -32'sd653623, 32'sd370230, 32'sd1798143, 32'sd1063884, -32'sd387385, -32'sd1741142, -32'sd1576108, -32'sd1097136, -32'sd716444, 32'sd1474103, -32'sd645810, -32'sd1209854, 32'sd881712, -32'sd1361520, 32'sd1066158, 32'sd515103, 32'sd487758, -32'sd416398, 32'sd479714, 32'sd1743391, 32'sd1099731, 32'sd2054313, 32'sd1810147, 32'sd582128, -32'sd147674, 32'sd130792, -32'sd830312, 32'sd74847, 32'sd948005, 32'sd307057, -32'sd129038, 32'sd1346388, 32'sd220314, 32'sd1157408, 32'sd1485981, 32'sd2150542, -32'sd373419, 32'sd1238594, 32'sd38167, -32'sd505574, 32'sd839269, 32'sd988133, -32'sd163031, 32'sd504231, 32'sd534398, -32'sd649273, 32'sd411669, -32'sd483206, 32'sd514492, 32'sd1598253, 32'sd2223532, 32'sd131559, -32'sd65018, -32'sd471645, -32'sd2066002, -32'sd1358588, -32'sd596706, 32'sd325100, -32'sd2807142, 32'sd2265178, 32'sd1240575, 32'sd1187501, 32'sd2810178, 32'sd350044, -32'sd24832, 32'sd1790706, 32'sd220043, -32'sd757732, -32'sd61849, 32'sd655956, 32'sd1508841, 32'sd0, 32'sd79664, 32'sd1235432, 32'sd1570939, 32'sd1108473, 32'sd2386209, 32'sd2623400, 32'sd1195339, -32'sd1053801, -32'sd2370927, -32'sd3270110, -32'sd3558316, -32'sd2285694, -32'sd1362721, -32'sd4295862, -32'sd3620498, -32'sd297715, 32'sd2040358, 32'sd1086152, 32'sd2229850, -32'sd238738, 32'sd1293262, 32'sd798775, 32'sd1442838, -32'sd221380, 32'sd1706791, -32'sd383276, 32'sd281348, 32'sd614955, -32'sd1556945, -32'sd592971, 32'sd209146, 32'sd1655443, 32'sd1594692, 32'sd963301, 32'sd1240321, 32'sd2138562, -32'sd255113, -32'sd188551, -32'sd1995774, -32'sd3662761, -32'sd3556141, -32'sd2605037, -32'sd2875529, -32'sd761788, 32'sd933271, 32'sd626977, 32'sd2855639, 32'sd1079562, -32'sd1329106, 32'sd754188, -32'sd320248, -32'sd806023, 32'sd434775, 32'sd537526, -32'sd570257, 32'sd124978, 32'sd6710, 32'sd644399, 32'sd695347, 32'sd125048, -32'sd1492234, -32'sd286149, -32'sd553784, 32'sd2373612, 32'sd417157, 32'sd160625, -32'sd1715324, -32'sd3141317, -32'sd3193814, -32'sd1808584, -32'sd2686734, 32'sd1362849, 32'sd1171068, 32'sd775427, -32'sd480475, -32'sd1119577, -32'sd1188124, 32'sd1068460, -32'sd2871132, -32'sd796277, 32'sd1098009, 32'sd45349, 32'sd314455, 32'sd0, 32'sd528373, 32'sd1212473, 32'sd33800, 32'sd608010, -32'sd2511321, -32'sd2520027, 32'sd947654, 32'sd1153726, 32'sd1108331, -32'sd280219, -32'sd449459, -32'sd2013034, 32'sd643560, -32'sd930199, -32'sd101417, 32'sd658928, -32'sd2445268, 32'sd757797, -32'sd193071, -32'sd865166, -32'sd2071167, -32'sd667125, -32'sd744739, -32'sd1127275, -32'sd1325788, 32'sd120189, 32'sd0, 32'sd0, 32'sd0, -32'sd789192, -32'sd1680305, -32'sd708403, -32'sd722264, -32'sd1417233, -32'sd2298401, -32'sd1079720, 32'sd1358744, 32'sd350865, 32'sd54663, -32'sd1440291, -32'sd53729, -32'sd1661314, -32'sd2151760, -32'sd507044, 32'sd200548, 32'sd1541024, -32'sd1040446, -32'sd25302, 32'sd805995, -32'sd902243, -32'sd1137543, -32'sd1755282, -32'sd268514, 32'sd1352297, 32'sd0, 32'sd0, 32'sd0, 32'sd621878, 32'sd350234, 32'sd51832, -32'sd1168205, -32'sd36258, -32'sd632992, 32'sd980267, -32'sd580907, -32'sd4157113, -32'sd4018289, -32'sd3783216, -32'sd2819625, -32'sd2677319, -32'sd1165143, -32'sd1332890, -32'sd2260055, -32'sd718124, -32'sd2762476, -32'sd1933281, 32'sd818075, 32'sd126644, 32'sd387701, 32'sd368866, 32'sd838334, 32'sd67463, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd920699, -32'sd74337, -32'sd231896, -32'sd827392, 32'sd129453, 32'sd956220, -32'sd299195, -32'sd1361558, 32'sd495171, -32'sd496327, 32'sd242393, -32'sd457935, -32'sd1302189, -32'sd271231, -32'sd539681, -32'sd2470562, -32'sd310423, 32'sd125720, 32'sd134837, 32'sd671315, -32'sd258173, 32'sd619948, 32'sd393146, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd130657, 32'sd698077, 32'sd160868, 32'sd1042444, -32'sd809583, -32'sd239441, 32'sd480575, -32'sd166782, 32'sd324378, -32'sd1133401, 32'sd1133279, -32'sd1214893, -32'sd90699, -32'sd1249208, 32'sd732645, 32'sd251218, -32'sd514358, 32'sd1062092, 32'sd2129330, 32'sd540680, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd281528, -32'sd1220395, 32'sd770669, 32'sd576497, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1710779, -32'sd329847, 32'sd1513091, 32'sd1435254, 32'sd192055, -32'sd10151, 32'sd428571, 32'sd968256, 32'sd464316, -32'sd42050, 32'sd257811, -32'sd858689, -32'sd1448198, -32'sd104124, 32'sd1132121, 32'sd1058078, 32'sd80882, 32'sd1186488, -32'sd1103123, 32'sd964767, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1073561, 32'sd781502, 32'sd1232848, 32'sd576576, 32'sd211309, 32'sd1099010, 32'sd1371474, 32'sd1083324, -32'sd498820, 32'sd13636, 32'sd417584, 32'sd2326149, 32'sd1185461, -32'sd565890, -32'sd103256, -32'sd952301, -32'sd1603083, -32'sd57318, 32'sd774906, -32'sd571141, 32'sd1284814, -32'sd125260, 32'sd250045, 32'sd410799, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd806779, 32'sd1316470, -32'sd221083, 32'sd955935, 32'sd1605473, 32'sd1135944, -32'sd588436, 32'sd126541, 32'sd107351, -32'sd1491407, -32'sd1310730, -32'sd1333553, -32'sd801785, -32'sd2123739, -32'sd2731768, -32'sd1135885, -32'sd2819621, 32'sd2511385, 32'sd2762061, 32'sd993760, 32'sd2060913, 32'sd50801, 32'sd919160, -32'sd1825907, 32'sd873463, 32'sd0, 32'sd0, 32'sd1217178, 32'sd813913, -32'sd386596, 32'sd475372, 32'sd744268, 32'sd390279, 32'sd362830, 32'sd1442434, 32'sd1616770, -32'sd1327614, -32'sd1044646, -32'sd1444912, 32'sd1963942, -32'sd896734, 32'sd815416, 32'sd2273721, 32'sd1413168, -32'sd40673, 32'sd1441763, 32'sd2093798, 32'sd2953066, 32'sd1019060, 32'sd46129, -32'sd568590, 32'sd462543, 32'sd248919, 32'sd468845, 32'sd0, 32'sd784429, -32'sd1251715, 32'sd970484, 32'sd318081, 32'sd113973, -32'sd110551, 32'sd318182, 32'sd1580585, 32'sd3296395, 32'sd2662419, -32'sd2412387, -32'sd2749655, -32'sd1528824, -32'sd2221397, -32'sd260611, -32'sd589025, 32'sd218424, 32'sd52815, 32'sd267694, 32'sd1446158, -32'sd960794, -32'sd877429, -32'sd100747, -32'sd249008, 32'sd954816, 32'sd1107806, 32'sd741508, 32'sd0, 32'sd418650, -32'sd280681, 32'sd582264, 32'sd2111324, 32'sd1235077, 32'sd1479261, -32'sd1189421, 32'sd746863, -32'sd8767, -32'sd1257342, -32'sd1866675, -32'sd2506590, -32'sd1684559, -32'sd1456978, -32'sd1191734, -32'sd2259891, 32'sd230804, -32'sd1234636, -32'sd605901, 32'sd503157, 32'sd1300001, 32'sd1397618, 32'sd1240667, -32'sd298297, -32'sd56421, -32'sd615165, 32'sd515480, 32'sd560026, 32'sd682648, 32'sd1154461, -32'sd501866, -32'sd380120, 32'sd252645, 32'sd919724, 32'sd1610606, 32'sd2812, -32'sd763747, 32'sd1698024, -32'sd696641, -32'sd843069, -32'sd2616473, -32'sd1792379, -32'sd2139670, -32'sd1415634, -32'sd1429319, -32'sd606198, 32'sd948141, -32'sd319016, 32'sd1611057, -32'sd136754, 32'sd892702, 32'sd335811, 32'sd1150470, 32'sd1298888, 32'sd1148707, 32'sd123150, -32'sd625775, 32'sd158888, 32'sd1216362, -32'sd186097, 32'sd974301, 32'sd1071722, 32'sd840948, -32'sd585791, 32'sd2587761, 32'sd753298, 32'sd1819216, 32'sd146163, -32'sd2634350, -32'sd2470690, -32'sd1208102, 32'sd880572, 32'sd541064, 32'sd606574, -32'sd465367, 32'sd1116630, 32'sd2247519, 32'sd286987, 32'sd542136, 32'sd1962604, 32'sd803060, 32'sd1531835, -32'sd1375225, 32'sd543832, 32'sd782217, 32'sd813821, -32'sd969859, 32'sd1954105, -32'sd653837, 32'sd915962, -32'sd215296, 32'sd1817734, 32'sd991208, 32'sd1132979, 32'sd825041, 32'sd634012, -32'sd1476564, -32'sd3602392, -32'sd829405, 32'sd1224400, 32'sd632147, -32'sd1337188, -32'sd535322, 32'sd1291240, 32'sd1832104, 32'sd47086, 32'sd1334318, 32'sd376412, 32'sd957780, -32'sd584120, 32'sd466432, 32'sd1436680, 32'sd952753, 32'sd645532, 32'sd1313165, 32'sd68899, -32'sd309688, -32'sd554788, 32'sd350258, 32'sd1057917, 32'sd2161535, 32'sd1340683, 32'sd1624057, 32'sd103396, -32'sd1218667, -32'sd3509963, 32'sd446434, -32'sd1908961, -32'sd439071, -32'sd740185, 32'sd204309, -32'sd1669385, -32'sd381943, 32'sd354366, -32'sd1732882, -32'sd795031, 32'sd467676, 32'sd709443, 32'sd417070, 32'sd1053959, -32'sd214828, 32'sd1115744, 32'sd479366, -32'sd1922508, 32'sd685879, 32'sd2143542, 32'sd1337452, 32'sd1730214, 32'sd2710900, 32'sd1595089, 32'sd1075830, 32'sd1712453, -32'sd4133014, -32'sd4301682, -32'sd231166, -32'sd1078881, 32'sd318063, -32'sd1098508, -32'sd2203598, -32'sd812813, -32'sd1213307, -32'sd1028697, -32'sd1002485, -32'sd1645540, 32'sd933765, -32'sd83037, -32'sd240638, -32'sd155167, -32'sd1240414, 32'sd1035490, 32'sd234777, 32'sd54718, 32'sd758649, 32'sd597960, 32'sd1777531, 32'sd1803629, 32'sd431868, 32'sd3611439, 32'sd2870868, -32'sd1148817, -32'sd2674801, -32'sd2053578, -32'sd1832556, 32'sd445812, -32'sd1308530, -32'sd428569, -32'sd65966, -32'sd842179, -32'sd2318508, -32'sd317434, -32'sd564248, -32'sd2031952, -32'sd1962715, -32'sd2460719, -32'sd610815, 32'sd848816, -32'sd1369878, -32'sd305400, -32'sd1437492, -32'sd482092, 32'sd1389610, 32'sd2193420, 32'sd3259996, 32'sd611065, -32'sd190336, 32'sd2804322, 32'sd88205, -32'sd1550037, -32'sd3503261, -32'sd2541353, -32'sd601878, 32'sd124171, 32'sd192414, -32'sd875403, 32'sd1369880, -32'sd925220, -32'sd130769, -32'sd1074130, -32'sd1155618, -32'sd1442945, 32'sd962956, -32'sd766974, -32'sd168111, 32'sd2360510, 32'sd173292, 32'sd460910, -32'sd998831, 32'sd731422, 32'sd1509199, 32'sd96462, -32'sd118207, 32'sd571423, 32'sd1025050, 32'sd2415100, 32'sd484839, -32'sd1162717, -32'sd2492515, -32'sd1670635, -32'sd1000351, 32'sd831870, 32'sd38809, 32'sd562394, 32'sd1338294, 32'sd269144, -32'sd401879, 32'sd1886865, -32'sd370576, -32'sd318441, -32'sd2196172, 32'sd237426, 32'sd712593, -32'sd425801, 32'sd140296, 32'sd1049571, -32'sd673118, 32'sd882106, -32'sd1612247, 32'sd459434, 32'sd302376, 32'sd1016846, 32'sd625030, 32'sd2213888, 32'sd669064, -32'sd1807457, -32'sd2596487, -32'sd2596175, 32'sd1664167, 32'sd288461, -32'sd86336, 32'sd1727496, 32'sd2133037, -32'sd363105, -32'sd605709, 32'sd2549750, 32'sd11637, -32'sd2162397, -32'sd1169572, -32'sd1468437, 32'sd1013640, 32'sd508896, 32'sd516762, 32'sd388912, 32'sd618856, 32'sd1288996, -32'sd325785, 32'sd1786529, 32'sd813423, 32'sd2283623, 32'sd1661186, 32'sd426188, -32'sd1156562, -32'sd304566, -32'sd4126598, -32'sd2978960, 32'sd677614, -32'sd727085, 32'sd1237402, 32'sd486362, 32'sd950968, 32'sd2091765, -32'sd368938, -32'sd519530, 32'sd489400, -32'sd76762, -32'sd1489442, -32'sd2677450, -32'sd873255, 32'sd0, 32'sd1054455, -32'sd612315, 32'sd702913, -32'sd127298, -32'sd148712, 32'sd1163650, 32'sd1782205, 32'sd1947686, -32'sd326495, 32'sd1400416, -32'sd1159077, -32'sd3801553, -32'sd4209905, -32'sd1427601, 32'sd1321302, 32'sd1924178, 32'sd1413583, 32'sd2306816, -32'sd658098, 32'sd649686, 32'sd724845, -32'sd1187057, -32'sd2274660, -32'sd417235, 32'sd644845, -32'sd287317, 32'sd730063, 32'sd158426, -32'sd1135248, 32'sd1994477, -32'sd398842, -32'sd272837, -32'sd237385, -32'sd544978, -32'sd944614, -32'sd3196755, -32'sd1000580, -32'sd2550207, -32'sd2214495, -32'sd2760967, -32'sd1284232, 32'sd273789, 32'sd2152411, 32'sd2012238, 32'sd1919321, -32'sd176767, -32'sd939768, 32'sd2111581, 32'sd1222582, 32'sd639340, -32'sd1791235, 32'sd1350497, -32'sd1807762, 32'sd1553679, 32'sd382703, 32'sd965404, 32'sd371047, -32'sd1175912, 32'sd1589644, -32'sd559554, 32'sd198758, 32'sd242623, -32'sd3616960, -32'sd2207848, -32'sd1240267, -32'sd3313537, -32'sd3441481, -32'sd3979628, -32'sd1207623, 32'sd22621, 32'sd2596930, 32'sd259951, -32'sd537256, 32'sd841501, -32'sd519550, -32'sd1318627, -32'sd1373574, -32'sd1596461, 32'sd120659, -32'sd726358, -32'sd2108535, -32'sd482702, 32'sd603681, 32'sd0, 32'sd161911, 32'sd697101, 32'sd753978, -32'sd1895044, -32'sd1599246, 32'sd689390, -32'sd1128620, -32'sd1121460, -32'sd3091396, -32'sd2408118, -32'sd1565821, -32'sd1989764, -32'sd790662, -32'sd344908, 32'sd638226, 32'sd889094, 32'sd1869143, 32'sd308911, -32'sd650720, -32'sd56990, 32'sd561753, 32'sd640103, 32'sd1401111, -32'sd1445875, -32'sd1691295, 32'sd1253423, 32'sd1229763, 32'sd1490203, 32'sd674172, 32'sd748443, 32'sd744949, -32'sd363515, -32'sd1756836, -32'sd1829411, -32'sd2082047, -32'sd1381917, -32'sd1819784, -32'sd2465557, -32'sd2821398, 32'sd461076, 32'sd1924068, -32'sd1343775, 32'sd792377, -32'sd819847, 32'sd941997, 32'sd940321, 32'sd1486000, -32'sd317636, 32'sd184522, 32'sd1680609, -32'sd172646, -32'sd459695, 32'sd860982, -32'sd40931, -32'sd885478, 32'sd2699271, 32'sd822478, -32'sd31331, -32'sd1652678, 32'sd109303, -32'sd1485278, 32'sd542642, -32'sd376257, -32'sd41129, -32'sd1078726, -32'sd1151896, -32'sd2376646, -32'sd1034934, 32'sd849761, 32'sd271430, 32'sd898600, 32'sd482534, -32'sd111912, 32'sd1692790, 32'sd2161667, -32'sd92618, 32'sd2554888, -32'sd1444034, 32'sd1138335, 32'sd160924, 32'sd114699, -32'sd311653, 32'sd824220, 32'sd0, 32'sd1681567, 32'sd899186, -32'sd132421, 32'sd596108, 32'sd1777577, 32'sd979606, 32'sd132415, -32'sd75785, -32'sd523639, 32'sd789588, 32'sd837648, 32'sd904333, 32'sd303338, 32'sd608833, -32'sd850913, 32'sd1955441, 32'sd523115, 32'sd374359, -32'sd552012, 32'sd969533, -32'sd131438, -32'sd669711, 32'sd628950, 32'sd534115, 32'sd42263, 32'sd761209, 32'sd0, 32'sd0, 32'sd0, -32'sd621959, 32'sd1148748, -32'sd264218, 32'sd2024371, 32'sd1326902, 32'sd349485, 32'sd459597, -32'sd811276, -32'sd2649960, 32'sd1185288, 32'sd897974, 32'sd626417, 32'sd1121557, -32'sd582336, 32'sd1563379, 32'sd1822606, 32'sd623735, 32'sd1012567, 32'sd636747, 32'sd1198164, 32'sd594620, 32'sd196741, 32'sd1823704, 32'sd1124500, -32'sd414166, 32'sd0, 32'sd0, 32'sd0, 32'sd340650, 32'sd577809, -32'sd138631, 32'sd576180, 32'sd446892, -32'sd2008542, -32'sd807518, 32'sd565231, -32'sd1467002, 32'sd1926091, 32'sd2197997, -32'sd321149, 32'sd715482, 32'sd506160, 32'sd488680, 32'sd416241, 32'sd385191, -32'sd1000317, 32'sd759538, 32'sd1116643, 32'sd1209364, 32'sd1465393, -32'sd140505, -32'sd1189528, 32'sd423, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1255915, 32'sd772092, 32'sd480998, -32'sd1484516, -32'sd1275634, -32'sd885245, -32'sd123790, -32'sd684519, -32'sd732168, -32'sd359278, -32'sd898454, -32'sd1307755, 32'sd1192872, 32'sd915129, -32'sd179413, -32'sd856060, -32'sd788645, -32'sd997363, -32'sd1136815, 32'sd906975, 32'sd776541, -32'sd265703, 32'sd1112725, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1384110, 32'sd427725, 32'sd18716, 32'sd1014629, 32'sd380760, 32'sd910379, 32'sd370508, 32'sd355858, 32'sd1262676, -32'sd1360820, -32'sd820106, -32'sd1783189, -32'sd240484, 32'sd1576358, -32'sd876480, 32'sd463206, -32'sd1864000, 32'sd604061, 32'sd1653678, 32'sd2004540, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd158338, -32'sd586926, -32'sd211020, 32'sd672578, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd254175, -32'sd338550, 32'sd41841, -32'sd399009, 32'sd183305, -32'sd1402159, 32'sd254212, 32'sd570318, -32'sd600807, -32'sd676392, -32'sd1072689, -32'sd488176, -32'sd180217, 32'sd462991, -32'sd778315, 32'sd504378, 32'sd33602, 32'sd639640, -32'sd1214252, 32'sd687462, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd556657, 32'sd331903, -32'sd506405, -32'sd159710, 32'sd199044, -32'sd1597344, -32'sd594715, -32'sd2176957, 32'sd537389, -32'sd241900, -32'sd929139, 32'sd919660, -32'sd1448737, 32'sd921935, 32'sd422402, 32'sd1184667, 32'sd1741432, -32'sd181772, 32'sd255939, 32'sd1127152, 32'sd1064645, 32'sd277743, 32'sd1067883, -32'sd201667, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd150976, -32'sd74447, 32'sd993707, -32'sd352591, -32'sd749257, -32'sd46502, 32'sd2626789, -32'sd1763381, 32'sd1500145, -32'sd1992312, -32'sd1956399, -32'sd589874, -32'sd2188431, -32'sd510971, -32'sd177312, -32'sd1775905, -32'sd2283689, -32'sd2035950, -32'sd651123, -32'sd527151, 32'sd258847, 32'sd87304, 32'sd428310, -32'sd496423, -32'sd174428, 32'sd0, 32'sd0, -32'sd275787, 32'sd511871, -32'sd419015, 32'sd460278, 32'sd445117, 32'sd348460, 32'sd738607, 32'sd59719, -32'sd328790, 32'sd2165939, 32'sd1108630, 32'sd1339472, 32'sd1561645, -32'sd788928, 32'sd16144, -32'sd477954, -32'sd239370, 32'sd1773289, 32'sd735960, -32'sd2600011, 32'sd537526, 32'sd420761, -32'sd723473, 32'sd1748473, -32'sd751258, 32'sd294106, 32'sd577367, 32'sd0, 32'sd1071684, 32'sd592974, 32'sd1583035, -32'sd1379022, -32'sd337630, -32'sd532838, -32'sd190645, 32'sd732949, 32'sd713913, 32'sd1013301, 32'sd1797904, 32'sd378543, 32'sd165761, -32'sd2114061, -32'sd1667328, -32'sd683010, 32'sd879619, 32'sd723669, 32'sd1191759, 32'sd941256, 32'sd1087825, -32'sd1915038, -32'sd1465361, 32'sd682514, 32'sd235154, -32'sd341607, -32'sd198444, 32'sd0, -32'sd197596, 32'sd34325, 32'sd709774, -32'sd1054312, 32'sd951753, 32'sd466014, -32'sd1040506, 32'sd659178, 32'sd937441, 32'sd211851, 32'sd2330609, 32'sd553148, 32'sd288484, 32'sd1814973, 32'sd1404993, -32'sd574977, -32'sd27916, 32'sd1097837, -32'sd1331313, -32'sd1329651, 32'sd995757, -32'sd1864615, 32'sd773508, 32'sd807406, -32'sd1695564, -32'sd1527, -32'sd979523, 32'sd110621, -32'sd864332, 32'sd59845, -32'sd575337, -32'sd47264, 32'sd808787, 32'sd25041, 32'sd642323, 32'sd1911651, 32'sd733305, -32'sd527320, 32'sd883465, 32'sd939536, 32'sd2739510, 32'sd544773, 32'sd1319399, 32'sd1555645, -32'sd1434501, 32'sd535210, -32'sd1292264, 32'sd903159, 32'sd1184152, -32'sd1195231, -32'sd3353918, -32'sd1016457, -32'sd1156796, -32'sd966374, -32'sd307848, 32'sd722144, -32'sd857809, -32'sd1338454, 32'sd338663, -32'sd260220, 32'sd372573, -32'sd647786, 32'sd862650, 32'sd2623095, 32'sd2197441, 32'sd1082324, -32'sd771693, 32'sd1863078, 32'sd1082865, 32'sd1202117, -32'sd1082410, -32'sd1398312, 32'sd185290, -32'sd1005407, -32'sd946193, -32'sd796827, -32'sd2154279, -32'sd2080036, 32'sd228164, -32'sd1039152, -32'sd938228, 32'sd621473, -32'sd128856, 32'sd325779, 32'sd37857, 32'sd1293824, -32'sd1127516, 32'sd93141, 32'sd1112564, 32'sd1013135, 32'sd397690, 32'sd2136188, -32'sd445175, -32'sd1533654, -32'sd354286, -32'sd53954, 32'sd763781, -32'sd444138, 32'sd1091290, 32'sd1058494, -32'sd1419170, -32'sd1415238, -32'sd924998, 32'sd553196, -32'sd1474020, -32'sd2037497, -32'sd248803, 32'sd919467, 32'sd15877, -32'sd1174426, 32'sd1232505, -32'sd324792, 32'sd151489, -32'sd803643, 32'sd1866366, 32'sd65786, 32'sd2257900, 32'sd705051, 32'sd3171933, 32'sd278449, -32'sd1310043, -32'sd2237751, -32'sd2716966, -32'sd2651280, 32'sd296211, 32'sd741966, 32'sd1222656, -32'sd477014, 32'sd665746, 32'sd215539, -32'sd1382055, 32'sd1147103, 32'sd157571, -32'sd17836, -32'sd73002, -32'sd2232010, 32'sd780011, 32'sd37139, -32'sd536524, 32'sd729499, -32'sd1292549, -32'sd1211003, 32'sd941785, 32'sd512428, 32'sd138213, -32'sd996088, 32'sd2084248, 32'sd209053, -32'sd2890900, -32'sd1572779, 32'sd1361197, 32'sd990218, 32'sd241536, 32'sd1252184, 32'sd568968, 32'sd956416, 32'sd1095388, 32'sd1351976, -32'sd1306859, 32'sd140911, -32'sd1632787, -32'sd1031747, -32'sd2276634, 32'sd76657, 32'sd664749, -32'sd289498, 32'sd170023, -32'sd191645, 32'sd681170, -32'sd406062, 32'sd210684, -32'sd390855, 32'sd392939, 32'sd1383152, -32'sd1652731, 32'sd261199, 32'sd365280, 32'sd191745, 32'sd1891940, 32'sd100496, 32'sd1932680, 32'sd3272110, 32'sd735939, 32'sd805591, 32'sd955931, 32'sd740902, -32'sd973305, -32'sd1125268, -32'sd1363595, -32'sd3112671, -32'sd916080, -32'sd443989, -32'sd62390, -32'sd524221, 32'sd856283, 32'sd355476, -32'sd520961, -32'sd1609168, 32'sd68582, -32'sd2065184, -32'sd421640, 32'sd766961, -32'sd791265, 32'sd714611, -32'sd900413, -32'sd630153, 32'sd1239800, 32'sd1771784, 32'sd2132267, 32'sd1767281, -32'sd1489020, -32'sd893993, 32'sd1231956, 32'sd126487, -32'sd625652, -32'sd858294, -32'sd989436, -32'sd1355502, -32'sd509510, 32'sd919807, -32'sd1227399, -32'sd412826, -32'sd475513, 32'sd320503, -32'sd14225, -32'sd925684, -32'sd1789978, -32'sd2112849, -32'sd234112, -32'sd1030989, 32'sd624727, 32'sd633963, 32'sd236467, -32'sd1821057, -32'sd442357, 32'sd641309, 32'sd1700253, 32'sd2131324, -32'sd443921, -32'sd1163789, -32'sd729048, 32'sd577207, 32'sd51747, -32'sd48297, -32'sd1625241, -32'sd1365104, -32'sd779734, 32'sd21084, -32'sd1136272, -32'sd1553122, 32'sd771703, -32'sd34310, -32'sd423359, -32'sd815733, -32'sd1186090, -32'sd1014854, -32'sd1721190, 32'sd227332, -32'sd1446667, 32'sd1503291, 32'sd390799, -32'sd282222, 32'sd885258, 32'sd1083672, 32'sd135685, 32'sd2198535, 32'sd1716632, 32'sd1435659, 32'sd1265193, -32'sd757752, 32'sd1458644, 32'sd438851, -32'sd629713, 32'sd463508, 32'sd1071954, 32'sd1694499, 32'sd1917208, 32'sd681744, 32'sd326407, -32'sd549012, -32'sd694858, -32'sd1262694, -32'sd1220560, -32'sd1177001, -32'sd876773, -32'sd191808, 32'sd85747, -32'sd2502854, -32'sd1683106, -32'sd1872232, -32'sd780172, -32'sd949054, 32'sd924469, 32'sd1603686, -32'sd857125, 32'sd271663, -32'sd507370, 32'sd1641937, 32'sd914051, 32'sd1859710, 32'sd768647, 32'sd1448851, 32'sd276916, 32'sd2150159, 32'sd1873043, 32'sd234825, 32'sd23638, 32'sd0, -32'sd690109, 32'sd400154, -32'sd941964, -32'sd560996, -32'sd994787, 32'sd79444, 32'sd1039214, -32'sd332610, -32'sd2416238, -32'sd3370222, -32'sd3688620, -32'sd3247443, -32'sd1946084, -32'sd2279215, -32'sd2343471, -32'sd1082997, -32'sd1276350, 32'sd2014097, 32'sd3573505, 32'sd2000363, 32'sd1172355, 32'sd1970273, 32'sd1191882, 32'sd527930, -32'sd1829091, 32'sd715364, 32'sd1769417, -32'sd242826, 32'sd176918, 32'sd663769, 32'sd1181460, -32'sd1274099, -32'sd306389, -32'sd1370654, -32'sd326807, -32'sd733903, -32'sd1583079, -32'sd4170858, -32'sd4566490, -32'sd3536619, -32'sd3332371, -32'sd3281537, -32'sd3040903, -32'sd1543343, 32'sd209447, 32'sd2146568, 32'sd2971809, 32'sd2525875, 32'sd3224338, -32'sd361433, -32'sd826118, -32'sd1748245, -32'sd996234, 32'sd2169363, 32'sd1469947, -32'sd88598, -32'sd825498, -32'sd674991, 32'sd1289800, -32'sd1411164, 32'sd832089, 32'sd474693, -32'sd561854, -32'sd1483770, -32'sd277343, 32'sd458611, -32'sd403628, -32'sd1041671, -32'sd2265564, -32'sd2882421, -32'sd3006947, -32'sd1386046, -32'sd1914375, 32'sd1231860, 32'sd1302339, 32'sd2333141, 32'sd2942459, 32'sd1481507, -32'sd357383, -32'sd1181286, 32'sd819880, 32'sd1608977, 32'sd1343767, 32'sd0, 32'sd498825, 32'sd147195, 32'sd595792, -32'sd248080, -32'sd922825, -32'sd309736, -32'sd514579, -32'sd487365, -32'sd448369, 32'sd332195, -32'sd499053, 32'sd74033, -32'sd1992484, -32'sd2771217, -32'sd2273079, 32'sd252903, -32'sd1187999, 32'sd1721158, 32'sd2476147, 32'sd2133678, 32'sd2252693, 32'sd2037917, 32'sd1110919, -32'sd420255, -32'sd966581, 32'sd1037497, 32'sd18270, 32'sd70474, -32'sd406082, 32'sd1976436, -32'sd1034588, 32'sd165701, -32'sd589270, -32'sd567241, 32'sd941744, -32'sd585258, -32'sd28400, 32'sd1201694, 32'sd828192, 32'sd1180917, 32'sd1078573, 32'sd347332, -32'sd105438, 32'sd1743723, 32'sd177900, -32'sd99892, -32'sd599859, 32'sd1203803, 32'sd619473, 32'sd903536, -32'sd703059, -32'sd771762, -32'sd2119200, -32'sd486262, -32'sd9642, -32'sd247194, -32'sd303410, 32'sd135983, 32'sd855564, 32'sd610154, 32'sd1300978, 32'sd640815, -32'sd216394, 32'sd1199640, 32'sd437366, 32'sd1755080, 32'sd421721, -32'sd70155, -32'sd176062, -32'sd943913, 32'sd40244, 32'sd1493316, -32'sd1115594, 32'sd529215, 32'sd440134, 32'sd1537607, 32'sd113281, 32'sd722383, -32'sd1089345, -32'sd1403534, -32'sd38707, 32'sd893274, -32'sd351594, 32'sd0, 32'sd180357, -32'sd550480, 32'sd57162, 32'sd776638, 32'sd805041, -32'sd419431, 32'sd340011, 32'sd932405, 32'sd206755, -32'sd598775, 32'sd1690818, 32'sd1364222, 32'sd946957, 32'sd1059163, 32'sd2929847, 32'sd1124400, -32'sd318182, -32'sd542887, 32'sd1011818, -32'sd1084843, -32'sd1238357, 32'sd149090, 32'sd192112, 32'sd985953, -32'sd637820, 32'sd1038722, 32'sd0, 32'sd0, 32'sd0, 32'sd1553018, 32'sd1584423, 32'sd955840, 32'sd612677, 32'sd2098679, 32'sd1268387, -32'sd594427, 32'sd802751, 32'sd1809085, 32'sd1878501, 32'sd1324564, 32'sd1998833, 32'sd840642, 32'sd586617, -32'sd2284962, 32'sd401307, -32'sd966528, -32'sd630425, -32'sd1897787, -32'sd1017699, -32'sd1913684, 32'sd773231, 32'sd417956, 32'sd699441, -32'sd557066, 32'sd0, 32'sd0, 32'sd0, 32'sd11804, 32'sd100502, 32'sd387453, 32'sd428579, -32'sd839585, 32'sd425706, 32'sd697230, -32'sd1354626, 32'sd1635709, 32'sd1268345, 32'sd501733, 32'sd2665632, 32'sd463468, -32'sd940044, -32'sd337930, -32'sd741769, -32'sd3526369, -32'sd1964269, -32'sd1600678, -32'sd3240096, -32'sd2187383, -32'sd393134, -32'sd2704757, -32'sd21613, 32'sd241156, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd60166, -32'sd1485085, 32'sd760820, -32'sd743026, 32'sd579074, 32'sd414794, 32'sd570135, 32'sd1808358, 32'sd708199, 32'sd202554, -32'sd293892, -32'sd1554049, 32'sd504357, -32'sd1248017, 32'sd1724123, 32'sd2256123, -32'sd1644458, -32'sd1892745, -32'sd150144, -32'sd679850, 32'sd94967, 32'sd1135210, -32'sd103882, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd556059, 32'sd1064520, -32'sd682534, -32'sd269682, -32'sd596771, -32'sd498058, -32'sd116568, -32'sd1450276, -32'sd713428, -32'sd480868, 32'sd730883, -32'sd1548615, -32'sd44320, -32'sd1737294, -32'sd646331, 32'sd848332, -32'sd1184200, 32'sd506285, -32'sd132044, -32'sd697986, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd656372, 32'sd486747, 32'sd194635, 32'sd1452752, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd709477, -32'sd485528, -32'sd579215, -32'sd8520, -32'sd120779, 32'sd364450, -32'sd341631, -32'sd1150123, -32'sd908877, -32'sd687690, 32'sd395310, -32'sd25904, 32'sd787255, 32'sd375887, -32'sd30246, -32'sd585769, 32'sd292301, -32'sd799329, -32'sd1530832, 32'sd963324, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd65759, 32'sd597795, -32'sd174068, -32'sd1738534, -32'sd1172722, 32'sd672419, -32'sd1035497, -32'sd133643, -32'sd60886, -32'sd192556, -32'sd308366, -32'sd2411966, -32'sd1183261, -32'sd1918300, -32'sd292077, -32'sd359298, -32'sd983630, 32'sd965355, 32'sd232263, -32'sd119238, -32'sd855743, -32'sd752522, 32'sd1020839, -32'sd168920, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1174652, -32'sd1366127, 32'sd1291123, 32'sd923, 32'sd1030338, -32'sd1037902, -32'sd600784, -32'sd1004182, 32'sd1702293, -32'sd979369, 32'sd235063, -32'sd3445688, -32'sd239803, -32'sd336597, -32'sd698984, 32'sd1072594, 32'sd2866915, -32'sd654692, 32'sd77045, -32'sd1499721, 32'sd180661, 32'sd258019, -32'sd538021, 32'sd454578, -32'sd453521, 32'sd0, 32'sd0, 32'sd269570, 32'sd729993, -32'sd277143, -32'sd2646483, -32'sd1490251, 32'sd1686293, 32'sd98462, 32'sd145370, -32'sd1090798, 32'sd115564, -32'sd483845, -32'sd2329133, -32'sd889644, -32'sd2370962, 32'sd108799, -32'sd287357, 32'sd161485, -32'sd1277085, -32'sd183633, -32'sd1027243, -32'sd170380, 32'sd519847, -32'sd899040, -32'sd1228901, 32'sd1030219, 32'sd442652, 32'sd1073650, 32'sd0, 32'sd553111, -32'sd552349, 32'sd170674, 32'sd376320, -32'sd364916, 32'sd570292, 32'sd2420609, 32'sd1875574, -32'sd339177, 32'sd1561796, 32'sd67148, 32'sd1460503, 32'sd760869, 32'sd844949, -32'sd1009589, -32'sd884321, -32'sd562882, -32'sd462620, -32'sd2036140, -32'sd1776002, -32'sd1491324, 32'sd112216, -32'sd716421, 32'sd504381, 32'sd1048947, 32'sd213741, -32'sd1302272, 32'sd0, -32'sd94184, -32'sd705680, -32'sd137890, 32'sd600120, 32'sd700958, -32'sd391941, 32'sd1117318, -32'sd255993, 32'sd2564976, 32'sd181579, 32'sd64190, -32'sd256699, 32'sd2180010, 32'sd2593398, -32'sd665169, 32'sd1031405, 32'sd1466573, 32'sd176922, 32'sd448167, -32'sd838351, 32'sd1504809, 32'sd1155964, -32'sd835387, 32'sd402468, -32'sd1560814, -32'sd1116085, -32'sd1151152, 32'sd279385, -32'sd376646, 32'sd598201, 32'sd317422, 32'sd412600, -32'sd1579680, 32'sd1545957, -32'sd449524, -32'sd84877, 32'sd1348814, 32'sd179576, 32'sd271949, 32'sd568528, 32'sd3975836, 32'sd1756963, -32'sd2385812, 32'sd602213, -32'sd1233588, -32'sd1840089, -32'sd856848, 32'sd2163604, -32'sd447263, -32'sd1576287, 32'sd184811, 32'sd67666, -32'sd2296211, -32'sd386239, -32'sd756118, -32'sd437730, 32'sd1256072, 32'sd1999639, -32'sd1107349, 32'sd473029, 32'sd1342100, 32'sd367807, 32'sd808536, 32'sd1340284, 32'sd2405234, 32'sd742711, 32'sd2689023, 32'sd1296850, -32'sd360770, 32'sd1504378, 32'sd1269759, -32'sd1106928, -32'sd111811, -32'sd434539, -32'sd707220, 32'sd741119, -32'sd881507, -32'sd1915946, -32'sd353959, -32'sd462271, -32'sd293320, -32'sd267588, 32'sd608028, 32'sd662508, 32'sd1638161, 32'sd676345, -32'sd396601, 32'sd979400, 32'sd2115166, 32'sd1870793, -32'sd404214, -32'sd862520, 32'sd422058, 32'sd1572481, 32'sd1448881, 32'sd1487104, -32'sd253335, 32'sd3110750, 32'sd1674996, 32'sd638358, 32'sd1282659, 32'sd963014, -32'sd1827594, -32'sd292923, -32'sd1403180, 32'sd1103022, -32'sd1906126, -32'sd49664, 32'sd189171, -32'sd1266069, 32'sd618007, 32'sd774224, 32'sd396487, 32'sd1200005, -32'sd1110617, 32'sd491196, -32'sd103437, 32'sd1960298, -32'sd1634275, 32'sd2104730, -32'sd786235, 32'sd388539, -32'sd1541033, -32'sd2044006, 32'sd280719, 32'sd2332824, 32'sd2662418, 32'sd1484980, -32'sd1015662, 32'sd1038685, -32'sd991100, -32'sd751543, -32'sd1851752, 32'sd345700, 32'sd697966, 32'sd884732, 32'sd2013657, 32'sd480973, 32'sd192306, 32'sd712917, 32'sd567997, 32'sd1474169, 32'sd1665669, 32'sd1475452, -32'sd246336, 32'sd1371735, 32'sd2864410, 32'sd1148401, 32'sd963732, -32'sd522434, 32'sd694910, -32'sd318784, 32'sd794060, 32'sd1914063, 32'sd2219516, 32'sd3399336, -32'sd449881, -32'sd607737, -32'sd256982, -32'sd477175, -32'sd1762801, -32'sd248489, 32'sd497703, -32'sd188403, 32'sd1230046, 32'sd624276, -32'sd1051204, 32'sd86039, 32'sd628063, -32'sd810061, -32'sd311254, -32'sd2381545, -32'sd2784885, -32'sd1379567, -32'sd454716, 32'sd1649186, 32'sd70442, -32'sd514105, -32'sd1434874, -32'sd483932, 32'sd1217566, 32'sd293403, 32'sd3785917, 32'sd1499692, -32'sd87580, 32'sd502958, -32'sd1957419, -32'sd2464764, -32'sd2051236, -32'sd2125953, -32'sd1109774, -32'sd1421133, 32'sd895847, 32'sd496181, -32'sd564110, 32'sd117565, -32'sd1182923, 32'sd521300, -32'sd530138, -32'sd3279983, -32'sd1436623, -32'sd1228794, -32'sd51449, 32'sd1519134, -32'sd301177, -32'sd489797, -32'sd1839395, -32'sd1027011, -32'sd251885, -32'sd2298443, -32'sd383106, 32'sd2105864, 32'sd301949, -32'sd571861, -32'sd2980751, -32'sd3281947, -32'sd1554577, -32'sd260583, 32'sd1170851, 32'sd259545, 32'sd228167, 32'sd349362, 32'sd110698, -32'sd366685, -32'sd430195, 32'sd629764, -32'sd1649342, -32'sd1479798, -32'sd2715006, -32'sd871748, -32'sd1054635, -32'sd955091, 32'sd270611, 32'sd1434885, 32'sd583196, -32'sd185237, -32'sd2469918, -32'sd868355, -32'sd742482, 32'sd493259, 32'sd1378964, -32'sd621239, -32'sd2346000, -32'sd1541313, -32'sd159596, -32'sd988980, -32'sd370443, -32'sd1304712, -32'sd546785, 32'sd522403, -32'sd966509, -32'sd426793, 32'sd794088, -32'sd88385, -32'sd1265759, -32'sd679053, -32'sd3389173, -32'sd4028841, -32'sd693504, -32'sd1071081, 32'sd1607771, 32'sd2822754, 32'sd2250159, 32'sd328340, -32'sd1624956, 32'sd841014, 32'sd1407246, 32'sd968826, 32'sd3526037, 32'sd803079, -32'sd2246237, 32'sd737557, 32'sd562458, 32'sd1342830, 32'sd267116, 32'sd119273, -32'sd1122881, -32'sd464348, -32'sd192285, 32'sd102059, -32'sd793990, 32'sd376016, -32'sd2038240, -32'sd579437, -32'sd1877685, -32'sd1535104, 32'sd1333568, 32'sd1774547, 32'sd1937221, 32'sd1086128, 32'sd2340348, 32'sd2354367, 32'sd2251695, 32'sd638023, 32'sd3402720, 32'sd2962730, 32'sd3062177, 32'sd200291, 32'sd93743, 32'sd463114, 32'sd1052233, 32'sd656641, 32'sd1338327, -32'sd2141952, -32'sd1179445, 32'sd652402, 32'sd157823, 32'sd0, -32'sd445090, -32'sd250261, -32'sd1140025, -32'sd159709, -32'sd412077, 32'sd1468791, 32'sd1952828, 32'sd1275258, 32'sd215493, 32'sd465594, 32'sd136398, 32'sd796808, -32'sd439357, 32'sd418056, 32'sd2519867, 32'sd233862, 32'sd591863, 32'sd340416, -32'sd1517923, 32'sd745683, 32'sd2100365, 32'sd2152937, -32'sd579528, 32'sd774566, 32'sd119295, 32'sd244455, 32'sd150301, -32'sd679520, 32'sd305130, 32'sd904341, -32'sd1498337, -32'sd1337974, -32'sd975939, -32'sd1910961, -32'sd120763, -32'sd1574097, -32'sd897518, -32'sd940527, -32'sd1780860, -32'sd1864428, 32'sd320094, 32'sd793939, 32'sd2004314, 32'sd784297, 32'sd1276842, -32'sd3052654, -32'sd421692, 32'sd1219346, -32'sd963201, -32'sd854407, -32'sd654082, -32'sd438357, -32'sd1594355, 32'sd1682282, -32'sd1407659, 32'sd900670, -32'sd86567, -32'sd77681, -32'sd112807, -32'sd1266249, 32'sd277111, -32'sd3637683, -32'sd3077884, -32'sd3520110, -32'sd2712484, -32'sd4136680, -32'sd3667084, -32'sd1503619, -32'sd336168, -32'sd1006983, 32'sd407992, -32'sd1666486, -32'sd1441893, -32'sd1844240, -32'sd998737, -32'sd944318, -32'sd672934, -32'sd1169600, 32'sd592658, -32'sd972398, -32'sd1603285, -32'sd1243182, -32'sd86768, 32'sd0, 32'sd37580, -32'sd986605, -32'sd831507, -32'sd1038645, -32'sd3323922, -32'sd3963206, -32'sd1768753, -32'sd3016375, -32'sd1969804, -32'sd2608039, -32'sd2163580, -32'sd405866, 32'sd1036013, -32'sd1785281, -32'sd2433171, -32'sd2446506, -32'sd3661997, -32'sd2018400, -32'sd3059804, -32'sd297648, -32'sd658716, 32'sd359099, -32'sd191261, 32'sd36149, -32'sd801596, -32'sd2028612, 32'sd184810, 32'sd376100, 32'sd402469, -32'sd1218757, 32'sd747824, 32'sd1905158, -32'sd960800, -32'sd3222539, -32'sd1881311, -32'sd2390230, 32'sd544417, -32'sd1283951, -32'sd552346, 32'sd1838936, -32'sd723534, -32'sd1992488, -32'sd1473454, -32'sd212948, -32'sd1630526, -32'sd5157149, -32'sd1992912, -32'sd2291519, -32'sd1143621, 32'sd1507493, 32'sd592874, -32'sd199092, -32'sd270410, -32'sd204677, 32'sd584469, -32'sd167268, 32'sd664830, 32'sd180661, -32'sd515121, 32'sd77693, 32'sd779966, 32'sd717145, -32'sd797350, 32'sd246425, -32'sd213887, 32'sd3417551, 32'sd1110404, 32'sd1592807, -32'sd2035086, -32'sd1246539, -32'sd152608, -32'sd1036241, -32'sd1342504, -32'sd2958249, -32'sd1705675, -32'sd2586075, -32'sd2230796, 32'sd1238740, -32'sd1526904, -32'sd336911, 32'sd912259, -32'sd120454, -32'sd726035, 32'sd0, 32'sd1254487, -32'sd611646, 32'sd1324068, -32'sd652745, 32'sd248317, 32'sd1517253, 32'sd1007907, 32'sd608448, 32'sd1187442, 32'sd585804, 32'sd789044, 32'sd522370, -32'sd230406, 32'sd129969, 32'sd226692, 32'sd188083, 32'sd831188, -32'sd1285434, -32'sd1810273, -32'sd1462316, 32'sd122775, -32'sd436970, 32'sd241624, 32'sd766399, -32'sd227907, -32'sd1199751, 32'sd0, 32'sd0, 32'sd0, -32'sd380037, 32'sd414378, -32'sd1196544, 32'sd1156046, 32'sd1234314, 32'sd740621, 32'sd1195004, -32'sd356735, 32'sd1449275, 32'sd225809, 32'sd307201, -32'sd766676, 32'sd39666, -32'sd1304697, -32'sd64174, -32'sd914904, -32'sd1090711, 32'sd906255, 32'sd175114, 32'sd331899, 32'sd1245664, 32'sd464159, 32'sd382139, -32'sd84005, 32'sd498121, 32'sd0, 32'sd0, 32'sd0, 32'sd1430428, 32'sd923455, -32'sd438239, 32'sd1380261, -32'sd71878, 32'sd147189, -32'sd169006, 32'sd275463, 32'sd1135864, -32'sd1136107, -32'sd422721, -32'sd1855565, -32'sd2185383, -32'sd839251, -32'sd941435, 32'sd1012520, -32'sd1056664, -32'sd462803, -32'sd760662, -32'sd107457, -32'sd1233531, -32'sd316379, 32'sd327974, 32'sd814978, -32'sd443356, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd189779, 32'sd90513, -32'sd118340, -32'sd911275, 32'sd204196, 32'sd1010200, 32'sd605828, 32'sd2843243, 32'sd972106, 32'sd1049101, 32'sd503567, 32'sd272819, 32'sd409044, -32'sd415914, 32'sd748921, -32'sd27354, 32'sd1087354, 32'sd162200, -32'sd399189, 32'sd715555, 32'sd1139471, 32'sd1102512, 32'sd860775, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1037982, -32'sd37442, -32'sd18652, 32'sd1372761, -32'sd1377304, -32'sd424079, 32'sd950257, -32'sd270296, -32'sd1135703, 32'sd627948, 32'sd2021693, 32'sd850295, 32'sd2325352, 32'sd952053, 32'sd789467, 32'sd841697, -32'sd420479, 32'sd1456661, 32'sd1689177, 32'sd1992655, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd522226, 32'sd617847, 32'sd1637122, -32'sd221470, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd214246, 32'sd1009615, -32'sd104613, 32'sd69175, 32'sd169761, 32'sd947766, -32'sd1417954, 32'sd262449, -32'sd531132, -32'sd78440, 32'sd615760, 32'sd905722, 32'sd560573, 32'sd748859, -32'sd649414, -32'sd215843, 32'sd920239, -32'sd585314, 32'sd409506, 32'sd11285, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd942499, 32'sd68310, 32'sd1060044, 32'sd565121, 32'sd107179, -32'sd450088, -32'sd697098, -32'sd787065, 32'sd984427, 32'sd659176, -32'sd754988, -32'sd2962535, 32'sd870256, 32'sd384726, 32'sd2199533, 32'sd1991439, 32'sd320961, 32'sd121505, -32'sd1623455, 32'sd391000, 32'sd555053, 32'sd1133370, -32'sd1023464, 32'sd894892, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1197813, -32'sd584621, -32'sd495055, -32'sd499076, 32'sd1362381, 32'sd933875, 32'sd153460, 32'sd2732, 32'sd1029190, 32'sd207525, -32'sd314470, -32'sd2354600, -32'sd1679899, -32'sd1575593, -32'sd548553, 32'sd944512, 32'sd725748, 32'sd521917, 32'sd370898, 32'sd1888427, -32'sd267818, 32'sd580085, -32'sd1213584, -32'sd507422, 32'sd394468, 32'sd0, 32'sd0, 32'sd256603, -32'sd259536, 32'sd1374034, 32'sd616863, -32'sd1622707, -32'sd2015456, -32'sd1635792, -32'sd1334494, -32'sd1715547, -32'sd488594, 32'sd1810910, 32'sd337230, -32'sd212431, -32'sd2099631, -32'sd1384387, -32'sd412201, -32'sd1498000, -32'sd1261352, -32'sd770353, 32'sd1134165, 32'sd2024506, -32'sd90219, -32'sd220784, -32'sd888701, -32'sd1240851, -32'sd748364, -32'sd90877, 32'sd0, 32'sd1025371, 32'sd425400, 32'sd1151248, 32'sd442431, 32'sd1019015, 32'sd1544496, -32'sd258121, 32'sd1774502, 32'sd283621, -32'sd543390, 32'sd347589, -32'sd2252797, -32'sd2406494, -32'sd2668929, -32'sd2623751, -32'sd717893, -32'sd601621, -32'sd802552, 32'sd50057, -32'sd152593, 32'sd1035563, 32'sd239135, -32'sd1255211, -32'sd359061, -32'sd686802, -32'sd658573, 32'sd650821, 32'sd0, -32'sd144147, -32'sd322162, -32'sd734364, 32'sd2125775, 32'sd1867220, 32'sd1205296, 32'sd810227, -32'sd1670089, 32'sd859653, 32'sd1690179, -32'sd1369582, 32'sd2116119, 32'sd967235, -32'sd1078247, -32'sd616562, 32'sd555160, 32'sd2172148, 32'sd847349, 32'sd947155, -32'sd1406966, 32'sd1943979, 32'sd241669, -32'sd761203, -32'sd1452791, -32'sd855532, -32'sd1083787, 32'sd681093, 32'sd579725, -32'sd377596, 32'sd1037285, -32'sd966313, 32'sd838122, -32'sd930847, 32'sd1318534, 32'sd901696, -32'sd97930, 32'sd2166469, 32'sd1312088, 32'sd1020766, 32'sd1643032, 32'sd1568831, -32'sd739361, -32'sd904933, 32'sd2121829, 32'sd168702, 32'sd1587449, 32'sd1188672, 32'sd1733431, -32'sd8055, 32'sd1460838, -32'sd25978, 32'sd682278, 32'sd971064, -32'sd1114671, -32'sd1573505, -32'sd521576, -32'sd306509, 32'sd1111761, 32'sd594438, -32'sd807123, -32'sd544747, -32'sd985077, 32'sd967443, 32'sd668033, 32'sd3273403, 32'sd2432675, 32'sd2113347, -32'sd297893, 32'sd845681, -32'sd284161, 32'sd2047339, 32'sd861593, 32'sd1774293, 32'sd1549403, 32'sd1142994, -32'sd577072, -32'sd738734, 32'sd1789547, -32'sd1347735, 32'sd859451, -32'sd752527, -32'sd1676415, 32'sd2760, 32'sd973093, 32'sd1139235, -32'sd1008768, -32'sd712116, -32'sd632980, 32'sd83173, 32'sd1408583, 32'sd393030, 32'sd950691, 32'sd936912, 32'sd1472857, 32'sd509607, 32'sd767531, 32'sd1567168, 32'sd1134678, -32'sd495744, 32'sd170856, 32'sd151586, -32'sd100195, -32'sd1752566, -32'sd630073, 32'sd881853, -32'sd257448, -32'sd163422, -32'sd461661, -32'sd2955446, -32'sd89405, -32'sd192993, 32'sd1366282, -32'sd929141, 32'sd503155, -32'sd2551764, -32'sd662096, 32'sd1311636, 32'sd480596, 32'sd47058, -32'sd702064, -32'sd580345, 32'sd1068227, 32'sd1887864, 32'sd33389, 32'sd1031568, -32'sd1512467, -32'sd1691636, -32'sd1112147, 32'sd583882, 32'sd2160026, 32'sd1251441, -32'sd171160, 32'sd402993, -32'sd738786, 32'sd655345, 32'sd812120, -32'sd2081959, -32'sd10729, 32'sd204664, 32'sd699987, -32'sd52131, -32'sd1913328, -32'sd270316, -32'sd165156, -32'sd3908, 32'sd755467, 32'sd1957969, -32'sd366787, 32'sd1933768, 32'sd648603, 32'sd2303989, 32'sd1318139, -32'sd267620, 32'sd31895, 32'sd132155, -32'sd863175, 32'sd2155830, 32'sd3349434, -32'sd513680, 32'sd918456, -32'sd1294382, -32'sd740162, 32'sd531728, 32'sd755507, -32'sd187614, 32'sd663331, 32'sd149236, -32'sd39546, 32'sd346558, -32'sd230054, -32'sd351506, -32'sd2177474, -32'sd602469, 32'sd526225, -32'sd911003, 32'sd667856, -32'sd593640, 32'sd1028651, 32'sd540552, -32'sd1275337, -32'sd1797346, -32'sd2879283, 32'sd1620606, 32'sd2474637, 32'sd1493636, 32'sd657067, -32'sd951837, -32'sd696783, 32'sd336600, -32'sd841732, -32'sd2200809, 32'sd1142142, 32'sd1115628, -32'sd1063186, 32'sd935315, 32'sd226802, -32'sd68736, 32'sd884289, -32'sd2427591, -32'sd1385807, -32'sd703365, -32'sd213653, 32'sd123331, 32'sd1025225, -32'sd1125334, 32'sd1268630, 32'sd959161, -32'sd1483858, -32'sd3673416, -32'sd2325541, 32'sd211745, 32'sd2269511, -32'sd597743, -32'sd308408, -32'sd2422428, -32'sd1583746, 32'sd373309, -32'sd98796, -32'sd592942, -32'sd1851812, -32'sd1784755, -32'sd1008589, 32'sd1434886, 32'sd186731, 32'sd231229, -32'sd75998, -32'sd194579, -32'sd440713, -32'sd1391570, -32'sd1901746, 32'sd266539, 32'sd328002, -32'sd90661, 32'sd605237, -32'sd609587, -32'sd2055412, -32'sd1894948, -32'sd741159, -32'sd1301329, 32'sd1216176, 32'sd1410090, -32'sd647596, -32'sd792155, 32'sd882516, -32'sd1858318, -32'sd1932871, -32'sd3182859, -32'sd1745822, 32'sd1309418, -32'sd177238, 32'sd689142, -32'sd536226, 32'sd482373, -32'sd259688, -32'sd900551, -32'sd1405003, -32'sd2094542, -32'sd1078151, 32'sd561478, -32'sd361175, -32'sd1026767, 32'sd88747, -32'sd690208, -32'sd1914326, -32'sd2472458, -32'sd1158079, -32'sd1268039, 32'sd1295699, 32'sd1705051, 32'sd1126521, -32'sd2575962, 32'sd339381, -32'sd853726, -32'sd1421745, -32'sd1749706, 32'sd473464, 32'sd1183915, 32'sd1481835, -32'sd621327, 32'sd536509, 32'sd589563, 32'sd1432833, -32'sd654923, 32'sd735336, -32'sd88809, 32'sd262572, 32'sd2891566, 32'sd2104082, -32'sd535017, 32'sd1886531, -32'sd861637, -32'sd434435, -32'sd636411, -32'sd126911, 32'sd1004364, 32'sd2838862, 32'sd1392562, -32'sd1514804, -32'sd610698, 32'sd704346, 32'sd212205, 32'sd627154, 32'sd132331, 32'sd541655, -32'sd685409, -32'sd770966, 32'sd1110238, 32'sd0, 32'sd369409, -32'sd409726, -32'sd318661, 32'sd102270, 32'sd1711732, 32'sd243436, 32'sd1908208, 32'sd1068161, -32'sd639520, 32'sd233600, 32'sd311563, -32'sd2246607, -32'sd2431453, 32'sd16923, 32'sd2622729, 32'sd1389106, 32'sd331838, 32'sd736465, -32'sd21067, 32'sd1980670, 32'sd3045750, 32'sd3552653, 32'sd1049904, -32'sd111825, 32'sd850280, 32'sd977017, 32'sd595252, 32'sd894120, -32'sd20028, 32'sd53633, -32'sd1874402, 32'sd2300367, -32'sd651611, 32'sd19827, -32'sd551319, 32'sd14087, -32'sd1635994, -32'sd1946563, -32'sd3499616, -32'sd2878335, -32'sd1785447, -32'sd274810, 32'sd265443, 32'sd1743973, 32'sd696661, 32'sd408652, -32'sd1185636, -32'sd389582, 32'sd875846, 32'sd2869888, 32'sd1388726, 32'sd971638, 32'sd1762694, 32'sd1287050, 32'sd934343, 32'sd604773, -32'sd623510, -32'sd1368093, 32'sd954396, 32'sd1435419, 32'sd312681, -32'sd695569, -32'sd466832, -32'sd1580519, -32'sd1661674, -32'sd1887440, -32'sd2542240, -32'sd2984548, -32'sd1553339, 32'sd854563, -32'sd1583944, -32'sd1623232, -32'sd1450579, -32'sd1580765, 32'sd84780, 32'sd857363, 32'sd2329808, 32'sd2794540, 32'sd2699345, 32'sd273785, 32'sd407815, 32'sd773252, 32'sd706085, 32'sd0, -32'sd864049, -32'sd955881, 32'sd565137, 32'sd2314653, 32'sd976392, -32'sd1210526, -32'sd287652, -32'sd774119, -32'sd1702709, -32'sd2295825, -32'sd1077590, -32'sd315334, -32'sd1348230, -32'sd126762, -32'sd766530, -32'sd1126915, -32'sd1570693, -32'sd2537527, -32'sd943190, -32'sd1118573, 32'sd598649, 32'sd1742609, 32'sd2280662, 32'sd2783446, 32'sd22502, 32'sd187413, 32'sd471868, 32'sd1003220, 32'sd299484, 32'sd1057683, -32'sd39773, 32'sd112689, 32'sd803362, -32'sd1563503, -32'sd119103, -32'sd2694470, 32'sd192653, -32'sd1556264, 32'sd229868, 32'sd866937, 32'sd975547, -32'sd107883, -32'sd1964947, -32'sd2135019, -32'sd2118053, -32'sd3358174, -32'sd1465696, -32'sd3023729, -32'sd1217481, 32'sd1063721, -32'sd55888, -32'sd1693396, 32'sd199388, 32'sd342607, 32'sd498932, -32'sd217171, -32'sd662961, 32'sd649474, -32'sd861168, -32'sd706503, -32'sd1600283, -32'sd157000, -32'sd753342, -32'sd646115, -32'sd1328416, 32'sd600113, -32'sd198871, 32'sd567345, -32'sd240646, -32'sd206633, -32'sd2246786, -32'sd305567, -32'sd1714039, -32'sd1750913, -32'sd2405302, -32'sd2194806, -32'sd1184608, 32'sd349261, -32'sd2582427, -32'sd915622, -32'sd471751, 32'sd634033, 32'sd1472855, 32'sd0, 32'sd199515, -32'sd1372553, -32'sd1576466, -32'sd1023489, 32'sd532426, 32'sd1223411, -32'sd665179, -32'sd907985, -32'sd459352, -32'sd715847, 32'sd197349, 32'sd827673, -32'sd872857, -32'sd1242604, 32'sd414041, -32'sd594686, -32'sd1037356, -32'sd901723, -32'sd1818710, -32'sd2229238, -32'sd917784, -32'sd732039, 32'sd296341, 32'sd323156, -32'sd300607, -32'sd803449, 32'sd0, 32'sd0, 32'sd0, -32'sd953067, -32'sd1568250, 32'sd1889742, 32'sd1074584, -32'sd851084, -32'sd237129, -32'sd467335, -32'sd493028, 32'sd1351163, 32'sd431944, 32'sd596472, -32'sd551631, -32'sd575410, -32'sd1203699, -32'sd37551, 32'sd472074, -32'sd1939267, 32'sd877058, -32'sd646768, 32'sd861082, -32'sd546124, -32'sd744383, -32'sd971255, -32'sd764569, 32'sd941225, 32'sd0, 32'sd0, 32'sd0, 32'sd236600, 32'sd73594, 32'sd795259, 32'sd1625651, -32'sd1776758, 32'sd170435, 32'sd1154014, -32'sd1109907, 32'sd221962, 32'sd2278780, 32'sd544666, -32'sd776759, 32'sd556486, -32'sd1288514, -32'sd704380, 32'sd676617, -32'sd825902, 32'sd540113, -32'sd269211, 32'sd796027, -32'sd551628, -32'sd459818, -32'sd166179, -32'sd18935, 32'sd996473, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1155089, -32'sd2240950, 32'sd607942, -32'sd611616, 32'sd1059375, -32'sd50198, 32'sd242510, 32'sd504775, 32'sd792791, 32'sd1867737, 32'sd2525838, 32'sd2366690, 32'sd6226, 32'sd998073, -32'sd1029710, 32'sd354250, 32'sd625442, 32'sd32976, 32'sd1015224, 32'sd961066, 32'sd1448585, 32'sd393108, 32'sd615475, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd272774, 32'sd652109, 32'sd829524, -32'sd344452, 32'sd393320, -32'sd690923, 32'sd1196807, 32'sd1298923, 32'sd204206, 32'sd1137078, 32'sd1994876, 32'sd601358, 32'sd1415776, 32'sd262545, -32'sd522877, -32'sd1138196, 32'sd178021, 32'sd131470, 32'sd1443247, -32'sd54284, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1008619, -32'sd479956, 32'sd282286, -32'sd655566, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd449342, -32'sd614928, -32'sd1025005, -32'sd1095308, -32'sd228776, 32'sd1860077, 32'sd1004922, -32'sd1455673, -32'sd2351598, -32'sd103098, 32'sd344280, 32'sd171130, -32'sd2048578, -32'sd128795, -32'sd124791, 32'sd144739, -32'sd1594867, 32'sd636322, -32'sd708045, -32'sd1952, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd249033, 32'sd105842, -32'sd1186395, 32'sd1321501, 32'sd1296720, -32'sd635864, -32'sd772161, 32'sd75243, -32'sd138272, 32'sd587738, 32'sd838224, -32'sd372985, 32'sd1953999, 32'sd1176447, -32'sd75671, 32'sd133031, -32'sd455017, 32'sd389818, -32'sd408778, -32'sd895600, -32'sd1231466, -32'sd48828, -32'sd431744, -32'sd578467, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd234794, 32'sd1063080, 32'sd477370, -32'sd1369492, -32'sd1125115, -32'sd411767, -32'sd790356, 32'sd297784, -32'sd658647, -32'sd752929, -32'sd221251, -32'sd439484, -32'sd1576983, 32'sd558851, 32'sd376034, -32'sd1135030, -32'sd1155561, 32'sd606447, 32'sd867632, 32'sd395167, -32'sd901634, -32'sd554792, -32'sd614618, -32'sd691404, -32'sd1576184, 32'sd0, 32'sd0, 32'sd266965, 32'sd699110, -32'sd217302, 32'sd48574, -32'sd435364, 32'sd180730, 32'sd570736, -32'sd224459, -32'sd1861227, -32'sd1610111, -32'sd961378, -32'sd1582796, -32'sd310316, -32'sd1867201, -32'sd1581719, -32'sd2068013, -32'sd1429407, -32'sd301330, -32'sd2065301, -32'sd253090, 32'sd17443, -32'sd560154, -32'sd2423741, 32'sd1220004, 32'sd1100813, 32'sd1470133, -32'sd304852, 32'sd0, -32'sd665753, -32'sd746665, -32'sd591290, 32'sd943804, -32'sd1313731, -32'sd1181822, -32'sd1544660, -32'sd1498414, -32'sd2228079, 32'sd1029439, -32'sd533423, -32'sd155852, -32'sd319940, -32'sd810022, -32'sd2876784, 32'sd94204, -32'sd2176614, -32'sd1470991, 32'sd1373472, 32'sd804278, 32'sd544693, -32'sd1561705, -32'sd1556430, 32'sd1507373, 32'sd1831762, 32'sd815738, -32'sd877146, 32'sd0, -32'sd379930, 32'sd251691, -32'sd315423, 32'sd437530, -32'sd1687899, -32'sd1605648, -32'sd1634595, 32'sd127412, -32'sd1105033, -32'sd238905, 32'sd1619402, 32'sd1745047, 32'sd714324, -32'sd1679558, -32'sd607465, 32'sd2059432, 32'sd1556269, 32'sd391220, 32'sd1730405, -32'sd241734, -32'sd1092888, -32'sd2505184, -32'sd1387027, -32'sd1156559, 32'sd717413, 32'sd1511759, -32'sd80007, -32'sd700679, -32'sd174989, -32'sd1017983, 32'sd262586, -32'sd258874, -32'sd1309788, -32'sd2095484, -32'sd955905, -32'sd2073036, -32'sd1227684, 32'sd726429, -32'sd980916, 32'sd705798, 32'sd614928, 32'sd380774, 32'sd271254, -32'sd1855446, -32'sd1273340, 32'sd898587, 32'sd2860557, 32'sd358953, -32'sd112414, 32'sd736691, -32'sd2746125, -32'sd631898, -32'sd1011589, -32'sd1765002, 32'sd927633, -32'sd472015, 32'sd357236, -32'sd553376, -32'sd75585, 32'sd718828, -32'sd117546, 32'sd91781, -32'sd1313468, -32'sd1038822, -32'sd2427563, -32'sd2127061, 32'sd36956, -32'sd1467551, -32'sd1293642, 32'sd346371, -32'sd227387, -32'sd1945746, -32'sd1175478, 32'sd1257389, -32'sd914653, -32'sd229345, 32'sd1451372, -32'sd1045169, -32'sd1092939, 32'sd753023, -32'sd1709251, -32'sd164880, -32'sd1042003, 32'sd717380, 32'sd2087421, -32'sd1753185, 32'sd654805, 32'sd903236, -32'sd1562306, 32'sd1441140, -32'sd349866, -32'sd1223984, 32'sd1193504, -32'sd1501707, 32'sd60975, -32'sd1950525, 32'sd1309501, 32'sd1283983, 32'sd530235, -32'sd153638, 32'sd29663, -32'sd787427, -32'sd642512, -32'sd1354051, 32'sd2434962, -32'sd522250, -32'sd1859263, -32'sd1496884, -32'sd1820168, -32'sd1507587, -32'sd1267513, 32'sd1290614, -32'sd1036566, -32'sd1884697, 32'sd99737, -32'sd719420, -32'sd508165, 32'sd105042, -32'sd1852577, -32'sd226034, -32'sd352471, 32'sd1325141, -32'sd1300944, -32'sd1406517, -32'sd242128, 32'sd1740730, -32'sd391346, -32'sd388369, -32'sd3182085, -32'sd184637, 32'sd209654, -32'sd1195756, 32'sd1212913, -32'sd1266873, -32'sd1101718, -32'sd248377, -32'sd2374975, -32'sd173036, -32'sd1682259, 32'sd706259, -32'sd3431530, -32'sd348592, -32'sd511510, -32'sd14132, 32'sd1266505, 32'sd922914, 32'sd1069135, 32'sd1656695, 32'sd344007, -32'sd1044793, -32'sd3247146, -32'sd3989857, -32'sd2718463, -32'sd254427, -32'sd331196, -32'sd3882724, -32'sd2262036, 32'sd677732, -32'sd1010622, -32'sd90312, 32'sd246426, 32'sd542170, 32'sd563280, -32'sd280878, 32'sd459604, 32'sd1263171, 32'sd1069592, -32'sd1151695, -32'sd917114, 32'sd229175, -32'sd76224, 32'sd24667, 32'sd752263, 32'sd601024, -32'sd90714, 32'sd2337382, 32'sd1508417, -32'sd235910, -32'sd2205155, -32'sd5018838, -32'sd3659760, -32'sd1248916, -32'sd2803732, -32'sd2504480, 32'sd983059, 32'sd777223, -32'sd476322, 32'sd1348829, 32'sd2761451, -32'sd365772, 32'sd257151, 32'sd1388432, -32'sd901088, -32'sd1207448, -32'sd191698, -32'sd117959, -32'sd230044, -32'sd278338, -32'sd1615706, -32'sd1071423, 32'sd1840273, 32'sd1106351, 32'sd1084610, 32'sd1964418, 32'sd619869, 32'sd1376256, -32'sd123124, -32'sd1930566, -32'sd1756752, -32'sd770793, 32'sd2305681, 32'sd1272254, 32'sd1445812, 32'sd1400871, 32'sd1374675, 32'sd689375, 32'sd2543973, 32'sd1676713, 32'sd574958, -32'sd958359, 32'sd1973912, -32'sd30667, -32'sd507366, -32'sd482572, -32'sd991415, -32'sd794592, -32'sd732099, 32'sd251271, -32'sd675649, 32'sd2329318, 32'sd79371, 32'sd124776, 32'sd1455542, 32'sd4475854, 32'sd3137916, 32'sd1014848, 32'sd951891, 32'sd1557094, -32'sd176301, 32'sd1316231, 32'sd1959833, 32'sd807996, 32'sd643487, -32'sd711067, -32'sd389860, -32'sd992767, 32'sd331688, -32'sd421465, 32'sd1126744, 32'sd535096, -32'sd1067278, 32'sd188090, -32'sd550411, -32'sd102433, -32'sd446267, 32'sd263460, 32'sd743222, 32'sd2065277, 32'sd595252, 32'sd1646842, 32'sd3501713, 32'sd3883626, 32'sd2685672, 32'sd3873004, 32'sd1105126, 32'sd1420679, 32'sd586722, 32'sd411439, 32'sd1945246, 32'sd2537216, 32'sd667927, -32'sd744579, -32'sd910455, 32'sd436720, 32'sd872354, 32'sd420619, 32'sd2044658, 32'sd1787621, 32'sd719556, -32'sd615181, 32'sd486460, -32'sd1795512, -32'sd505881, 32'sd61812, 32'sd320408, 32'sd1888006, 32'sd1616332, 32'sd966897, 32'sd1151076, 32'sd258150, 32'sd1676498, 32'sd2772877, 32'sd3472677, -32'sd129879, -32'sd1537220, 32'sd1893715, 32'sd1387789, 32'sd446961, -32'sd676641, 32'sd1153665, -32'sd548785, 32'sd498005, 32'sd21509, 32'sd38978, -32'sd758974, -32'sd304980, 32'sd351729, 32'sd0, -32'sd498453, 32'sd340987, -32'sd14550, 32'sd704594, 32'sd191429, -32'sd340249, -32'sd169726, -32'sd200372, -32'sd1738063, -32'sd1010187, -32'sd607876, 32'sd2131284, 32'sd754984, 32'sd180581, 32'sd1756715, 32'sd397488, 32'sd608547, -32'sd1251391, -32'sd940177, 32'sd1053335, -32'sd203185, -32'sd1416768, -32'sd1358396, 32'sd586349, 32'sd467771, 32'sd85388, 32'sd112915, -32'sd530311, 32'sd782988, -32'sd1065393, -32'sd601891, 32'sd605080, 32'sd938584, 32'sd2836162, 32'sd1764823, -32'sd1325189, -32'sd2356175, 32'sd769172, -32'sd602195, -32'sd301312, 32'sd2357278, 32'sd2243664, -32'sd171050, 32'sd436817, -32'sd1094173, 32'sd796528, -32'sd1499754, -32'sd68443, -32'sd683608, 32'sd158352, -32'sd1137751, -32'sd801254, -32'sd1748669, -32'sd52247, -32'sd659536, -32'sd984484, 32'sd33259, 32'sd866034, 32'sd517736, -32'sd49617, 32'sd1187296, 32'sd100615, 32'sd817375, -32'sd1153349, -32'sd19007, -32'sd268836, 32'sd940496, 32'sd1985621, 32'sd2845255, 32'sd2515159, -32'sd753294, -32'sd373641, -32'sd1074991, -32'sd226713, 32'sd1094230, -32'sd1762736, 32'sd1445994, -32'sd362151, 32'sd535140, -32'sd2102155, 32'sd176027, 32'sd534586, -32'sd862602, 32'sd0, 32'sd254880, 32'sd1603076, -32'sd1901363, -32'sd1638923, -32'sd106655, -32'sd349920, 32'sd692758, -32'sd570242, -32'sd196459, 32'sd523208, 32'sd929830, 32'sd563094, 32'sd1559216, -32'sd836814, -32'sd1059895, -32'sd47336, 32'sd345391, 32'sd2203774, 32'sd68041, -32'sd545794, -32'sd503145, -32'sd462734, 32'sd509220, 32'sd181270, -32'sd67404, -32'sd670590, -32'sd933352, 32'sd37053, 32'sd476840, 32'sd2175406, -32'sd397813, 32'sd686999, 32'sd2859487, 32'sd1222346, -32'sd1432868, 32'sd1092293, -32'sd89591, 32'sd877265, 32'sd547707, -32'sd909751, -32'sd8683, 32'sd1497620, -32'sd26484, -32'sd2122623, 32'sd52760, -32'sd1364633, 32'sd177409, 32'sd249554, 32'sd21642, -32'sd1221070, 32'sd1312972, 32'sd2021320, -32'sd2141269, -32'sd295333, -32'sd154587, -32'sd410381, 32'sd1013475, 32'sd1361210, -32'sd967272, 32'sd1656839, -32'sd895532, -32'sd947631, 32'sd178358, -32'sd60733, -32'sd1214451, -32'sd1748785, -32'sd1160064, -32'sd474898, -32'sd1424141, -32'sd2250729, -32'sd2581159, -32'sd387165, -32'sd90489, -32'sd1065894, -32'sd1053557, -32'sd619808, -32'sd1206124, 32'sd1160993, 32'sd2265804, 32'sd427671, -32'sd325110, -32'sd409127, -32'sd466124, 32'sd0, -32'sd279006, 32'sd342237, 32'sd572845, 32'sd2066788, 32'sd2466059, -32'sd610613, 32'sd188545, -32'sd379202, -32'sd1170029, 32'sd320519, -32'sd117394, -32'sd1846185, -32'sd1249785, 32'sd162251, 32'sd621567, 32'sd1183604, 32'sd772340, 32'sd643100, -32'sd1093125, 32'sd1712935, 32'sd456393, 32'sd1361936, 32'sd1072700, -32'sd40050, -32'sd188383, -32'sd693632, 32'sd0, 32'sd0, 32'sd0, -32'sd333183, -32'sd290206, 32'sd1395500, -32'sd1013890, 32'sd203576, 32'sd558838, 32'sd293305, 32'sd1039213, -32'sd982547, -32'sd1487192, 32'sd587641, 32'sd105089, 32'sd9406, 32'sd1085891, -32'sd1248179, 32'sd164305, 32'sd1397090, 32'sd135034, 32'sd48291, -32'sd387214, 32'sd1820885, -32'sd67845, -32'sd126065, -32'sd580459, 32'sd1447043, 32'sd0, 32'sd0, 32'sd0, -32'sd836221, 32'sd337621, -32'sd518205, -32'sd1648109, 32'sd918758, -32'sd1161057, -32'sd615548, 32'sd16139, 32'sd1949007, 32'sd637263, -32'sd1636659, -32'sd2882576, -32'sd387182, -32'sd1945470, 32'sd457739, -32'sd1050886, 32'sd181957, 32'sd180133, 32'sd35773, 32'sd408804, 32'sd295771, 32'sd283515, -32'sd335732, 32'sd233166, 32'sd1371346, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd364310, 32'sd1475913, -32'sd1318131, 32'sd283471, -32'sd662509, -32'sd325312, 32'sd407591, -32'sd153863, -32'sd2153274, -32'sd1185790, 32'sd1631560, -32'sd354642, -32'sd1455249, 32'sd2510324, 32'sd1039809, 32'sd1537128, -32'sd2395, -32'sd157070, -32'sd1223409, 32'sd132711, 32'sd784989, -32'sd216665, -32'sd865073, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1077074, -32'sd536838, 32'sd1146042, 32'sd1011717, -32'sd327884, -32'sd311243, 32'sd1052724, 32'sd835928, -32'sd223561, -32'sd352651, 32'sd969231, -32'sd69303, -32'sd1458376, -32'sd665612, 32'sd414874, 32'sd626769, -32'sd121320, -32'sd255764, -32'sd984746, -32'sd781040, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd389150, 32'sd663008, 32'sd1148212, -32'sd130944, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1227313, 32'sd413243, 32'sd266429, 32'sd1259773, 32'sd1455900, 32'sd929599, -32'sd1180102, 32'sd115199, 32'sd363646, 32'sd893297, -32'sd1151469, 32'sd1209629, 32'sd886273, 32'sd1872515, 32'sd1104323, -32'sd187965, -32'sd307364, 32'sd262407, -32'sd81055, 32'sd372959, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd143826, 32'sd89802, 32'sd788606, 32'sd342564, 32'sd413502, 32'sd246686, -32'sd1754282, 32'sd1394291, -32'sd164771, -32'sd268949, -32'sd133008, -32'sd411338, 32'sd530079, 32'sd2497883, 32'sd838584, 32'sd1135936, -32'sd920691, 32'sd1290270, -32'sd430956, 32'sd1035593, -32'sd934059, -32'sd684628, 32'sd329012, 32'sd1068785, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd404417, -32'sd611872, -32'sd64478, -32'sd1249863, 32'sd108753, 32'sd347959, -32'sd1497382, -32'sd242793, -32'sd715852, -32'sd1440204, -32'sd234430, -32'sd558968, -32'sd426762, -32'sd727852, 32'sd482811, -32'sd784207, -32'sd1418911, 32'sd947706, -32'sd126066, -32'sd775733, -32'sd425155, 32'sd754986, 32'sd1265942, 32'sd301616, 32'sd657395, 32'sd0, 32'sd0, 32'sd165229, 32'sd146373, -32'sd1878464, -32'sd174811, 32'sd1755648, -32'sd1137631, -32'sd1620497, -32'sd1347054, -32'sd519941, -32'sd20732, 32'sd1305872, -32'sd726017, -32'sd1081185, -32'sd1573706, -32'sd1391640, 32'sd1899983, -32'sd1417670, -32'sd1511840, -32'sd2057594, -32'sd1252852, -32'sd531273, -32'sd302867, 32'sd210502, -32'sd174897, -32'sd802773, -32'sd1425438, 32'sd182168, 32'sd0, -32'sd349826, 32'sd499274, 32'sd1779186, 32'sd1973288, 32'sd39118, 32'sd1121223, 32'sd2078407, 32'sd938817, 32'sd454212, 32'sd947873, -32'sd66218, 32'sd24096, 32'sd1423790, 32'sd1007531, 32'sd2710974, 32'sd2778910, -32'sd267649, -32'sd1431433, -32'sd3825586, -32'sd592277, -32'sd1740410, 32'sd262120, -32'sd478768, -32'sd372566, -32'sd1044297, 32'sd151669, -32'sd357844, 32'sd0, 32'sd1092147, -32'sd167795, -32'sd389851, -32'sd661296, 32'sd170314, 32'sd583111, 32'sd217805, -32'sd316840, 32'sd1618505, 32'sd1291245, 32'sd271184, 32'sd1585239, 32'sd784510, 32'sd1802512, 32'sd2740119, 32'sd2939374, 32'sd54211, -32'sd497170, -32'sd1945174, -32'sd1633131, 32'sd871547, -32'sd751387, -32'sd589247, -32'sd616268, -32'sd809186, 32'sd541273, -32'sd1057374, -32'sd91018, -32'sd55011, 32'sd420715, 32'sd515148, -32'sd935978, -32'sd275792, -32'sd1075026, 32'sd1381181, -32'sd2589518, -32'sd1347724, 32'sd793868, 32'sd626276, 32'sd1262462, 32'sd1934620, 32'sd568726, -32'sd261236, 32'sd2299974, -32'sd697770, -32'sd3364405, -32'sd2037936, -32'sd2952720, -32'sd2155379, -32'sd2247626, -32'sd2086793, -32'sd849834, 32'sd363642, 32'sd485170, 32'sd28506, 32'sd448677, -32'sd1085956, -32'sd873504, -32'sd490051, 32'sd796081, -32'sd167816, -32'sd2051355, -32'sd479738, -32'sd2602557, -32'sd2066281, -32'sd55403, 32'sd579410, -32'sd253458, 32'sd2128381, 32'sd3444899, 32'sd4428921, 32'sd2481123, 32'sd506751, -32'sd3271643, -32'sd2823328, -32'sd2741187, -32'sd2281581, -32'sd3147867, -32'sd857714, 32'sd1532026, 32'sd675828, 32'sd1349427, -32'sd872262, 32'sd521967, 32'sd1692538, -32'sd705613, -32'sd1410432, 32'sd1335750, -32'sd696299, 32'sd1085182, -32'sd1970706, -32'sd2017447, -32'sd1623281, -32'sd2729341, -32'sd3089507, 32'sd1640822, 32'sd1127949, 32'sd1392359, 32'sd3908450, 32'sd2842629, -32'sd496976, -32'sd2341099, -32'sd2410427, -32'sd2555254, -32'sd3555300, -32'sd1776357, -32'sd1332642, 32'sd1396261, 32'sd1516637, 32'sd1413339, 32'sd18886, 32'sd392945, 32'sd328833, -32'sd1452186, -32'sd2224737, -32'sd798307, -32'sd502460, 32'sd106068, -32'sd2176011, -32'sd1462013, -32'sd2516482, -32'sd1058369, -32'sd1243156, -32'sd513564, 32'sd1668193, 32'sd2368092, 32'sd4019005, 32'sd1002368, -32'sd1710701, -32'sd3330688, -32'sd3065891, -32'sd1922100, -32'sd1421828, -32'sd1470203, -32'sd1968305, -32'sd722690, 32'sd2227993, 32'sd1689608, 32'sd846029, 32'sd5986, 32'sd112231, -32'sd827013, -32'sd1381702, -32'sd484512, 32'sd1498689, -32'sd239726, -32'sd473247, 32'sd1261393, -32'sd638588, -32'sd1323253, 32'sd379104, 32'sd1466707, 32'sd1677838, 32'sd3553429, 32'sd1156048, -32'sd352247, -32'sd1673101, -32'sd2823314, -32'sd596148, -32'sd842392, -32'sd2046330, -32'sd517113, -32'sd901258, -32'sd1569059, -32'sd1046439, 32'sd779034, -32'sd645650, 32'sd342046, -32'sd854191, -32'sd1437698, -32'sd867997, -32'sd827240, 32'sd881858, -32'sd433326, 32'sd428410, 32'sd691085, -32'sd1524821, 32'sd567868, -32'sd1130245, 32'sd520798, 32'sd2812830, 32'sd1032345, -32'sd868205, -32'sd821251, -32'sd2362569, -32'sd1736463, -32'sd2205007, -32'sd2465458, -32'sd1838392, 32'sd919657, -32'sd808130, -32'sd379149, 32'sd454876, -32'sd81407, -32'sd128119, -32'sd61249, -32'sd736789, 32'sd165841, -32'sd1614570, -32'sd2175463, -32'sd310135, 32'sd528907, -32'sd2139599, 32'sd305433, 32'sd250143, 32'sd1881121, 32'sd1664343, 32'sd1077637, 32'sd1036669, 32'sd742926, -32'sd1373589, -32'sd1421398, -32'sd348813, -32'sd1682077, -32'sd45655, -32'sd72039, 32'sd1379122, 32'sd9585, 32'sd564745, -32'sd1010113, -32'sd577888, 32'sd953668, 32'sd699582, -32'sd855400, 32'sd1173540, 32'sd1031993, 32'sd1598847, -32'sd2404058, 32'sd1668578, 32'sd471575, 32'sd1171095, 32'sd248541, -32'sd533531, -32'sd211482, 32'sd1706361, 32'sd774154, 32'sd1197485, 32'sd2882543, -32'sd485235, 32'sd1324435, -32'sd2531537, -32'sd567536, -32'sd729630, -32'sd256245, 32'sd2477359, 32'sd926001, 32'sd1579580, 32'sd604244, 32'sd669179, 32'sd225065, -32'sd736276, 32'sd325373, 32'sd319408, -32'sd1495279, 32'sd2114793, -32'sd1857891, 32'sd96419, 32'sd2179469, 32'sd2205520, 32'sd119998, -32'sd350798, -32'sd827366, 32'sd2546234, 32'sd113317, 32'sd1175057, 32'sd1996615, 32'sd2034718, -32'sd312073, -32'sd2488397, -32'sd1061071, 32'sd904094, 32'sd219835, 32'sd718900, 32'sd3020150, -32'sd1168824, -32'sd919518, -32'sd1025017, -32'sd392419, -32'sd336879, 32'sd921120, -32'sd876875, -32'sd1085611, 32'sd224796, 32'sd821613, 32'sd1109389, 32'sd1172355, 32'sd2835860, 32'sd1496439, -32'sd131179, 32'sd238568, 32'sd1686416, 32'sd1860164, 32'sd544294, 32'sd2315124, 32'sd2442161, 32'sd2507268, -32'sd1097914, -32'sd362807, 32'sd433133, -32'sd173205, 32'sd424192, 32'sd905922, -32'sd272074, -32'sd198107, -32'sd4649882, 32'sd376328, -32'sd105163, 32'sd0, -32'sd57949, -32'sd774374, -32'sd1519973, -32'sd833970, -32'sd376346, 32'sd170444, 32'sd702933, -32'sd444826, -32'sd48834, -32'sd1588607, -32'sd1880361, 32'sd39293, 32'sd3059413, 32'sd3134534, 32'sd1429932, 32'sd2303957, -32'sd619519, -32'sd1277659, -32'sd1060483, 32'sd1755936, 32'sd1803424, 32'sd1031594, 32'sd523657, -32'sd226801, -32'sd945622, 32'sd498316, -32'sd83216, -32'sd613946, -32'sd996190, 32'sd853179, -32'sd377973, 32'sd1249951, -32'sd1206655, -32'sd1876847, -32'sd748335, -32'sd359079, -32'sd1110379, -32'sd713021, -32'sd702053, 32'sd1045880, 32'sd3283493, 32'sd323901, -32'sd1248851, -32'sd746022, -32'sd956820, 32'sd727736, -32'sd1956762, 32'sd1564361, 32'sd1794465, -32'sd99424, -32'sd852890, -32'sd1346682, -32'sd1950859, -32'sd763265, -32'sd1348746, 32'sd226987, 32'sd1006337, -32'sd974718, 32'sd690934, 32'sd1353990, -32'sd2018442, 32'sd300549, 32'sd91093, -32'sd1775799, 32'sd600418, -32'sd1494823, 32'sd1388782, 32'sd709610, 32'sd1142668, -32'sd707576, -32'sd531752, 32'sd372744, -32'sd158241, 32'sd464276, -32'sd842372, 32'sd697345, -32'sd37666, 32'sd1967910, -32'sd252809, -32'sd1773805, -32'sd266422, 32'sd574178, 32'sd168922, 32'sd0, 32'sd667040, -32'sd638811, -32'sd492546, -32'sd492030, -32'sd570922, -32'sd180806, -32'sd716491, -32'sd844170, -32'sd515270, -32'sd1316492, 32'sd1034735, -32'sd48076, 32'sd1844240, 32'sd1166626, -32'sd773002, 32'sd372397, 32'sd279296, 32'sd1178840, 32'sd637984, -32'sd831471, 32'sd174966, 32'sd810272, -32'sd1206630, -32'sd710963, -32'sd884945, 32'sd634468, -32'sd364880, 32'sd353380, -32'sd1468763, -32'sd255777, 32'sd432450, -32'sd833932, 32'sd552052, -32'sd691482, -32'sd1174708, -32'sd684900, 32'sd78022, 32'sd1200375, -32'sd875330, -32'sd173695, -32'sd632287, 32'sd2156149, -32'sd914533, -32'sd206019, 32'sd126734, -32'sd432271, -32'sd791746, -32'sd734398, 32'sd189919, 32'sd766010, 32'sd638103, -32'sd998548, -32'sd235959, 32'sd945606, -32'sd156389, -32'sd1092982, -32'sd317383, -32'sd543608, 32'sd952063, 32'sd418400, 32'sd1050590, -32'sd1320898, -32'sd1338878, 32'sd808590, -32'sd1228328, 32'sd455356, -32'sd1724609, 32'sd305528, -32'sd6345, -32'sd576153, 32'sd166648, -32'sd1011170, -32'sd599271, 32'sd1471973, -32'sd1026494, 32'sd565970, -32'sd1191544, 32'sd1706194, -32'sd1264923, 32'sd536434, -32'sd337181, -32'sd264172, 32'sd6905, 32'sd0, 32'sd405751, 32'sd404194, 32'sd2259384, 32'sd110657, -32'sd885620, -32'sd769334, 32'sd16355, -32'sd686882, 32'sd588975, 32'sd1991504, -32'sd726857, -32'sd1437829, 32'sd1513801, 32'sd899172, 32'sd71435, -32'sd2429647, -32'sd1670577, -32'sd407001, 32'sd681626, -32'sd1595385, -32'sd2015790, -32'sd1619901, 32'sd360686, -32'sd1673939, -32'sd714920, 32'sd1449094, 32'sd0, 32'sd0, 32'sd0, 32'sd1344760, -32'sd197093, 32'sd1206081, -32'sd2748713, 32'sd590145, 32'sd222172, 32'sd251145, 32'sd1311955, 32'sd2660588, 32'sd1629772, -32'sd527925, -32'sd655014, -32'sd568675, 32'sd81516, -32'sd933054, -32'sd959937, -32'sd1003073, 32'sd195815, -32'sd1663780, 32'sd879429, 32'sd1286030, -32'sd715793, 32'sd1133900, -32'sd482371, 32'sd240147, 32'sd0, 32'sd0, 32'sd0, 32'sd185930, 32'sd392582, -32'sd1660651, -32'sd181023, 32'sd263437, 32'sd2379700, 32'sd2629559, 32'sd1120688, 32'sd1678598, 32'sd381635, 32'sd1382629, 32'sd517752, -32'sd1950946, -32'sd1141168, -32'sd164124, -32'sd396439, -32'sd244785, -32'sd1706117, -32'sd2694573, -32'sd1422655, -32'sd676680, 32'sd1753850, -32'sd721004, -32'sd699765, 32'sd67215, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd172495, -32'sd519358, 32'sd399965, 32'sd265637, -32'sd1351943, -32'sd697804, 32'sd117139, 32'sd328684, -32'sd113505, -32'sd447968, 32'sd662769, -32'sd180628, -32'sd1917471, -32'sd719515, -32'sd282669, -32'sd174442, -32'sd864710, -32'sd1743481, -32'sd208969, -32'sd44301, -32'sd760516, 32'sd65030, 32'sd638967, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd104536, 32'sd217703, -32'sd142380, 32'sd1027761, 32'sd798742, 32'sd1091759, -32'sd1580088, -32'sd168792, -32'sd1259372, -32'sd1348287, -32'sd2329184, 32'sd412572, 32'sd404377, -32'sd388705, -32'sd668091, -32'sd1420807, 32'sd168248, 32'sd56658, 32'sd81356, 32'sd1744031, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1438666, 32'sd1787818, -32'sd1130436, 32'sd1137633, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd797460, 32'sd559345, 32'sd27225, -32'sd1943501, -32'sd1128570, -32'sd1381152, -32'sd8743, -32'sd875733, 32'sd1496664, 32'sd785843, -32'sd202069, 32'sd338212, -32'sd529598, 32'sd1013984, 32'sd564148, 32'sd906699, 32'sd297715, 32'sd1752530, 32'sd990643, 32'sd118421, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1475372, -32'sd689085, 32'sd1376168, 32'sd357550, -32'sd1850272, -32'sd952722, -32'sd696506, 32'sd785399, -32'sd1194521, 32'sd1305331, 32'sd1716385, 32'sd1449679, 32'sd275149, 32'sd3088232, 32'sd2507514, 32'sd671477, 32'sd996984, -32'sd411471, -32'sd288700, 32'sd289826, -32'sd268031, -32'sd439683, 32'sd2286645, 32'sd1082027, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd518002, 32'sd1572481, -32'sd234944, -32'sd24726, -32'sd1315003, -32'sd1170604, 32'sd656672, -32'sd546653, 32'sd778180, 32'sd542792, -32'sd286477, 32'sd1276743, 32'sd787257, 32'sd1531525, 32'sd1579637, 32'sd2469141, 32'sd1158729, 32'sd3442439, -32'sd104431, -32'sd684431, -32'sd1160266, -32'sd387300, 32'sd12423, -32'sd348018, 32'sd712144, 32'sd0, 32'sd0, 32'sd1039914, 32'sd1243093, -32'sd391312, 32'sd1090787, -32'sd59632, -32'sd2709349, -32'sd732720, 32'sd23725, -32'sd374259, -32'sd270379, -32'sd980641, 32'sd1195308, 32'sd582222, 32'sd1269132, -32'sd491752, -32'sd1213791, -32'sd347965, 32'sd1642408, -32'sd251439, -32'sd829240, 32'sd1633459, 32'sd781336, 32'sd328218, 32'sd701048, -32'sd1153980, -32'sd1063585, -32'sd872940, 32'sd0, 32'sd1344593, -32'sd405599, -32'sd570146, 32'sd402680, 32'sd95368, -32'sd1447986, -32'sd34715, 32'sd293795, 32'sd241174, 32'sd236601, 32'sd182013, -32'sd1220229, 32'sd858287, 32'sd1768458, 32'sd1152533, 32'sd1590241, -32'sd194161, 32'sd984140, -32'sd788113, -32'sd604117, -32'sd467693, -32'sd1343412, 32'sd576160, -32'sd175631, 32'sd498807, 32'sd746921, 32'sd1240650, 32'sd0, 32'sd1110871, -32'sd174263, -32'sd1218592, 32'sd290509, 32'sd7480, -32'sd1825605, -32'sd2366067, -32'sd3713348, -32'sd688413, -32'sd1615657, 32'sd180430, 32'sd890920, 32'sd818553, 32'sd393446, 32'sd68100, -32'sd809649, -32'sd856151, 32'sd1436122, 32'sd76754, 32'sd201682, 32'sd1051724, -32'sd1419137, -32'sd211545, -32'sd668124, -32'sd110692, 32'sd1735557, -32'sd284993, 32'sd680519, -32'sd722558, 32'sd1120541, -32'sd213914, -32'sd645169, -32'sd1666165, -32'sd1546863, -32'sd126403, -32'sd2737177, -32'sd623749, -32'sd366778, -32'sd973366, 32'sd575806, -32'sd147440, 32'sd1350636, -32'sd2218288, -32'sd568708, -32'sd39605, -32'sd1292333, -32'sd735648, -32'sd268253, 32'sd573756, 32'sd293497, -32'sd683349, -32'sd1736742, -32'sd1149291, 32'sd1798985, 32'sd49653, 32'sd1064830, -32'sd118158, -32'sd1310310, 32'sd1030123, 32'sd525978, -32'sd575206, 32'sd100806, 32'sd483433, -32'sd1711018, -32'sd852696, -32'sd1971842, -32'sd2769167, -32'sd1008784, -32'sd424718, 32'sd1133708, -32'sd835626, -32'sd2223970, 32'sd786194, -32'sd2772406, -32'sd701901, -32'sd1586281, -32'sd2000407, -32'sd1974010, -32'sd510609, -32'sd950532, -32'sd1967468, 32'sd1698821, -32'sd358557, 32'sd1841346, -32'sd176428, -32'sd478743, -32'sd400859, 32'sd1760924, 32'sd243167, 32'sd850990, 32'sd1382374, -32'sd613931, -32'sd2553531, -32'sd4335595, -32'sd2796066, 32'sd504618, 32'sd1330257, 32'sd1412805, 32'sd927627, 32'sd720075, -32'sd1056815, -32'sd2290770, -32'sd1231800, -32'sd1597192, -32'sd2620086, -32'sd2038745, -32'sd1388850, -32'sd647865, -32'sd1235635, 32'sd1533535, 32'sd602524, 32'sd144823, 32'sd1913240, -32'sd1740179, -32'sd1134922, 32'sd307875, -32'sd198530, 32'sd1847283, -32'sd199476, -32'sd1366792, -32'sd1192376, -32'sd2141357, -32'sd1623399, 32'sd576552, 32'sd2868941, 32'sd2919904, 32'sd2262540, 32'sd1039595, -32'sd21935, -32'sd568943, -32'sd1935825, -32'sd1854551, -32'sd838482, -32'sd1482725, -32'sd2885876, -32'sd243879, -32'sd1599938, 32'sd1377447, -32'sd265627, 32'sd188958, 32'sd44031, -32'sd3057153, -32'sd1613475, 32'sd949010, 32'sd219450, -32'sd137547, 32'sd566266, -32'sd1755557, -32'sd2783203, -32'sd2557568, -32'sd36923, 32'sd2316090, 32'sd2123468, 32'sd2613141, 32'sd2205025, -32'sd1821157, -32'sd2174095, -32'sd1424144, 32'sd748890, -32'sd1066197, -32'sd1172656, -32'sd1381818, -32'sd2028011, -32'sd3181039, 32'sd207204, 32'sd1216033, -32'sd369945, 32'sd458390, -32'sd1450624, 32'sd705149, 32'sd435047, 32'sd1175227, 32'sd256659, -32'sd1549202, -32'sd2470792, -32'sd3474976, -32'sd953917, 32'sd1712020, 32'sd801710, 32'sd2962819, 32'sd2388134, 32'sd1285535, 32'sd2380576, -32'sd1051062, -32'sd565064, 32'sd317413, 32'sd1322344, -32'sd726428, 32'sd899853, -32'sd1451378, 32'sd1348824, -32'sd288267, -32'sd1536692, -32'sd1399186, -32'sd1760665, 32'sd243236, -32'sd45406, -32'sd271661, 32'sd1090308, 32'sd68771, 32'sd1705968, 32'sd205038, 32'sd69586, -32'sd836060, 32'sd761358, 32'sd2679050, 32'sd1015581, -32'sd369085, -32'sd533805, 32'sd475283, 32'sd1264236, 32'sd162015, 32'sd878850, 32'sd351311, 32'sd2036511, 32'sd1942343, 32'sd1593398, -32'sd129412, 32'sd2126155, 32'sd125753, -32'sd1734220, -32'sd628169, 32'sd79678, 32'sd1929249, -32'sd188270, 32'sd241696, 32'sd811836, -32'sd353816, -32'sd203741, 32'sd901762, -32'sd1947199, -32'sd719084, -32'sd349501, 32'sd2804881, 32'sd1300088, 32'sd904711, 32'sd670294, 32'sd1013691, -32'sd1374834, 32'sd683881, -32'sd82156, 32'sd1164733, 32'sd3085974, 32'sd596875, 32'sd2717949, 32'sd1547655, 32'sd2286327, -32'sd102858, -32'sd728272, -32'sd2351853, 32'sd266038, 32'sd1567981, -32'sd1125810, -32'sd466809, -32'sd694099, -32'sd535330, 32'sd17111, 32'sd1783991, 32'sd1560022, -32'sd79182, 32'sd203140, 32'sd1855937, 32'sd726292, 32'sd97295, -32'sd400550, 32'sd276162, -32'sd740993, -32'sd585159, 32'sd1090213, 32'sd2620836, 32'sd2919183, 32'sd1489649, 32'sd1075795, 32'sd1779846, 32'sd2853953, 32'sd761151, -32'sd618466, -32'sd215056, 32'sd220427, -32'sd371335, 32'sd115248, 32'sd603832, -32'sd659599, -32'sd630180, -32'sd1433975, 32'sd580155, 32'sd2608756, 32'sd1500345, 32'sd963541, 32'sd1594071, 32'sd1328325, 32'sd766696, 32'sd849058, -32'sd244208, -32'sd715509, 32'sd676888, -32'sd923384, 32'sd2046827, 32'sd1790692, 32'sd128525, 32'sd2569423, 32'sd115359, 32'sd721367, 32'sd1232209, -32'sd2922772, 32'sd812810, 32'sd825155, 32'sd0, 32'sd759326, -32'sd326595, 32'sd126822, 32'sd2780618, 32'sd690577, 32'sd127082, 32'sd1491052, -32'sd169003, -32'sd1069510, 32'sd818716, -32'sd1096702, -32'sd998917, 32'sd255681, 32'sd688548, -32'sd2044083, 32'sd1833163, 32'sd280454, -32'sd760046, -32'sd10579, 32'sd890968, 32'sd1824653, 32'sd303366, 32'sd1003257, 32'sd593454, -32'sd1042946, 32'sd1387074, -32'sd1656652, -32'sd656952, 32'sd568573, -32'sd1288908, 32'sd1159944, 32'sd1191431, -32'sd148206, 32'sd5808, 32'sd912689, -32'sd1529988, -32'sd158281, -32'sd720424, -32'sd1621704, -32'sd1711381, 32'sd2775240, 32'sd656154, 32'sd177776, -32'sd719363, -32'sd515370, -32'sd199750, 32'sd324966, -32'sd977209, -32'sd204820, 32'sd582123, -32'sd1979376, -32'sd601794, -32'sd496173, 32'sd1419491, -32'sd201652, 32'sd371987, 32'sd420591, -32'sd763238, -32'sd305361, 32'sd269612, 32'sd269921, 32'sd125782, -32'sd848115, -32'sd2312896, 32'sd2095858, -32'sd1697408, -32'sd982164, 32'sd2281421, 32'sd904421, -32'sd261512, 32'sd602833, -32'sd428199, -32'sd615459, 32'sd817812, 32'sd87488, -32'sd1508258, -32'sd1095069, -32'sd2115564, -32'sd1510060, -32'sd1508195, -32'sd2219177, -32'sd655825, -32'sd471423, 32'sd0, -32'sd720031, 32'sd206431, -32'sd371363, -32'sd41584, -32'sd28201, -32'sd423371, -32'sd105101, -32'sd1729106, -32'sd880961, -32'sd207553, 32'sd710210, 32'sd174550, 32'sd2664335, 32'sd1668604, 32'sd1556797, 32'sd2193760, -32'sd2141140, 32'sd913009, -32'sd2160546, -32'sd159224, -32'sd1278204, -32'sd1363014, -32'sd2465898, -32'sd1389666, -32'sd1937425, 32'sd1083348, -32'sd362810, 32'sd1296888, 32'sd1160566, 32'sd896854, -32'sd1849336, -32'sd1632992, -32'sd1743417, -32'sd800451, -32'sd1171587, -32'sd638809, -32'sd1244278, -32'sd264377, -32'sd27737, 32'sd583114, 32'sd199802, 32'sd1619495, 32'sd1560499, 32'sd1941518, 32'sd233386, 32'sd1325894, -32'sd242072, -32'sd1623447, -32'sd2827284, -32'sd1577219, -32'sd1076712, 32'sd258625, 32'sd129855, 32'sd1000898, 32'sd123904, -32'sd22875, 32'sd1515630, 32'sd1147554, -32'sd553946, -32'sd1289787, 32'sd843978, -32'sd1630141, -32'sd1910329, -32'sd1292921, -32'sd2120322, -32'sd31563, 32'sd127941, 32'sd336199, 32'sd95608, -32'sd789201, 32'sd73055, 32'sd711170, -32'sd1030199, -32'sd951070, -32'sd909192, -32'sd347804, -32'sd1078092, 32'sd902543, -32'sd1219282, -32'sd1724427, -32'sd722493, 32'sd807943, 32'sd446836, 32'sd0, 32'sd1411863, 32'sd155158, 32'sd1409851, 32'sd1497693, 32'sd880986, 32'sd438050, 32'sd648842, 32'sd595967, 32'sd1176709, 32'sd1281675, 32'sd2473005, 32'sd854918, 32'sd50625, 32'sd734751, 32'sd1691542, -32'sd1251017, -32'sd1255273, -32'sd1511141, 32'sd456722, -32'sd192434, 32'sd466741, 32'sd708692, -32'sd806648, -32'sd955060, 32'sd938990, -32'sd1163186, 32'sd0, 32'sd0, 32'sd0, -32'sd126848, -32'sd1195312, -32'sd727392, -32'sd618063, -32'sd1302424, 32'sd801357, -32'sd1443882, 32'sd2068914, -32'sd30084, 32'sd4115, -32'sd708672, -32'sd657929, 32'sd1451509, -32'sd402922, -32'sd854216, -32'sd1139356, -32'sd635921, 32'sd299918, 32'sd621870, -32'sd1635210, -32'sd1402735, 32'sd808371, 32'sd1119370, 32'sd440361, 32'sd578669, 32'sd0, 32'sd0, 32'sd0, 32'sd146726, 32'sd472589, 32'sd1687108, 32'sd1026214, 32'sd1482116, 32'sd1194887, -32'sd377148, 32'sd808531, 32'sd529881, 32'sd1154162, 32'sd462179, 32'sd1004045, -32'sd1864442, 32'sd81209, 32'sd1252041, -32'sd2009264, -32'sd397090, -32'sd1606867, -32'sd1553977, -32'sd2697808, -32'sd1938358, 32'sd298721, 32'sd513726, 32'sd431875, 32'sd1240126, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd308948, -32'sd2036044, -32'sd1675781, -32'sd368817, -32'sd1612649, -32'sd3121018, -32'sd1589651, -32'sd125658, 32'sd328142, -32'sd522110, 32'sd1611024, 32'sd785861, 32'sd1507552, 32'sd807200, -32'sd769201, -32'sd83208, -32'sd381656, -32'sd1035511, -32'sd1494338, -32'sd336952, -32'sd585230, 32'sd467219, 32'sd1137268, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1711449, 32'sd982430, 32'sd27621, 32'sd976036, -32'sd792293, 32'sd1186042, -32'sd830814, 32'sd289545, 32'sd461932, -32'sd457342, 32'sd1589503, -32'sd361184, 32'sd109537, 32'sd61468, -32'sd226016, -32'sd1549397, 32'sd871939, -32'sd856179, 32'sd419785, 32'sd39318, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd503793, -32'sd244924, 32'sd547700, 32'sd644936, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd240084, -32'sd602276, -32'sd935471, 32'sd274400, 32'sd67559, -32'sd948885, 32'sd801806, 32'sd527428, -32'sd1710221, -32'sd870541, -32'sd611825, -32'sd989904, 32'sd1087267, -32'sd323211, -32'sd331578, 32'sd1064532, -32'sd677265, 32'sd254014, 32'sd365319, 32'sd522954, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd266892, 32'sd766322, -32'sd79286, 32'sd135517, 32'sd1185603, -32'sd680231, 32'sd327259, -32'sd66231, 32'sd228315, 32'sd1250079, -32'sd198949, -32'sd874617, -32'sd1103793, 32'sd129499, 32'sd1136110, 32'sd487819, 32'sd1919797, 32'sd446288, 32'sd257631, -32'sd262487, 32'sd1277147, 32'sd195161, 32'sd233051, 32'sd667324, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1071148, 32'sd577536, 32'sd409835, 32'sd538674, 32'sd1124098, 32'sd977312, 32'sd1166459, 32'sd651870, 32'sd1706664, 32'sd1122447, 32'sd3184409, 32'sd2118261, 32'sd1395910, 32'sd1458163, 32'sd2364549, -32'sd94750, -32'sd1010367, 32'sd283052, 32'sd21859, -32'sd1344490, 32'sd327375, 32'sd1117255, -32'sd434975, 32'sd128022, -32'sd106572, 32'sd0, 32'sd0, 32'sd683851, -32'sd1325428, 32'sd29037, -32'sd1511451, -32'sd623985, 32'sd385924, 32'sd857941, 32'sd989893, 32'sd118244, -32'sd1446142, 32'sd341253, 32'sd921637, 32'sd2545768, 32'sd1694475, 32'sd2888856, 32'sd1143994, 32'sd72957, -32'sd1167727, 32'sd1533086, 32'sd1864888, -32'sd42882, 32'sd661089, 32'sd1354133, -32'sd60038, 32'sd840381, 32'sd1011450, -32'sd656272, 32'sd0, 32'sd622729, 32'sd834907, -32'sd1753312, 32'sd240855, -32'sd726620, -32'sd931233, -32'sd1327711, -32'sd574813, -32'sd217017, -32'sd1062550, 32'sd2847485, 32'sd1893992, 32'sd602321, 32'sd225491, 32'sd787785, 32'sd1404558, 32'sd487965, 32'sd667381, 32'sd1125265, 32'sd334989, -32'sd50515, -32'sd790361, 32'sd862011, -32'sd527962, -32'sd995384, 32'sd1152464, 32'sd1554977, 32'sd0, 32'sd1309690, -32'sd73953, 32'sd1078617, 32'sd688070, -32'sd1117777, 32'sd529910, -32'sd1374691, -32'sd477818, 32'sd2551154, -32'sd383408, 32'sd725135, -32'sd48006, 32'sd1338651, 32'sd53986, -32'sd78741, 32'sd1190374, 32'sd480559, 32'sd1149019, -32'sd1113286, -32'sd2514586, 32'sd147171, -32'sd1704592, 32'sd138798, 32'sd1566465, 32'sd1309396, 32'sd1138825, 32'sd103134, 32'sd256017, -32'sd378588, 32'sd920546, -32'sd543275, 32'sd1102518, 32'sd143290, 32'sd352476, -32'sd520849, 32'sd485096, 32'sd561564, 32'sd824307, 32'sd4321727, 32'sd1637186, 32'sd1334710, -32'sd52677, 32'sd1466851, 32'sd1721488, -32'sd71497, 32'sd141456, -32'sd11994, -32'sd463174, -32'sd793530, -32'sd750874, -32'sd1280608, 32'sd710853, 32'sd2144819, -32'sd758639, -32'sd798579, 32'sd539273, 32'sd641464, -32'sd1858482, -32'sd705077, -32'sd43791, -32'sd527889, -32'sd797153, 32'sd1288608, 32'sd3715402, 32'sd1226232, 32'sd150360, 32'sd1554666, 32'sd320447, 32'sd189851, -32'sd607807, -32'sd2182453, -32'sd2822508, -32'sd2031016, -32'sd1234831, 32'sd560176, -32'sd507470, 32'sd85261, -32'sd1076921, -32'sd18805, -32'sd1559438, 32'sd1221932, 32'sd899312, 32'sd866763, -32'sd885602, -32'sd633618, 32'sd109835, -32'sd1259220, 32'sd119649, 32'sd1519493, 32'sd1012010, 32'sd1033552, 32'sd2087574, 32'sd1647076, 32'sd610280, 32'sd568746, 32'sd116869, -32'sd461757, -32'sd1308158, -32'sd191609, -32'sd438053, -32'sd1394428, -32'sd618703, -32'sd1283631, -32'sd1030181, -32'sd606293, 32'sd734872, -32'sd388184, -32'sd2060955, -32'sd1339602, 32'sd339648, -32'sd1505308, 32'sd115044, -32'sd2299999, -32'sd493148, 32'sd1079543, 32'sd1388779, 32'sd297265, 32'sd844577, 32'sd181324, -32'sd2077600, -32'sd99199, 32'sd806658, -32'sd1247554, 32'sd780201, 32'sd950882, 32'sd1071405, -32'sd283113, 32'sd993303, 32'sd358184, -32'sd650137, 32'sd465158, -32'sd1400217, -32'sd1131907, -32'sd940112, -32'sd1011027, 32'sd839390, 32'sd70517, -32'sd733836, 32'sd945448, -32'sd394478, 32'sd673270, -32'sd158328, 32'sd343776, 32'sd478050, 32'sd194746, 32'sd69033, -32'sd276745, -32'sd2504965, -32'sd3126907, 32'sd1373475, 32'sd2228112, 32'sd1379131, 32'sd1259743, 32'sd1910862, -32'sd43806, 32'sd2128520, -32'sd238919, -32'sd1683779, -32'sd2143281, -32'sd2846078, -32'sd1132891, -32'sd1559994, -32'sd821451, -32'sd174137, -32'sd445596, -32'sd623305, 32'sd1717206, 32'sd656774, -32'sd1210925, -32'sd335373, -32'sd968888, 32'sd1050227, -32'sd491397, -32'sd2348216, -32'sd1244699, -32'sd1066167, -32'sd345284, 32'sd403731, -32'sd301397, 32'sd571996, 32'sd1063022, 32'sd717398, 32'sd387751, -32'sd84464, 32'sd240962, -32'sd170158, -32'sd180039, 32'sd1641289, 32'sd1140288, -32'sd1350991, -32'sd269221, -32'sd1000995, -32'sd617758, -32'sd800810, 32'sd2283, 32'sd657450, 32'sd869181, -32'sd90268, -32'sd355685, 32'sd4056, 32'sd707469, -32'sd2274857, -32'sd1329369, -32'sd2308452, -32'sd1014692, -32'sd1138406, 32'sd237585, 32'sd475583, -32'sd191425, -32'sd897559, -32'sd3338816, -32'sd1393844, 32'sd206399, 32'sd1507855, 32'sd1979162, 32'sd2599361, 32'sd3117088, -32'sd613416, 32'sd445819, 32'sd791701, 32'sd665224, -32'sd522813, 32'sd1146470, 32'sd1080044, -32'sd383749, -32'sd1336490, 32'sd997344, -32'sd3411448, -32'sd1473157, -32'sd2075049, -32'sd923600, -32'sd3568937, -32'sd2927777, -32'sd4594297, -32'sd2479323, -32'sd1041278, 32'sd152968, 32'sd395770, -32'sd747830, 32'sd780529, -32'sd1994472, 32'sd1133435, -32'sd104380, 32'sd1311684, 32'sd583838, 32'sd239949, 32'sd507048, -32'sd1728839, -32'sd436975, -32'sd463288, 32'sd1862488, 32'sd1756714, 32'sd1115274, 32'sd1735079, -32'sd549756, -32'sd3432963, -32'sd2892287, -32'sd3415260, -32'sd3004153, -32'sd3705206, -32'sd5854100, -32'sd3795718, -32'sd3613857, -32'sd1354342, -32'sd911148, 32'sd2535182, 32'sd1996887, 32'sd1218778, 32'sd613699, -32'sd999849, 32'sd843382, 32'sd661309, 32'sd270656, 32'sd316498, 32'sd685182, -32'sd1177193, -32'sd545889, -32'sd256159, 32'sd696363, 32'sd614310, -32'sd1255837, 32'sd471349, 32'sd827785, -32'sd1898767, -32'sd1419939, -32'sd3579228, -32'sd4097529, -32'sd6083522, -32'sd4961425, -32'sd3438496, -32'sd5383277, -32'sd2304464, 32'sd315862, 32'sd2051727, 32'sd1972150, 32'sd255296, 32'sd1238448, -32'sd522072, 32'sd817297, 32'sd134054, 32'sd1158199, 32'sd1659265, -32'sd350859, -32'sd995263, 32'sd1754080, 32'sd824400, -32'sd582959, 32'sd0, 32'sd747014, -32'sd801916, -32'sd728750, -32'sd2615871, -32'sd202301, -32'sd2702797, -32'sd3199701, -32'sd1959167, -32'sd4211921, -32'sd4085740, -32'sd4168593, -32'sd4524743, -32'sd128910, 32'sd544201, 32'sd709845, -32'sd1914608, 32'sd149140, 32'sd522033, -32'sd1228141, 32'sd331636, 32'sd949753, -32'sd1220377, -32'sd1595269, -32'sd701916, 32'sd2470181, 32'sd1260723, 32'sd917548, -32'sd173749, 32'sd1193280, 32'sd1453483, 32'sd1490236, -32'sd56553, -32'sd172781, -32'sd1170494, -32'sd2128790, -32'sd1386649, -32'sd2051744, -32'sd1793650, -32'sd2331356, -32'sd3541437, -32'sd507298, -32'sd1012487, 32'sd419786, 32'sd1441928, 32'sd466238, -32'sd524732, 32'sd252654, -32'sd1006257, 32'sd648137, -32'sd313712, 32'sd751190, -32'sd1310016, 32'sd451232, -32'sd943, -32'sd766301, 32'sd436919, -32'sd341173, 32'sd102279, 32'sd1268320, -32'sd126861, -32'sd21719, 32'sd806353, -32'sd229168, 32'sd291188, -32'sd988047, 32'sd2371093, 32'sd895053, -32'sd1431927, -32'sd127751, -32'sd1145379, -32'sd898190, 32'sd2415799, 32'sd922901, -32'sd993007, -32'sd271794, -32'sd513731, -32'sd2063003, 32'sd184246, 32'sd730031, -32'sd826119, -32'sd548198, 32'sd1536102, 32'sd278535, 32'sd0, 32'sd820745, 32'sd581266, -32'sd1360153, 32'sd228727, 32'sd804357, 32'sd2104863, 32'sd802774, 32'sd2480936, 32'sd1571974, 32'sd3421326, 32'sd3192728, 32'sd3077351, 32'sd2401921, -32'sd926373, -32'sd279128, 32'sd2765264, 32'sd550866, 32'sd78786, -32'sd416171, -32'sd843908, 32'sd448464, 32'sd942030, -32'sd1275778, 32'sd480775, 32'sd151875, 32'sd1774902, -32'sd505950, 32'sd1658766, -32'sd129399, 32'sd822425, -32'sd917022, 32'sd1010689, 32'sd1448876, 32'sd814844, 32'sd1430383, 32'sd1798528, 32'sd3160771, 32'sd4510244, 32'sd4277277, 32'sd3889956, 32'sd3900080, -32'sd130830, -32'sd99641, 32'sd1645084, 32'sd2460312, 32'sd2329428, 32'sd389902, 32'sd2620143, 32'sd1091136, -32'sd865334, 32'sd1564668, 32'sd2222733, -32'sd245857, -32'sd493127, 32'sd513582, 32'sd873453, 32'sd668779, -32'sd154493, 32'sd1525770, 32'sd1059334, -32'sd1356886, 32'sd587689, 32'sd2232880, 32'sd2170845, 32'sd1936876, 32'sd2174929, 32'sd1524641, 32'sd2119592, 32'sd2689702, 32'sd2628704, 32'sd3050548, 32'sd1618713, 32'sd771714, 32'sd1973826, -32'sd701561, 32'sd1616411, 32'sd693112, 32'sd1221221, 32'sd3330751, 32'sd250874, 32'sd1940388, 32'sd532232, 32'sd927806, 32'sd0, 32'sd1327751, 32'sd1783437, 32'sd795193, -32'sd277545, -32'sd996190, 32'sd485282, -32'sd334146, 32'sd2555154, 32'sd1886236, 32'sd1976523, 32'sd3019101, 32'sd2242692, 32'sd2601159, 32'sd2311819, 32'sd2572857, 32'sd2295864, -32'sd644520, -32'sd525324, 32'sd958844, -32'sd284156, 32'sd1764669, 32'sd1372232, 32'sd615932, -32'sd511535, -32'sd1332892, -32'sd598190, 32'sd0, 32'sd0, 32'sd0, -32'sd434970, -32'sd2270667, -32'sd2511075, -32'sd12746, 32'sd1553239, 32'sd1213794, -32'sd706754, -32'sd1329409, -32'sd613611, 32'sd379355, -32'sd554281, -32'sd525122, 32'sd2337540, -32'sd1105698, 32'sd890415, 32'sd400824, 32'sd1908143, 32'sd1987334, -32'sd460147, 32'sd923148, 32'sd72192, 32'sd772455, 32'sd950679, -32'sd428621, 32'sd267191, 32'sd0, 32'sd0, 32'sd0, -32'sd14809, 32'sd1138465, -32'sd1807958, -32'sd1801863, 32'sd1030091, -32'sd517699, -32'sd978472, -32'sd1368004, -32'sd804363, 32'sd355320, 32'sd1223361, 32'sd1988755, 32'sd2359169, 32'sd826980, -32'sd552569, 32'sd944759, -32'sd1117752, 32'sd250001, 32'sd154031, -32'sd1598237, -32'sd1549048, -32'sd1345876, 32'sd781706, -32'sd33501, 32'sd1278610, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1329983, 32'sd491381, -32'sd470426, -32'sd472672, 32'sd1056802, 32'sd947181, -32'sd875410, -32'sd777476, 32'sd994384, -32'sd323105, 32'sd200061, -32'sd1464434, -32'sd1659788, -32'sd884835, 32'sd330590, -32'sd359788, -32'sd1604129, -32'sd603883, -32'sd20199, 32'sd769731, -32'sd199690, 32'sd615753, -32'sd568833, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd218719, 32'sd732338, 32'sd1746, 32'sd1244041, 32'sd1554522, 32'sd1430936, -32'sd344062, -32'sd164587, 32'sd965666, -32'sd528599, 32'sd1029224, -32'sd538051, 32'sd1282126, 32'sd104728, 32'sd244760, 32'sd558542, -32'sd909840, 32'sd254482, -32'sd205469, 32'sd538175, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd26620, -32'sd1134394, -32'sd722416, 32'sd408928, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd13652, 32'sd52377, 32'sd179987, -32'sd848714, -32'sd689825, -32'sd879185, -32'sd1527266, -32'sd1581028, -32'sd1463415, -32'sd269335, 32'sd290011, -32'sd122755, 32'sd245244, -32'sd1758186, 32'sd633542, -32'sd1171330, 32'sd572191, 32'sd1151393, -32'sd418759, -32'sd1112670, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd44846, -32'sd83766, -32'sd1497043, -32'sd810756, -32'sd385222, -32'sd1141228, -32'sd791546, 32'sd490049, 32'sd698997, 32'sd224832, 32'sd2093665, -32'sd1279576, -32'sd560667, 32'sd378968, -32'sd1776808, 32'sd348639, -32'sd263799, -32'sd256780, -32'sd799415, 32'sd1253808, 32'sd1100126, -32'sd1495578, -32'sd163929, -32'sd1226560, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd226211, -32'sd900962, -32'sd1407742, -32'sd1313108, -32'sd1799997, -32'sd2339393, -32'sd761792, 32'sd73062, 32'sd437765, 32'sd418775, -32'sd252289, 32'sd897051, 32'sd2241568, 32'sd712198, 32'sd477856, -32'sd983498, -32'sd97160, -32'sd33118, -32'sd1234188, 32'sd2012327, -32'sd767255, 32'sd221492, 32'sd814674, 32'sd91698, -32'sd320771, 32'sd0, 32'sd0, 32'sd271928, -32'sd1300212, -32'sd125101, -32'sd1843589, -32'sd313090, -32'sd296976, 32'sd623392, -32'sd317679, 32'sd2226950, 32'sd334487, -32'sd464848, -32'sd1422777, 32'sd827602, 32'sd328670, 32'sd1370834, 32'sd810841, 32'sd2284580, 32'sd856553, -32'sd459866, 32'sd1332126, 32'sd1827918, 32'sd1587175, -32'sd423112, 32'sd1613582, -32'sd516315, -32'sd5626, 32'sd343491, 32'sd0, 32'sd559846, -32'sd281230, -32'sd307298, -32'sd1434919, -32'sd807297, 32'sd1516242, -32'sd273950, -32'sd462722, -32'sd703100, -32'sd1098613, -32'sd950023, 32'sd1551970, 32'sd2645624, 32'sd1348889, 32'sd1380712, 32'sd1552058, 32'sd1678068, 32'sd282479, 32'sd1629980, 32'sd2706149, 32'sd1879253, 32'sd468873, 32'sd191163, 32'sd597967, 32'sd127038, 32'sd216860, 32'sd214731, 32'sd0, 32'sd390451, 32'sd1236357, -32'sd884939, -32'sd1099488, 32'sd309691, 32'sd175879, -32'sd1343699, 32'sd161501, -32'sd154019, -32'sd259940, 32'sd628949, 32'sd1177662, 32'sd532322, 32'sd796207, -32'sd2188283, -32'sd419172, 32'sd836642, -32'sd120851, 32'sd1642240, -32'sd474356, -32'sd131320, 32'sd2351719, -32'sd250419, 32'sd466168, 32'sd1020868, 32'sd522640, -32'sd7344, 32'sd246120, 32'sd401124, 32'sd1300645, 32'sd1556656, 32'sd433513, -32'sd1766935, -32'sd43304, 32'sd744306, -32'sd347571, 32'sd1336575, 32'sd861955, -32'sd1110813, 32'sd1128136, 32'sd942123, -32'sd1807339, 32'sd198550, -32'sd2089401, -32'sd916120, 32'sd1803073, -32'sd1660463, -32'sd561961, -32'sd865308, -32'sd638148, 32'sd716413, 32'sd569917, 32'sd1272070, -32'sd450366, 32'sd974477, 32'sd92796, 32'sd757786, -32'sd477080, -32'sd1117385, 32'sd873928, -32'sd639757, 32'sd758503, -32'sd710113, -32'sd1224549, 32'sd665852, 32'sd68667, -32'sd901166, -32'sd436475, 32'sd1605727, -32'sd109192, -32'sd1450464, -32'sd1351819, -32'sd1474875, 32'sd1641683, 32'sd960243, 32'sd164062, 32'sd563768, 32'sd224903, 32'sd708311, -32'sd757938, 32'sd456705, 32'sd605695, 32'sd278338, -32'sd1018882, -32'sd1306278, -32'sd2071458, -32'sd519506, 32'sd1497145, 32'sd1017909, -32'sd703045, -32'sd548251, -32'sd191544, 32'sd19351, -32'sd1707717, -32'sd667824, -32'sd657378, 32'sd704588, -32'sd390448, -32'sd2356444, -32'sd4137386, -32'sd1000362, 32'sd1137798, 32'sd2537958, 32'sd1539364, 32'sd1844098, 32'sd1637405, 32'sd2098694, -32'sd346754, 32'sd1079056, 32'sd718271, 32'sd767672, -32'sd1366994, -32'sd779944, 32'sd86352, 32'sd1938916, -32'sd1244949, 32'sd65367, 32'sd1014814, 32'sd109869, 32'sd966845, -32'sd1225030, -32'sd1835920, -32'sd1774204, -32'sd1235078, 32'sd652811, 32'sd3850838, 32'sd405842, -32'sd1117728, -32'sd2218191, 32'sd1377718, 32'sd733339, 32'sd2877381, 32'sd3027634, 32'sd1602637, 32'sd1058207, -32'sd3454673, -32'sd2680535, -32'sd789819, 32'sd428364, -32'sd721978, -32'sd77276, 32'sd1677436, 32'sd271940, -32'sd1182698, -32'sd441967, 32'sd956008, 32'sd1367518, -32'sd19559, -32'sd2826577, -32'sd1191035, -32'sd3304830, 32'sd681080, 32'sd2050462, 32'sd4244923, 32'sd3015552, -32'sd170169, -32'sd54296, 32'sd1438062, 32'sd3069249, 32'sd2663253, 32'sd872873, 32'sd1802625, 32'sd209666, -32'sd1875713, -32'sd792621, 32'sd141273, 32'sd50407, 32'sd820240, 32'sd1369390, 32'sd592356, -32'sd307472, -32'sd1266977, 32'sd1177731, 32'sd68274, -32'sd2332198, -32'sd2903467, -32'sd3158904, -32'sd2526356, -32'sd71934, 32'sd1285337, 32'sd2903747, 32'sd4896903, 32'sd4128871, 32'sd1094936, 32'sd2396218, 32'sd854051, 32'sd1301138, -32'sd312656, -32'sd439064, -32'sd593144, -32'sd2404564, -32'sd693547, -32'sd1366207, -32'sd18499, -32'sd1277707, -32'sd1066382, 32'sd769677, 32'sd668336, -32'sd1200660, -32'sd2070483, -32'sd1546790, -32'sd1817250, -32'sd1767437, -32'sd491398, -32'sd2241152, 32'sd283065, 32'sd3712676, 32'sd4040738, 32'sd3263496, 32'sd3974519, 32'sd1773060, 32'sd1045960, 32'sd1286810, 32'sd368061, -32'sd1691891, -32'sd2083288, -32'sd1349460, -32'sd1094010, -32'sd2783341, -32'sd2478824, -32'sd178237, 32'sd751061, 32'sd838941, -32'sd418506, -32'sd913943, -32'sd2032298, -32'sd233482, -32'sd752043, 32'sd1510608, -32'sd2380768, -32'sd2423264, -32'sd2404548, -32'sd1160725, 32'sd1367435, 32'sd1501403, 32'sd555967, -32'sd127535, 32'sd1467209, 32'sd975412, 32'sd2676826, 32'sd2735553, -32'sd1073900, -32'sd2798824, 32'sd229332, 32'sd93452, -32'sd425510, -32'sd1469682, -32'sd1268574, -32'sd818786, -32'sd1870209, -32'sd830598, -32'sd1252408, -32'sd241273, 32'sd59590, -32'sd603415, 32'sd513911, 32'sd112292, -32'sd191636, -32'sd1347813, -32'sd538567, 32'sd1779746, -32'sd546008, 32'sd973290, -32'sd2436631, -32'sd298709, 32'sd1391717, 32'sd1341300, 32'sd1596373, 32'sd122107, -32'sd925347, -32'sd1450577, 32'sd895130, 32'sd1851164, -32'sd303407, 32'sd2441312, 32'sd1133238, 32'sd1438420, -32'sd983588, -32'sd59906, 32'sd733973, -32'sd1053224, 32'sd539331, 32'sd1648990, -32'sd349393, 32'sd407922, -32'sd586875, 32'sd1059452, 32'sd1963520, 32'sd3432763, 32'sd987277, 32'sd1479363, 32'sd692368, 32'sd666695, -32'sd836634, 32'sd42037, 32'sd529689, -32'sd525604, -32'sd688848, 32'sd76684, 32'sd1714001, 32'sd1572311, 32'sd637830, 32'sd1609306, 32'sd1527511, -32'sd232196, -32'sd772650, 32'sd829368, 32'sd0, 32'sd82465, -32'sd251670, 32'sd1274751, 32'sd2047335, 32'sd86798, -32'sd86585, 32'sd1593706, 32'sd2618642, 32'sd2654790, 32'sd732759, 32'sd575532, -32'sd134366, -32'sd1491712, -32'sd952745, -32'sd1364648, -32'sd552052, -32'sd823449, -32'sd396960, -32'sd380117, 32'sd441078, 32'sd2095076, -32'sd282497, 32'sd2936967, 32'sd891088, -32'sd799913, 32'sd803629, -32'sd616574, -32'sd1204263, -32'sd1171493, -32'sd1166508, 32'sd734480, 32'sd452542, 32'sd986491, 32'sd1326578, 32'sd1377961, 32'sd651525, 32'sd1060225, 32'sd1276246, -32'sd2627, -32'sd2353260, -32'sd2744159, -32'sd2273159, 32'sd781257, -32'sd1772751, 32'sd56348, 32'sd803766, -32'sd1284381, -32'sd362685, 32'sd2239436, 32'sd11447, 32'sd991899, -32'sd609705, -32'sd3036005, -32'sd1222973, -32'sd1177735, -32'sd656287, -32'sd884181, -32'sd840326, -32'sd117490, 32'sd831600, 32'sd1728019, 32'sd1256035, 32'sd300276, 32'sd2336896, -32'sd67644, 32'sd1106926, -32'sd1708032, -32'sd3204094, -32'sd3197143, -32'sd567504, 32'sd723426, -32'sd626439, 32'sd555345, 32'sd588137, 32'sd1421959, -32'sd16977, -32'sd136621, 32'sd2220617, 32'sd1777120, -32'sd867445, -32'sd2327507, 32'sd156144, -32'sd1049229, 32'sd0, 32'sd795759, 32'sd655830, 32'sd407349, 32'sd295832, 32'sd371140, -32'sd517505, 32'sd1124923, 32'sd1397570, -32'sd231772, -32'sd518019, -32'sd2568737, -32'sd2410703, -32'sd404926, 32'sd960186, 32'sd1060510, -32'sd810530, -32'sd1828710, -32'sd1410695, 32'sd796792, -32'sd1604184, -32'sd1087910, -32'sd456715, 32'sd719501, -32'sd606545, -32'sd361126, -32'sd54080, -32'sd935835, -32'sd177407, 32'sd119075, -32'sd363854, -32'sd1662349, -32'sd1998372, 32'sd451882, 32'sd1884027, 32'sd2175709, 32'sd859602, -32'sd1064528, 32'sd1845062, 32'sd1306554, -32'sd588846, -32'sd1333943, 32'sd180738, 32'sd1636393, -32'sd248375, -32'sd572576, -32'sd2065296, -32'sd1449020, -32'sd584887, -32'sd221317, 32'sd419124, -32'sd1092314, -32'sd124629, -32'sd1924821, 32'sd17179, 32'sd152301, -32'sd902883, 32'sd490633, -32'sd1119510, -32'sd358901, -32'sd1915283, -32'sd1235114, 32'sd1866285, 32'sd1281810, -32'sd1919929, 32'sd280807, 32'sd951137, 32'sd313103, 32'sd2039112, 32'sd122898, 32'sd148464, 32'sd194600, 32'sd879805, 32'sd110775, -32'sd1283573, -32'sd658051, 32'sd1582187, -32'sd1360164, 32'sd373087, -32'sd2186237, 32'sd173769, -32'sd1675945, -32'sd750070, -32'sd838502, 32'sd0, 32'sd450617, 32'sd160467, -32'sd909850, 32'sd669680, 32'sd1241131, -32'sd1654138, -32'sd416323, 32'sd571711, -32'sd1266105, 32'sd435464, 32'sd1700501, 32'sd1549615, 32'sd2566756, 32'sd74204, 32'sd338501, -32'sd2211296, -32'sd1963647, -32'sd654492, 32'sd2738771, -32'sd229619, 32'sd309775, 32'sd859382, -32'sd352485, 32'sd1109812, 32'sd1222225, 32'sd1239709, 32'sd0, 32'sd0, 32'sd0, 32'sd1009245, 32'sd1806730, -32'sd1575780, -32'sd274451, 32'sd525084, -32'sd935761, -32'sd734905, 32'sd175760, -32'sd889314, -32'sd811654, 32'sd884421, -32'sd184915, -32'sd25784, -32'sd864739, 32'sd1220830, -32'sd231348, 32'sd40280, -32'sd1576709, -32'sd1537469, -32'sd1294391, -32'sd729871, 32'sd68010, -32'sd1022982, 32'sd35647, -32'sd362900, 32'sd0, 32'sd0, 32'sd0, -32'sd259511, -32'sd1228646, 32'sd514325, 32'sd416950, 32'sd930907, -32'sd612208, -32'sd2554879, 32'sd2136871, 32'sd1085390, 32'sd850385, -32'sd45447, -32'sd1082126, 32'sd471793, -32'sd352796, -32'sd48072, 32'sd220414, -32'sd908899, -32'sd626820, 32'sd206391, 32'sd496719, 32'sd1568759, -32'sd344905, -32'sd640, -32'sd1114540, -32'sd644566, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1000089, -32'sd101189, -32'sd119320, 32'sd801311, -32'sd1191268, -32'sd1350243, 32'sd891493, 32'sd1112494, -32'sd1037329, -32'sd2748470, -32'sd1384846, -32'sd2258237, -32'sd1073406, -32'sd283500, -32'sd1659470, -32'sd1365386, 32'sd1836644, 32'sd385407, 32'sd1613309, -32'sd490652, -32'sd1090380, -32'sd314321, 32'sd469421, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd105957, -32'sd1493253, -32'sd596897, 32'sd193456, -32'sd396243, 32'sd258490, -32'sd1400, -32'sd1815122, -32'sd1662846, -32'sd1607522, 32'sd2953059, 32'sd2673336, 32'sd934883, -32'sd873874, 32'sd614223, -32'sd1692889, -32'sd417709, -32'sd1569321, 32'sd555598, -32'sd1243911, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2764399, 32'sd1223424, 32'sd1176180, 32'sd1291610, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd944454, 32'sd1010906, -32'sd851820, 32'sd197849, 32'sd1245876, -32'sd170773, 32'sd428020, 32'sd936247, 32'sd1494100, 32'sd940910, 32'sd1546862, 32'sd2047449, -32'sd694076, 32'sd48291, 32'sd1451991, 32'sd809659, 32'sd1603454, 32'sd430939, 32'sd1028013, 32'sd493309, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd739251, 32'sd1154966, 32'sd1414989, -32'sd852650, -32'sd1045241, -32'sd1732845, 32'sd1018533, 32'sd2313069, -32'sd4789, 32'sd406224, 32'sd1044545, 32'sd2920994, 32'sd4134679, 32'sd2768712, 32'sd2679040, 32'sd786495, -32'sd1412384, -32'sd1328814, 32'sd279801, -32'sd5308, -32'sd784243, -32'sd1378295, 32'sd648801, 32'sd2076504, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2144972, 32'sd235976, -32'sd582142, 32'sd811747, 32'sd2611517, 32'sd1932437, 32'sd571464, 32'sd843400, 32'sd530183, 32'sd27774, 32'sd330501, 32'sd2058570, -32'sd951561, 32'sd43574, 32'sd958264, 32'sd1642919, 32'sd29708, -32'sd1035365, 32'sd640253, -32'sd2133981, 32'sd37237, -32'sd689619, -32'sd129824, 32'sd420313, 32'sd831195, 32'sd0, 32'sd0, 32'sd751581, -32'sd701638, 32'sd17309, 32'sd247436, 32'sd1125507, 32'sd1517688, -32'sd685698, 32'sd1291901, 32'sd1107082, 32'sd425147, 32'sd2976110, 32'sd2223162, 32'sd3518730, 32'sd1172109, -32'sd2069458, 32'sd872503, -32'sd781652, 32'sd2175030, 32'sd134657, -32'sd1459861, 32'sd32583, 32'sd317748, 32'sd2142346, -32'sd579926, 32'sd1083660, -32'sd240783, 32'sd210998, 32'sd0, 32'sd1058113, 32'sd970156, 32'sd770793, 32'sd883012, 32'sd936968, 32'sd214812, 32'sd1316977, 32'sd2566434, 32'sd2764315, 32'sd1558662, 32'sd899312, 32'sd35767, 32'sd121995, 32'sd403036, -32'sd2007089, -32'sd1780349, -32'sd625309, -32'sd436838, 32'sd901471, -32'sd504155, 32'sd33133, -32'sd1957337, -32'sd1259695, -32'sd278572, -32'sd241714, 32'sd442979, 32'sd901977, 32'sd0, 32'sd1266066, 32'sd108213, -32'sd1362266, 32'sd644107, 32'sd148252, 32'sd1798996, -32'sd486057, 32'sd165099, 32'sd1866021, 32'sd41311, -32'sd870385, -32'sd592000, -32'sd1645537, -32'sd1439204, -32'sd783193, -32'sd3151018, -32'sd2008840, 32'sd423861, -32'sd312240, 32'sd1419783, -32'sd1614970, -32'sd1525431, 32'sd172853, -32'sd19062, -32'sd237933, 32'sd402139, 32'sd492138, 32'sd907972, 32'sd644111, 32'sd690006, -32'sd1574588, -32'sd2719306, -32'sd2005478, 32'sd1144456, -32'sd1201495, -32'sd1683, -32'sd1251884, -32'sd310579, 32'sd276430, 32'sd1504342, 32'sd99141, 32'sd1701507, -32'sd2554296, -32'sd2432151, -32'sd2497101, 32'sd137078, -32'sd1232609, -32'sd907942, 32'sd790326, -32'sd1844429, 32'sd1425768, 32'sd1825673, -32'sd394173, 32'sd1037364, 32'sd218284, -32'sd404365, -32'sd735570, -32'sd512639, -32'sd266472, -32'sd1529234, -32'sd2621108, -32'sd1301082, -32'sd245951, 32'sd531074, 32'sd163488, -32'sd1217194, 32'sd1411848, 32'sd1194654, 32'sd2046374, -32'sd370814, 32'sd259514, -32'sd3445027, -32'sd2660686, 32'sd412733, -32'sd1898205, 32'sd478939, -32'sd616382, -32'sd138122, 32'sd746014, 32'sd873958, 32'sd1294812, 32'sd782858, -32'sd494882, 32'sd299746, 32'sd2051962, 32'sd322024, 32'sd666094, 32'sd84508, -32'sd1536123, -32'sd1316118, 32'sd1201448, -32'sd1344995, -32'sd2863712, -32'sd490798, 32'sd1481502, 32'sd2524652, -32'sd26736, -32'sd382192, -32'sd3926648, -32'sd3207552, -32'sd1061814, -32'sd682977, 32'sd320730, 32'sd2488717, 32'sd1624803, -32'sd277927, -32'sd983215, -32'sd1342609, 32'sd574911, 32'sd613587, -32'sd290581, 32'sd1498784, 32'sd2107834, 32'sd1922685, 32'sd921471, 32'sd903815, -32'sd77759, -32'sd136655, -32'sd626003, 32'sd628357, -32'sd1674402, 32'sd1455983, 32'sd2647178, 32'sd2498022, 32'sd719783, -32'sd2858813, -32'sd4699678, -32'sd2217926, -32'sd535969, 32'sd408693, 32'sd698493, -32'sd222192, 32'sd906778, 32'sd853312, -32'sd1374085, 32'sd824934, 32'sd1657064, -32'sd172461, -32'sd1451284, -32'sd485425, 32'sd626327, -32'sd852135, 32'sd1307069, 32'sd523462, -32'sd446184, 32'sd547708, -32'sd435035, 32'sd898223, 32'sd1984060, 32'sd730041, 32'sd2124574, 32'sd171379, -32'sd1075602, -32'sd2218901, -32'sd3387341, -32'sd1765454, 32'sd613369, 32'sd802161, 32'sd1546110, 32'sd1881538, 32'sd125695, 32'sd848686, 32'sd135311, -32'sd2145979, 32'sd71592, -32'sd1204298, 32'sd750699, 32'sd849877, 32'sd423312, 32'sd393919, -32'sd1609801, 32'sd1494760, 32'sd358849, -32'sd1920180, 32'sd702012, 32'sd1393922, 32'sd1849330, 32'sd1953935, 32'sd2797671, 32'sd1981881, -32'sd3462302, -32'sd3393444, 32'sd165712, 32'sd1351013, -32'sd1026227, 32'sd903660, 32'sd225613, 32'sd644844, -32'sd110109, 32'sd627790, -32'sd2147599, 32'sd2115, -32'sd37614, 32'sd841099, -32'sd1104844, 32'sd1224552, -32'sd174130, 32'sd1726615, -32'sd36221, 32'sd915931, 32'sd191401, 32'sd373510, -32'sd782833, 32'sd1469538, 32'sd575806, 32'sd833758, 32'sd1450276, -32'sd825452, -32'sd3613600, -32'sd1778729, 32'sd404681, 32'sd1320405, 32'sd3233270, 32'sd483942, 32'sd1854061, -32'sd1132971, 32'sd1605295, 32'sd483336, -32'sd1634705, -32'sd628412, -32'sd817228, -32'sd875622, 32'sd554116, 32'sd849537, -32'sd427052, 32'sd444917, 32'sd243181, 32'sd956408, -32'sd1225503, 32'sd263846, 32'sd1997772, 32'sd2253682, -32'sd32901, -32'sd1894934, -32'sd1560763, -32'sd2367373, -32'sd1155547, -32'sd636594, 32'sd1655356, 32'sd1404586, 32'sd2286108, 32'sd1224310, -32'sd33842, 32'sd1286393, -32'sd1045217, 32'sd1208472, -32'sd51264, -32'sd944143, -32'sd79254, -32'sd148214, 32'sd1035459, 32'sd840442, 32'sd531783, -32'sd284217, 32'sd894837, -32'sd901392, -32'sd536978, 32'sd1366254, 32'sd2091474, 32'sd1860463, -32'sd656249, 32'sd80224, -32'sd2073396, -32'sd2766470, -32'sd1698022, 32'sd471412, 32'sd2974036, 32'sd1335655, 32'sd566486, -32'sd2296453, 32'sd1646771, 32'sd3020770, 32'sd136646, 32'sd1023307, -32'sd321789, -32'sd1112847, 32'sd1578843, -32'sd1792569, 32'sd290512, 32'sd804078, -32'sd1006915, 32'sd1395746, -32'sd210100, 32'sd1388191, 32'sd630430, 32'sd2593521, 32'sd1189081, 32'sd683757, -32'sd715616, -32'sd2234498, -32'sd2311284, -32'sd1411286, 32'sd163071, 32'sd1830434, 32'sd3437575, 32'sd3962216, 32'sd1336877, 32'sd731303, 32'sd1359296, 32'sd2360307, 32'sd667100, -32'sd1323520, -32'sd518001, 32'sd371599, 32'sd1656924, 32'sd503040, 32'sd1006757, 32'sd0, -32'sd243962, -32'sd360145, 32'sd555726, 32'sd3109422, -32'sd1465379, 32'sd49393, -32'sd748359, -32'sd944054, -32'sd2125755, -32'sd3357364, -32'sd2402557, -32'sd1563423, 32'sd2199040, 32'sd1341443, 32'sd3588917, 32'sd2342687, 32'sd2316152, 32'sd2562992, 32'sd2122453, 32'sd1170791, 32'sd2003134, 32'sd267877, -32'sd110254, 32'sd308316, 32'sd1821508, 32'sd1273265, 32'sd11854, -32'sd540653, 32'sd643808, 32'sd372457, -32'sd918633, 32'sd2291140, 32'sd1272949, -32'sd138021, 32'sd142471, -32'sd1252359, -32'sd1120999, -32'sd3904461, -32'sd2129806, 32'sd510056, 32'sd1391904, 32'sd1883817, 32'sd1949780, 32'sd3931157, 32'sd2365421, 32'sd3305768, 32'sd1025027, -32'sd101852, 32'sd1228764, -32'sd1303552, -32'sd509361, 32'sd1092951, 32'sd2095816, 32'sd896396, 32'sd474741, 32'sd1279967, 32'sd40931, 32'sd361700, -32'sd1901112, -32'sd257445, -32'sd45231, -32'sd86967, 32'sd671105, 32'sd1186441, -32'sd599528, -32'sd3502846, -32'sd1518224, -32'sd290773, -32'sd1435189, 32'sd1579462, 32'sd2182395, 32'sd1511552, 32'sd1956703, 32'sd56135, -32'sd633158, -32'sd554767, -32'sd4546, -32'sd132033, -32'sd983888, 32'sd694058, 32'sd946068, 32'sd227066, 32'sd82477, 32'sd0, 32'sd185112, 32'sd603872, -32'sd512285, -32'sd1079576, -32'sd971938, -32'sd267415, 32'sd1218233, -32'sd382867, -32'sd1526192, -32'sd772493, -32'sd949742, -32'sd376021, -32'sd2163987, 32'sd980479, 32'sd784327, 32'sd1684735, 32'sd1613948, 32'sd1873297, -32'sd1675865, -32'sd2256777, -32'sd586047, -32'sd778131, 32'sd1087563, 32'sd1549674, 32'sd615706, 32'sd458669, -32'sd240533, 32'sd661041, 32'sd170437, 32'sd633077, -32'sd804466, -32'sd1072018, -32'sd271029, -32'sd115506, -32'sd349944, -32'sd1073766, 32'sd826874, 32'sd969827, -32'sd669349, -32'sd12017, 32'sd506763, -32'sd2700511, -32'sd1347700, -32'sd1491620, 32'sd144961, -32'sd93757, 32'sd858375, -32'sd1232670, -32'sd687579, 32'sd331730, -32'sd1233387, -32'sd50097, 32'sd1015121, 32'sd330820, 32'sd311711, 32'sd1264847, 32'sd348762, -32'sd619077, 32'sd1434858, -32'sd625025, 32'sd965872, -32'sd119844, -32'sd1468061, -32'sd642951, 32'sd880477, -32'sd468282, -32'sd2362638, -32'sd1603009, -32'sd1505755, -32'sd3087886, -32'sd651457, -32'sd476431, -32'sd1579499, 32'sd731872, 32'sd1530814, 32'sd1368359, 32'sd920120, -32'sd347238, -32'sd168679, -32'sd2108757, -32'sd1427438, 32'sd31038, 32'sd1415627, 32'sd0, 32'sd1153880, -32'sd569744, 32'sd613366, -32'sd839845, -32'sd634168, 32'sd304973, 32'sd850158, -32'sd1151508, 32'sd715551, -32'sd254118, -32'sd2678121, -32'sd1699694, -32'sd711484, -32'sd1483159, -32'sd1750455, -32'sd1159353, 32'sd47090, -32'sd1054708, 32'sd1293651, 32'sd1967371, 32'sd85392, 32'sd826322, 32'sd1917656, -32'sd681629, 32'sd936748, 32'sd788017, 32'sd0, 32'sd0, 32'sd0, 32'sd83196, 32'sd1229370, -32'sd101431, -32'sd1704551, 32'sd111393, 32'sd505234, 32'sd1115720, 32'sd1210428, 32'sd997675, 32'sd2035806, -32'sd151687, -32'sd189155, -32'sd303280, -32'sd433495, -32'sd1791493, -32'sd1512654, 32'sd435293, 32'sd585431, -32'sd394863, 32'sd731254, -32'sd886829, 32'sd425278, -32'sd876514, 32'sd1402641, 32'sd924778, 32'sd0, 32'sd0, 32'sd0, 32'sd471503, 32'sd142468, 32'sd112796, 32'sd23483, 32'sd812549, 32'sd797123, 32'sd27468, 32'sd2659718, 32'sd896173, 32'sd561864, 32'sd649168, -32'sd1744407, 32'sd3607, -32'sd1905477, -32'sd327650, -32'sd217468, 32'sd595886, -32'sd147484, -32'sd1784830, -32'sd1173556, -32'sd268517, -32'sd37737, 32'sd1168850, 32'sd919043, 32'sd551038, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1083371, 32'sd324011, -32'sd2440846, -32'sd1443216, -32'sd1787192, 32'sd14186, 32'sd919360, -32'sd1406145, -32'sd515175, -32'sd141719, 32'sd761241, -32'sd1048148, -32'sd1806520, -32'sd1447321, 32'sd24226, -32'sd436426, 32'sd791321, 32'sd819465, -32'sd307783, -32'sd346414, 32'sd854880, 32'sd73748, 32'sd940519, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1691282, 32'sd1531616, -32'sd523381, 32'sd1258338, 32'sd476280, 32'sd1324760, 32'sd354941, -32'sd543271, -32'sd461435, -32'sd836834, -32'sd1398490, -32'sd1617579, -32'sd1324726, 32'sd734931, -32'sd388901, -32'sd887216, 32'sd547938, 32'sd423791, 32'sd289336, 32'sd1310855, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1925572, -32'sd144367, 32'sd2203471, 32'sd1992589, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd540181, 32'sd971041, 32'sd878318, 32'sd1037999, 32'sd179707, 32'sd1694351, 32'sd235631, 32'sd1628670, 32'sd897473, 32'sd2266629, 32'sd579558, -32'sd588904, 32'sd275692, -32'sd265641, 32'sd1204201, 32'sd1318700, 32'sd608439, 32'sd1615849, 32'sd200157, 32'sd901433, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd554043, 32'sd711297, -32'sd742324, -32'sd629358, 32'sd439043, 32'sd2046688, 32'sd2146575, 32'sd2170276, 32'sd2102781, 32'sd2070196, 32'sd1616632, 32'sd537498, 32'sd1817197, -32'sd692271, -32'sd467739, 32'sd704942, 32'sd1521753, -32'sd1237001, -32'sd981292, 32'sd1288167, 32'sd1565968, -32'sd1294005, 32'sd2617796, 32'sd680486, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd669428, 32'sd958261, 32'sd685438, 32'sd883386, 32'sd823715, 32'sd456638, 32'sd843418, 32'sd1868367, -32'sd1101144, -32'sd897340, 32'sd1786725, 32'sd296091, -32'sd457142, -32'sd1040088, 32'sd565349, 32'sd813813, -32'sd1003404, 32'sd226304, -32'sd599158, -32'sd480560, -32'sd278503, 32'sd130986, 32'sd746182, -32'sd368770, -32'sd1760529, 32'sd0, 32'sd0, 32'sd523306, 32'sd917545, -32'sd331272, -32'sd358280, -32'sd642729, -32'sd1063147, 32'sd861734, -32'sd253208, 32'sd1176776, 32'sd2018180, 32'sd1639307, -32'sd298332, 32'sd1937102, 32'sd665097, -32'sd278292, 32'sd582417, 32'sd43010, 32'sd633240, -32'sd167627, -32'sd84115, -32'sd404316, -32'sd1421111, -32'sd658939, -32'sd448873, 32'sd184232, -32'sd131755, 32'sd1023374, 32'sd0, 32'sd301530, 32'sd1074182, -32'sd75537, 32'sd1554813, 32'sd418036, -32'sd1001142, 32'sd397732, 32'sd1699052, -32'sd708531, -32'sd247724, -32'sd1257453, 32'sd1424968, 32'sd2154390, -32'sd1092663, -32'sd466803, -32'sd519335, -32'sd2724019, -32'sd1403331, 32'sd596442, -32'sd30178, -32'sd294143, -32'sd2296708, 32'sd169719, 32'sd820541, -32'sd300780, 32'sd215404, 32'sd55877, 32'sd0, 32'sd1021986, -32'sd1352876, 32'sd1365277, -32'sd114826, 32'sd708593, -32'sd1237650, 32'sd415429, -32'sd851766, -32'sd248801, 32'sd1214563, 32'sd1362370, 32'sd888935, 32'sd1635554, 32'sd243719, -32'sd495253, -32'sd1105402, -32'sd1265546, -32'sd1127425, -32'sd1729129, -32'sd4747, -32'sd2107294, 32'sd192219, -32'sd1983849, -32'sd677790, -32'sd1064765, 32'sd374441, -32'sd1653069, 32'sd1138918, 32'sd1497934, -32'sd1720616, 32'sd1398410, -32'sd159449, -32'sd1418498, -32'sd2301472, -32'sd719235, -32'sd117787, 32'sd1549565, 32'sd153936, -32'sd194324, 32'sd1225227, 32'sd1208616, 32'sd625256, 32'sd2180287, -32'sd1608785, -32'sd579395, 32'sd584637, -32'sd766304, -32'sd2464483, -32'sd852891, 32'sd425389, -32'sd503763, -32'sd3134886, -32'sd446967, 32'sd1237378, 32'sd196012, 32'sd1401472, 32'sd1795845, -32'sd1763247, -32'sd5770, 32'sd1891595, -32'sd1578424, -32'sd1361313, -32'sd784083, 32'sd967183, 32'sd422504, 32'sd1657616, -32'sd593767, -32'sd438735, 32'sd1161495, 32'sd1022125, 32'sd801536, 32'sd951225, 32'sd69873, -32'sd1884232, -32'sd315345, -32'sd877480, -32'sd527498, -32'sd2279091, -32'sd269844, -32'sd2604726, 32'sd55612, 32'sd643723, -32'sd840730, 32'sd182075, -32'sd257120, -32'sd798760, -32'sd1192728, -32'sd858444, 32'sd1600602, 32'sd1194977, 32'sd863283, 32'sd807703, -32'sd244522, -32'sd2021673, -32'sd213762, -32'sd1566876, -32'sd268802, 32'sd952195, -32'sd1199021, -32'sd431602, 32'sd776805, 32'sd42733, -32'sd1346161, -32'sd1802219, -32'sd589923, -32'sd1439524, -32'sd1563827, -32'sd240400, -32'sd936778, -32'sd611336, 32'sd899749, 32'sd1181645, 32'sd1139377, 32'sd1371929, -32'sd1226321, -32'sd1734274, 32'sd1262188, 32'sd1249361, -32'sd449507, -32'sd1950842, -32'sd3159928, -32'sd2446120, -32'sd2228580, -32'sd1446696, -32'sd1506009, -32'sd1013359, -32'sd2198361, -32'sd1390168, -32'sd124765, 32'sd193036, 32'sd1102041, -32'sd996864, -32'sd724172, -32'sd1689951, -32'sd931543, -32'sd124703, -32'sd1187179, -32'sd1430481, 32'sd753464, 32'sd111754, -32'sd953495, -32'sd908719, -32'sd958122, -32'sd307295, -32'sd1082276, 32'sd838372, -32'sd1994213, -32'sd1156702, -32'sd3284070, -32'sd1007132, -32'sd2976491, -32'sd4295263, -32'sd818079, 32'sd780585, 32'sd1513460, -32'sd1072453, -32'sd1781276, -32'sd1061928, -32'sd2252334, -32'sd587980, -32'sd144538, -32'sd521502, -32'sd782759, -32'sd668570, 32'sd1213304, -32'sd640432, 32'sd17758, 32'sd605892, -32'sd1133020, -32'sd1754070, -32'sd957567, -32'sd837800, -32'sd2244781, -32'sd3522971, -32'sd3133700, -32'sd2290964, -32'sd2541620, -32'sd1976854, -32'sd1808787, -32'sd686971, -32'sd283799, 32'sd4002880, 32'sd1566347, -32'sd116418, -32'sd2193, 32'sd1206838, -32'sd1729198, -32'sd163579, 32'sd888339, -32'sd747332, 32'sd303071, -32'sd916136, 32'sd251865, -32'sd308967, 32'sd201286, 32'sd1064717, 32'sd92376, 32'sd248800, 32'sd62596, -32'sd163218, -32'sd1215422, -32'sd1880614, -32'sd2089240, -32'sd1180432, 32'sd191595, 32'sd1222506, -32'sd755394, 32'sd499577, 32'sd939080, 32'sd2498604, 32'sd1112699, -32'sd473999, -32'sd693864, 32'sd928228, 32'sd1685680, 32'sd699706, 32'sd1222056, 32'sd410961, -32'sd1287499, 32'sd1304750, 32'sd1226267, -32'sd811278, 32'sd431222, 32'sd508715, -32'sd380461, -32'sd1000842, 32'sd1315820, -32'sd721176, 32'sd476933, -32'sd1366039, -32'sd538968, -32'sd865296, 32'sd1371321, 32'sd1575557, 32'sd2775274, 32'sd2117463, 32'sd582323, 32'sd1327732, -32'sd2595924, 32'sd553119, -32'sd1878512, 32'sd260952, 32'sd2304595, 32'sd1312099, 32'sd1470750, 32'sd1081744, -32'sd1530252, -32'sd1156281, 32'sd435173, -32'sd1844113, 32'sd2034472, 32'sd1224142, 32'sd335576, -32'sd450884, 32'sd150444, 32'sd175623, -32'sd517797, -32'sd604000, 32'sd1309526, 32'sd718052, 32'sd1644085, 32'sd2674341, 32'sd3288532, 32'sd338726, 32'sd1402339, 32'sd186145, -32'sd3066369, -32'sd1755729, -32'sd2365249, 32'sd707073, 32'sd1059864, -32'sd761411, 32'sd971516, -32'sd1374537, 32'sd355270, 32'sd1046613, 32'sd763731, -32'sd1444676, 32'sd333149, 32'sd1173237, 32'sd108642, 32'sd518410, 32'sd895662, -32'sd380806, 32'sd1324946, -32'sd32824, 32'sd1694316, 32'sd1234160, 32'sd1985088, 32'sd2818715, 32'sd698214, 32'sd157202, -32'sd938631, -32'sd679013, -32'sd1970203, -32'sd2821714, -32'sd3654709, -32'sd2366040, -32'sd1554534, -32'sd173967, 32'sd189785, -32'sd659729, 32'sd526860, 32'sd145712, 32'sd449590, 32'sd679194, -32'sd510032, 32'sd0, 32'sd592350, 32'sd222992, -32'sd1386137, -32'sd2443667, -32'sd1369566, 32'sd586190, -32'sd568807, -32'sd389408, 32'sd1353897, 32'sd2246892, 32'sd791356, -32'sd344538, -32'sd1828459, -32'sd51509, -32'sd2283127, -32'sd448227, -32'sd1169733, -32'sd1279467, 32'sd139192, -32'sd1167870, 32'sd1478793, 32'sd2210404, 32'sd2167835, -32'sd112886, 32'sd1415628, 32'sd537629, 32'sd810611, -32'sd430970, 32'sd1434223, 32'sd451754, 32'sd382524, -32'sd766706, -32'sd1113873, -32'sd484039, 32'sd53243, 32'sd28879, 32'sd599370, 32'sd664948, 32'sd447809, -32'sd92069, 32'sd1814755, 32'sd903803, 32'sd780749, 32'sd521926, -32'sd275273, -32'sd763129, -32'sd745897, -32'sd711839, -32'sd281565, -32'sd43401, 32'sd61738, -32'sd791586, 32'sd1061343, 32'sd973281, 32'sd384974, 32'sd78340, -32'sd129138, -32'sd423658, -32'sd1907846, -32'sd194951, 32'sd33737, -32'sd1927534, -32'sd748927, -32'sd2318926, 32'sd670224, 32'sd1557925, 32'sd78927, -32'sd445714, -32'sd301205, 32'sd631782, -32'sd572466, 32'sd1674406, 32'sd2232164, 32'sd787151, -32'sd2186222, 32'sd77055, 32'sd77989, -32'sd151231, 32'sd565879, -32'sd743843, -32'sd1295009, 32'sd496400, 32'sd62738, 32'sd0, 32'sd20617, 32'sd94147, -32'sd563190, -32'sd1715068, 32'sd196609, -32'sd2291400, -32'sd2268380, 32'sd286035, 32'sd859092, 32'sd2148004, 32'sd39906, 32'sd2257391, 32'sd2040265, 32'sd2360701, 32'sd1360153, 32'sd913668, -32'sd351911, 32'sd645046, -32'sd2086565, -32'sd1452540, -32'sd417218, 32'sd1704070, 32'sd1151332, 32'sd417769, -32'sd871166, -32'sd403504, 32'sd654000, -32'sd11913, 32'sd826396, 32'sd241499, 32'sd401025, -32'sd83619, -32'sd2338133, -32'sd3424266, -32'sd508384, -32'sd682517, 32'sd1602140, 32'sd2151724, 32'sd2532565, 32'sd1032536, 32'sd2408468, 32'sd1784025, 32'sd1335221, 32'sd1173822, 32'sd1331446, 32'sd702364, -32'sd1176816, -32'sd1520870, -32'sd105631, 32'sd724210, 32'sd36150, -32'sd385602, -32'sd188981, -32'sd553105, 32'sd465512, 32'sd1486850, 32'sd371589, -32'sd379930, 32'sd802642, -32'sd1158736, -32'sd821187, -32'sd185115, -32'sd1138888, 32'sd123992, 32'sd1789140, 32'sd1224210, 32'sd774961, 32'sd1195090, 32'sd1072073, -32'sd140900, 32'sd1790336, -32'sd901850, -32'sd1598820, -32'sd393337, 32'sd1093687, 32'sd1455407, 32'sd1198819, 32'sd2124388, 32'sd234046, 32'sd260962, -32'sd470267, 32'sd10667, 32'sd386885, 32'sd0, 32'sd852814, -32'sd464567, 32'sd422630, -32'sd1147428, 32'sd756449, -32'sd38861, -32'sd1741382, -32'sd504014, 32'sd941156, 32'sd1397227, 32'sd741790, 32'sd438450, 32'sd1231733, 32'sd508989, 32'sd167484, 32'sd1598623, -32'sd319899, -32'sd1965903, 32'sd1073165, 32'sd1297300, 32'sd346204, 32'sd167121, -32'sd828712, -32'sd2168050, -32'sd1289123, -32'sd109448, 32'sd0, 32'sd0, 32'sd0, -32'sd806968, 32'sd116451, 32'sd463877, -32'sd734659, -32'sd2520857, -32'sd1393753, -32'sd2343662, -32'sd990536, -32'sd1106701, -32'sd806585, 32'sd250406, -32'sd306143, 32'sd664794, -32'sd2496840, -32'sd1336993, -32'sd837625, 32'sd106609, 32'sd28983, 32'sd613843, -32'sd1219133, -32'sd551454, -32'sd1846501, -32'sd2006187, 32'sd1543109, 32'sd737810, 32'sd0, 32'sd0, 32'sd0, 32'sd921958, -32'sd199810, 32'sd237691, -32'sd867147, 32'sd485502, 32'sd14185, 32'sd480370, -32'sd1742525, -32'sd930662, 32'sd1649242, 32'sd1816077, -32'sd830272, 32'sd105818, -32'sd3187466, -32'sd346536, 32'sd293191, 32'sd1460554, -32'sd1367468, 32'sd1168093, -32'sd281709, -32'sd2550869, -32'sd2601849, 32'sd597938, 32'sd810286, 32'sd531300, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd856976, 32'sd431603, 32'sd760624, -32'sd492119, 32'sd35121, 32'sd1574242, 32'sd553485, 32'sd1066460, -32'sd88816, -32'sd1549404, -32'sd1025063, 32'sd383050, -32'sd7635, -32'sd279030, 32'sd420213, 32'sd1111962, 32'sd94399, -32'sd1647175, -32'sd341825, 32'sd518567, 32'sd919073, -32'sd1027178, 32'sd869227, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd894759, 32'sd559816, 32'sd1197633, 32'sd992101, 32'sd807025, 32'sd1053419, 32'sd51562, 32'sd544666, 32'sd1368823, 32'sd486867, 32'sd435128, 32'sd1322828, 32'sd282108, 32'sd980736, -32'sd357761, 32'sd3018, 32'sd133965, -32'sd1223669, 32'sd872827, -32'sd139537, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd45110, -32'sd848929, 32'sd640926, 32'sd1336041, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1207334, 32'sd863856, 32'sd188936, -32'sd405870, 32'sd950227, 32'sd1108444, 32'sd824305, 32'sd90430, -32'sd748321, 32'sd336478, 32'sd208097, 32'sd1057499, 32'sd269192, 32'sd657579, 32'sd726851, 32'sd528838, 32'sd1327566, 32'sd1546166, -32'sd735802, -32'sd25375, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd194764, -32'sd231264, 32'sd1245492, 32'sd820437, 32'sd136845, -32'sd925564, 32'sd631069, 32'sd714706, -32'sd592897, 32'sd651982, 32'sd73103, 32'sd877963, 32'sd2067752, 32'sd1647461, 32'sd1122612, 32'sd1891962, 32'sd1845032, 32'sd2249621, 32'sd595025, 32'sd2772578, 32'sd1553779, 32'sd264562, 32'sd719993, 32'sd1104840, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd914447, -32'sd304429, -32'sd121975, -32'sd638088, 32'sd1060904, -32'sd2364520, -32'sd470460, -32'sd85761, -32'sd1916724, -32'sd197467, 32'sd1391404, 32'sd2905854, -32'sd177223, -32'sd176872, 32'sd14143, 32'sd2237835, 32'sd156023, 32'sd405999, -32'sd197412, -32'sd279957, -32'sd151254, 32'sd738859, 32'sd995627, -32'sd241990, 32'sd863007, 32'sd0, 32'sd0, 32'sd711114, -32'sd63346, 32'sd221236, -32'sd635480, -32'sd46102, -32'sd180146, -32'sd1453843, -32'sd1209821, -32'sd841743, 32'sd183362, -32'sd782389, -32'sd1183896, 32'sd249118, -32'sd352815, 32'sd762605, 32'sd1305397, 32'sd933236, -32'sd465327, -32'sd222909, -32'sd2198665, -32'sd399624, 32'sd353188, 32'sd224670, 32'sd38271, -32'sd1597584, 32'sd391496, 32'sd621072, 32'sd0, 32'sd307363, -32'sd1063761, 32'sd330392, -32'sd1807623, -32'sd679891, -32'sd1840873, -32'sd641609, -32'sd333256, -32'sd3004892, -32'sd1274258, -32'sd1139843, -32'sd3173999, -32'sd441640, 32'sd2948070, 32'sd2703560, 32'sd282303, 32'sd358194, -32'sd989382, -32'sd1714513, -32'sd700294, -32'sd49756, -32'sd1419945, 32'sd104112, 32'sd924687, 32'sd1349405, 32'sd800550, -32'sd908049, 32'sd0, 32'sd560028, -32'sd595053, -32'sd1675887, -32'sd3154517, -32'sd491895, -32'sd1087790, -32'sd807591, -32'sd2174263, -32'sd2111051, 32'sd127808, 32'sd236505, 32'sd104621, 32'sd2161563, 32'sd2787654, 32'sd2539260, -32'sd597743, -32'sd975587, -32'sd1735275, -32'sd3196383, -32'sd2395846, -32'sd1384666, 32'sd19133, -32'sd2204593, 32'sd764782, -32'sd1375722, 32'sd422617, -32'sd2105995, 32'sd681419, 32'sd115023, -32'sd1281464, -32'sd440556, -32'sd560044, -32'sd826879, -32'sd414237, -32'sd1208587, -32'sd521027, 32'sd1135581, -32'sd244298, 32'sd1944710, 32'sd1766182, 32'sd207053, 32'sd690132, 32'sd2301313, -32'sd444062, 32'sd192225, 32'sd767439, -32'sd705487, -32'sd3450360, -32'sd2619317, -32'sd300765, 32'sd206127, 32'sd2019412, 32'sd1010688, 32'sd211646, -32'sd1463484, -32'sd77247, 32'sd1285487, 32'sd1773778, -32'sd1003495, -32'sd1440790, -32'sd518068, -32'sd124665, 32'sd81949, 32'sd2443429, -32'sd834887, 32'sd711812, -32'sd456285, 32'sd295996, 32'sd120159, 32'sd3365613, 32'sd4167547, -32'sd812886, -32'sd352889, 32'sd928697, -32'sd1691304, -32'sd3354439, 32'sd73513, -32'sd337649, 32'sd933507, 32'sd1087895, 32'sd1268207, 32'sd670727, -32'sd727049, -32'sd267617, -32'sd20038, 32'sd2874648, -32'sd405575, -32'sd461019, 32'sd1455778, 32'sd1126039, 32'sd1231193, 32'sd755470, 32'sd61133, -32'sd1045328, -32'sd2019314, -32'sd1499066, 32'sd861920, 32'sd3104755, 32'sd883026, -32'sd1229690, -32'sd1072192, -32'sd1308683, -32'sd1135954, -32'sd67956, -32'sd154410, 32'sd1467248, 32'sd1448895, -32'sd516765, 32'sd1201273, -32'sd730892, 32'sd360887, 32'sd104261, 32'sd67716, 32'sd1318391, 32'sd397518, 32'sd762830, -32'sd216270, -32'sd199966, -32'sd483534, -32'sd1721082, -32'sd3068325, -32'sd3708560, -32'sd3064874, -32'sd492066, 32'sd1420624, 32'sd2124199, 32'sd1941471, -32'sd1106897, -32'sd1374925, -32'sd2247213, -32'sd1555609, 32'sd553750, 32'sd887305, 32'sd2429679, 32'sd1472208, -32'sd274908, 32'sd14073, 32'sd1096840, 32'sd1345790, -32'sd601091, 32'sd667384, 32'sd1629712, 32'sd1287145, 32'sd444235, -32'sd998685, 32'sd66055, -32'sd1429026, -32'sd2768931, -32'sd2861480, -32'sd3626897, -32'sd1929724, 32'sd2065243, 32'sd3506595, -32'sd49177, -32'sd2250678, -32'sd2580627, -32'sd1217219, -32'sd2817798, -32'sd1283887, 32'sd1075715, 32'sd4251, 32'sd2165706, 32'sd567197, 32'sd1081998, 32'sd1025290, 32'sd9423, -32'sd961796, -32'sd235000, -32'sd188589, -32'sd590529, -32'sd868250, -32'sd641000, -32'sd2002881, -32'sd1768662, -32'sd1609672, -32'sd3510445, -32'sd2367168, -32'sd730169, 32'sd193647, 32'sd3365134, 32'sd1634292, -32'sd1182317, -32'sd3458158, -32'sd3761880, -32'sd774574, -32'sd639393, -32'sd64625, -32'sd350693, 32'sd1224449, 32'sd1166186, -32'sd50978, 32'sd1772343, 32'sd611816, 32'sd286934, 32'sd1380665, 32'sd242816, 32'sd595506, -32'sd1096010, 32'sd1838928, -32'sd14211, -32'sd1604498, -32'sd1722054, -32'sd176857, 32'sd1403189, 32'sd765865, 32'sd1990526, 32'sd3108998, 32'sd2029373, 32'sd543912, -32'sd2536914, -32'sd3641711, -32'sd3474979, -32'sd812381, 32'sd747161, 32'sd1976967, -32'sd923772, 32'sd256963, -32'sd2062, 32'sd814568, 32'sd1596063, 32'sd492637, 32'sd1228653, 32'sd1379861, 32'sd41911, 32'sd419760, -32'sd470231, -32'sd476342, 32'sd279773, 32'sd1308490, -32'sd416075, -32'sd990443, 32'sd849997, 32'sd2107001, 32'sd1440092, 32'sd1604426, -32'sd181742, -32'sd3080380, -32'sd2787149, -32'sd2071648, -32'sd1382833, -32'sd890662, -32'sd170087, 32'sd1043483, -32'sd136273, -32'sd1223188, 32'sd22610, 32'sd348135, -32'sd2072, 32'sd720678, -32'sd658687, 32'sd1345278, 32'sd153171, -32'sd732632, -32'sd1184913, -32'sd58431, -32'sd2059812, 32'sd372165, -32'sd380879, 32'sd840261, 32'sd2194988, 32'sd1875970, 32'sd1925510, 32'sd1771831, -32'sd238576, -32'sd3314349, -32'sd3428983, -32'sd872461, 32'sd780441, 32'sd490436, -32'sd21865, 32'sd416183, 32'sd761951, 32'sd994742, 32'sd1459664, -32'sd1262893, -32'sd56643, 32'sd193558, -32'sd1172660, 32'sd861572, 32'sd316361, 32'sd697358, 32'sd95278, -32'sd101605, -32'sd566277, -32'sd97631, -32'sd1066984, 32'sd1242226, 32'sd343960, 32'sd2301236, 32'sd1904131, 32'sd2066813, -32'sd1504031, -32'sd1658088, -32'sd2735777, -32'sd37430, 32'sd867164, 32'sd42296, -32'sd1708972, -32'sd1332306, -32'sd651936, 32'sd445461, 32'sd1319060, 32'sd624401, 32'sd1291919, 32'sd771875, 32'sd604175, 32'sd1022504, 32'sd0, -32'sd253400, -32'sd922063, -32'sd1540105, 32'sd628015, 32'sd1113792, 32'sd1690751, 32'sd129489, -32'sd998125, 32'sd989315, -32'sd842595, -32'sd579406, -32'sd47863, -32'sd1296977, -32'sd590719, 32'sd222047, 32'sd1371987, -32'sd672253, -32'sd650817, 32'sd604616, -32'sd515812, -32'sd768205, 32'sd424338, 32'sd376989, -32'sd380728, 32'sd1209526, -32'sd1458144, 32'sd1114462, -32'sd327813, -32'sd1188492, -32'sd661046, -32'sd3310874, -32'sd402249, -32'sd733670, 32'sd226096, 32'sd289951, 32'sd1093415, 32'sd2573181, -32'sd563019, -32'sd530662, -32'sd1520567, -32'sd1074153, -32'sd2133308, 32'sd669494, 32'sd48562, -32'sd1342348, 32'sd1051048, -32'sd1272366, 32'sd609172, 32'sd419912, 32'sd1389482, -32'sd1011326, -32'sd395711, -32'sd717444, -32'sd2187897, -32'sd718284, 32'sd275214, 32'sd755089, -32'sd1575086, -32'sd2601442, 32'sd510523, 32'sd791406, -32'sd245339, 32'sd780314, 32'sd1550579, 32'sd953139, 32'sd633405, -32'sd213397, -32'sd891084, 32'sd568079, -32'sd1768122, 32'sd900716, 32'sd1126866, -32'sd732499, 32'sd125334, 32'sd232257, -32'sd1130751, 32'sd996485, 32'sd2667665, 32'sd1041523, -32'sd1549060, 32'sd811254, -32'sd376205, -32'sd957973, 32'sd0, -32'sd1265042, 32'sd173785, -32'sd1500612, -32'sd1551656, -32'sd1016034, 32'sd1408937, 32'sd3349620, 32'sd205891, 32'sd2569752, 32'sd1553677, 32'sd1345785, 32'sd2261297, -32'sd421055, -32'sd832805, 32'sd1379918, 32'sd436093, -32'sd117003, 32'sd1090174, -32'sd89920, 32'sd1830747, 32'sd504078, 32'sd289552, 32'sd1269870, -32'sd1728189, 32'sd703955, 32'sd763327, -32'sd462827, 32'sd312960, 32'sd908468, -32'sd252478, -32'sd1462084, 32'sd471916, -32'sd3992, -32'sd179797, -32'sd844979, 32'sd1592370, 32'sd714471, 32'sd197352, 32'sd1397018, 32'sd1309059, 32'sd670595, 32'sd843093, -32'sd205650, 32'sd504654, 32'sd290605, 32'sd632595, -32'sd138895, -32'sd1231687, 32'sd914339, 32'sd2008796, 32'sd648206, 32'sd354077, 32'sd66515, 32'sd948355, 32'sd169707, 32'sd1661274, 32'sd594147, -32'sd882225, 32'sd52103, -32'sd466806, 32'sd1071176, 32'sd719659, 32'sd292340, 32'sd2014294, 32'sd1172569, 32'sd1483903, 32'sd639015, 32'sd2746962, 32'sd72139, -32'sd2828607, -32'sd1461771, -32'sd2739761, -32'sd541423, -32'sd1345703, 32'sd283135, -32'sd1196710, -32'sd1041857, 32'sd1676752, -32'sd1372475, -32'sd611116, -32'sd242146, 32'sd2292430, 32'sd1047393, 32'sd0, -32'sd169945, 32'sd1377031, -32'sd2429380, -32'sd270981, -32'sd1145769, -32'sd563239, 32'sd2235627, 32'sd1024822, 32'sd1302867, 32'sd1778926, 32'sd1220646, 32'sd2167453, -32'sd2142988, -32'sd3089434, -32'sd1016958, -32'sd2121833, -32'sd273500, -32'sd1286861, -32'sd1369649, 32'sd53012, 32'sd396916, -32'sd684987, -32'sd1222921, -32'sd1517811, -32'sd1428688, 32'sd1164339, 32'sd0, 32'sd0, 32'sd0, 32'sd828051, -32'sd777727, 32'sd161501, -32'sd745575, -32'sd204092, 32'sd2378238, 32'sd1707639, 32'sd69587, -32'sd452009, -32'sd180681, 32'sd2351735, 32'sd1196560, 32'sd1155805, 32'sd187078, 32'sd1265600, -32'sd401851, 32'sd1092249, -32'sd1173483, -32'sd475010, 32'sd595828, 32'sd1165151, 32'sd54976, -32'sd570002, 32'sd821425, 32'sd330482, 32'sd0, 32'sd0, 32'sd0, -32'sd1014211, -32'sd63180, -32'sd2220760, -32'sd864029, -32'sd476518, -32'sd2497878, -32'sd1697876, 32'sd806482, -32'sd934152, 32'sd365493, 32'sd161864, -32'sd211501, 32'sd619278, -32'sd568426, -32'sd937153, -32'sd1336106, -32'sd137178, 32'sd313655, -32'sd746310, -32'sd945771, -32'sd725490, 32'sd317203, -32'sd2055218, 32'sd203363, 32'sd201790, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd386276, 32'sd46299, -32'sd484063, -32'sd996310, -32'sd2122504, -32'sd1830200, 32'sd269243, 32'sd563676, 32'sd1332866, -32'sd1353172, 32'sd679268, 32'sd2983668, 32'sd1424429, 32'sd163031, 32'sd480847, -32'sd648693, -32'sd1030903, -32'sd673752, -32'sd926779, -32'sd1980011, 32'sd145261, -32'sd267319, 32'sd359018, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd540803, 32'sd1052771, -32'sd449302, 32'sd1372658, -32'sd704129, 32'sd553149, -32'sd322143, -32'sd1610956, 32'sd396360, -32'sd11528, -32'sd1151731, -32'sd953203, -32'sd484143, 32'sd846992, 32'sd292653, -32'sd1226372, -32'sd1209744, 32'sd914502, -32'sd344426, 32'sd799861, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1136915, 32'sd403940, 32'sd1488199, 32'sd1772924, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd86920, 32'sd1051060, 32'sd1490435, 32'sd1153955, 32'sd2430811, 32'sd1546646, 32'sd1178907, 32'sd131948, -32'sd890769, -32'sd1209871, 32'sd907096, 32'sd1579318, 32'sd824584, 32'sd1349303, 32'sd1185912, -32'sd49959, 32'sd1200986, 32'sd325450, 32'sd793344, 32'sd413903, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd629780, -32'sd1119997, -32'sd296298, -32'sd586108, 32'sd82135, -32'sd225141, -32'sd875215, 32'sd602199, -32'sd673333, 32'sd232258, 32'sd284100, -32'sd742024, 32'sd838972, -32'sd116022, 32'sd290906, 32'sd484508, -32'sd454499, 32'sd1961845, 32'sd189125, 32'sd1375071, -32'sd724604, 32'sd248653, -32'sd418320, 32'sd1324921, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd590541, 32'sd635397, 32'sd611995, -32'sd444189, -32'sd471721, -32'sd857149, -32'sd1843323, -32'sd491436, -32'sd142433, -32'sd1860221, -32'sd2542848, 32'sd1634315, 32'sd433213, 32'sd1433492, 32'sd1700588, 32'sd1447859, 32'sd2046486, -32'sd1199692, 32'sd1136542, 32'sd1204726, 32'sd1285678, -32'sd125347, -32'sd305893, 32'sd1923379, -32'sd105877, 32'sd0, 32'sd0, 32'sd440250, 32'sd471373, -32'sd1534431, 32'sd363792, 32'sd349003, 32'sd930902, 32'sd1081503, 32'sd1434519, 32'sd1952159, 32'sd545116, -32'sd388882, -32'sd269702, 32'sd1687466, -32'sd1921397, 32'sd1192019, 32'sd1860273, 32'sd1019263, 32'sd1198520, 32'sd936404, 32'sd1841134, 32'sd1066347, 32'sd983319, 32'sd598263, -32'sd389895, -32'sd410947, -32'sd533755, 32'sd851059, 32'sd0, 32'sd251522, -32'sd973990, 32'sd1449916, 32'sd1887960, 32'sd1158356, 32'sd1292552, -32'sd1202665, 32'sd940284, 32'sd403541, 32'sd1903493, 32'sd1006602, -32'sd369812, 32'sd2855882, 32'sd2025966, 32'sd1987179, 32'sd429032, 32'sd114620, 32'sd1242884, 32'sd3263809, 32'sd1254710, 32'sd1353268, 32'sd2446999, -32'sd823662, -32'sd1462162, -32'sd39367, -32'sd62324, -32'sd637263, 32'sd0, 32'sd353171, 32'sd160156, 32'sd989850, -32'sd742059, -32'sd374769, 32'sd1037052, 32'sd2157174, 32'sd972750, 32'sd2118509, 32'sd1247008, 32'sd1827819, -32'sd526525, 32'sd95587, -32'sd2125761, 32'sd1543680, 32'sd1266560, 32'sd1780138, 32'sd1214395, 32'sd2287582, 32'sd2056696, 32'sd235946, 32'sd632855, -32'sd1016208, -32'sd380055, -32'sd57793, -32'sd1091486, 32'sd534247, 32'sd1165215, -32'sd980182, 32'sd396338, -32'sd1030346, 32'sd1234075, 32'sd1517591, 32'sd2611402, -32'sd228006, 32'sd46596, -32'sd466292, 32'sd2742149, 32'sd881828, -32'sd523117, -32'sd575088, -32'sd1905362, -32'sd996509, 32'sd899406, 32'sd1044169, 32'sd462335, 32'sd904873, 32'sd1090991, 32'sd627989, 32'sd1126407, -32'sd242369, -32'sd414927, 32'sd611186, -32'sd918890, 32'sd87935, 32'sd1077747, 32'sd1069704, 32'sd1589593, -32'sd992276, -32'sd432416, 32'sd3016456, 32'sd1413235, -32'sd817694, 32'sd1182918, -32'sd852085, 32'sd2201, -32'sd804321, -32'sd2244515, -32'sd2659631, -32'sd1027886, 32'sd1318733, -32'sd1305240, -32'sd123082, 32'sd1445472, 32'sd950067, 32'sd1015686, 32'sd1168162, 32'sd521586, 32'sd397452, -32'sd1021920, -32'sd229859, -32'sd1202991, 32'sd472199, -32'sd311890, 32'sd843958, -32'sd1147505, -32'sd2639184, -32'sd230185, 32'sd6499, 32'sd60236, -32'sd19555, 32'sd1991574, 32'sd35813, 32'sd260446, -32'sd1202215, -32'sd2928882, -32'sd571499, -32'sd2283680, -32'sd1328410, -32'sd3453912, -32'sd1369194, -32'sd457604, -32'sd94678, -32'sd778230, 32'sd1075741, 32'sd312913, -32'sd1590449, -32'sd487964, 32'sd1205315, -32'sd470358, 32'sd579771, 32'sd526545, 32'sd246083, 32'sd1460978, -32'sd864993, 32'sd2267283, -32'sd319831, -32'sd530388, 32'sd405788, 32'sd1864114, 32'sd1332346, 32'sd793055, -32'sd1337735, -32'sd1683878, -32'sd3553525, -32'sd3285290, -32'sd3227990, -32'sd2918713, -32'sd2218969, -32'sd2051024, -32'sd2530699, -32'sd3199121, 32'sd1188082, 32'sd429740, -32'sd82146, 32'sd576547, 32'sd988908, -32'sd1488534, 32'sd374615, -32'sd1097413, 32'sd1001590, 32'sd1727629, -32'sd654518, -32'sd1130509, 32'sd232453, -32'sd179111, 32'sd917694, -32'sd1515661, -32'sd850478, -32'sd1377499, -32'sd3433989, -32'sd1636272, -32'sd3472618, -32'sd3692032, -32'sd4238201, -32'sd2689573, -32'sd2532185, -32'sd1541887, -32'sd2654385, -32'sd2513627, -32'sd52180, 32'sd639965, 32'sd1735407, 32'sd1175675, -32'sd858511, -32'sd1549959, 32'sd769659, 32'sd378565, 32'sd881822, -32'sd462640, 32'sd1280517, -32'sd1359326, -32'sd57786, 32'sd655810, 32'sd1264151, 32'sd250977, -32'sd1533452, -32'sd812839, -32'sd2171738, -32'sd1382207, -32'sd3782856, -32'sd2915652, -32'sd2789237, -32'sd1611511, -32'sd1127035, -32'sd3600221, -32'sd241191, -32'sd554045, -32'sd17567, 32'sd1115124, -32'sd1153585, -32'sd207481, -32'sd745452, -32'sd630301, 32'sd1539991, 32'sd469652, -32'sd159258, 32'sd893847, 32'sd1733569, 32'sd1836455, -32'sd256230, -32'sd109902, -32'sd757479, -32'sd541248, -32'sd1547172, 32'sd230623, -32'sd319273, -32'sd2573968, -32'sd2479774, -32'sd2157528, -32'sd2062759, -32'sd1255188, -32'sd503040, -32'sd1710780, 32'sd984358, 32'sd144632, 32'sd1655222, 32'sd1658806, 32'sd537425, -32'sd697161, 32'sd582947, 32'sd209663, 32'sd1672227, 32'sd1626304, 32'sd548209, -32'sd577660, 32'sd1001101, 32'sd793262, 32'sd1313379, -32'sd507696, 32'sd1296522, 32'sd1029111, -32'sd50859, 32'sd111100, -32'sd473825, 32'sd489582, 32'sd1408635, 32'sd1297321, 32'sd623833, -32'sd1908236, -32'sd423890, -32'sd363302, 32'sd829489, 32'sd2103291, 32'sd1620708, 32'sd628516, 32'sd6041, 32'sd844371, -32'sd126714, 32'sd1880935, 32'sd573785, 32'sd1896632, 32'sd991733, 32'sd829767, 32'sd785928, -32'sd175937, -32'sd805461, -32'sd438422, -32'sd1123145, 32'sd714595, 32'sd1690927, 32'sd351003, 32'sd166551, 32'sd237007, 32'sd554892, 32'sd702674, 32'sd384403, -32'sd1461241, -32'sd1046236, 32'sd1003801, 32'sd2418989, 32'sd785589, 32'sd2282538, 32'sd1561699, -32'sd1094302, 32'sd526446, 32'sd1109032, -32'sd5748, -32'sd570796, 32'sd413202, -32'sd1019888, -32'sd628473, 32'sd287877, 32'sd635171, 32'sd725553, 32'sd656510, -32'sd570381, -32'sd88744, -32'sd615232, -32'sd1160791, 32'sd126200, -32'sd1352527, -32'sd1132451, -32'sd993813, -32'sd2365809, -32'sd3421224, -32'sd2570751, 32'sd695408, -32'sd288954, 32'sd2299267, 32'sd2578996, -32'sd537887, -32'sd773667, -32'sd1695444, 32'sd700124, 32'sd1319915, -32'sd263243, 32'sd0, -32'sd1516655, -32'sd2021593, -32'sd266328, -32'sd1060807, -32'sd341291, 32'sd1858741, 32'sd2655295, 32'sd703582, -32'sd1219019, -32'sd210591, -32'sd2190433, -32'sd668185, -32'sd2539506, -32'sd2756677, -32'sd4362782, -32'sd3462462, 32'sd419421, 32'sd1708297, -32'sd57878, 32'sd2059683, 32'sd220159, -32'sd401092, -32'sd1085238, -32'sd481435, -32'sd250969, 32'sd359715, 32'sd1238632, 32'sd305626, 32'sd713276, -32'sd1378798, 32'sd1848095, 32'sd774567, -32'sd1254582, 32'sd2529906, 32'sd3565264, -32'sd159794, 32'sd295100, 32'sd2247020, -32'sd1409047, -32'sd1859661, -32'sd3194266, -32'sd2293270, -32'sd2385873, -32'sd305847, 32'sd1932414, 32'sd1363824, 32'sd440434, 32'sd794936, -32'sd946305, -32'sd1427619, -32'sd2289855, -32'sd2139688, 32'sd285422, 32'sd1273830, 32'sd99151, 32'sd540898, 32'sd926228, -32'sd1256260, 32'sd2108327, -32'sd171768, -32'sd1412435, 32'sd3094321, 32'sd1513696, 32'sd332817, 32'sd2082534, 32'sd734277, -32'sd1295507, 32'sd246588, -32'sd2353806, 32'sd606235, 32'sd684819, 32'sd1087393, 32'sd1116481, 32'sd1546774, -32'sd201164, -32'sd1115712, 32'sd201919, 32'sd1428132, -32'sd1338454, -32'sd138984, 32'sd19023, -32'sd285209, -32'sd1526870, 32'sd0, -32'sd278434, 32'sd48845, 32'sd1099727, -32'sd466376, 32'sd1299687, 32'sd2412609, 32'sd1270074, 32'sd1340859, 32'sd1958905, -32'sd222829, 32'sd954640, -32'sd246721, -32'sd697779, -32'sd990603, -32'sd780516, 32'sd2290800, 32'sd2861883, 32'sd2737995, 32'sd1026344, -32'sd244675, 32'sd1569157, 32'sd738042, 32'sd457071, -32'sd659926, -32'sd1578664, 32'sd172509, 32'sd150585, 32'sd1092123, 32'sd1035336, 32'sd680055, 32'sd2762923, -32'sd838390, -32'sd942154, 32'sd1430210, 32'sd2089755, 32'sd755947, -32'sd310389, -32'sd1537448, -32'sd1104973, -32'sd232017, -32'sd43920, 32'sd1959358, 32'sd980569, 32'sd2504390, 32'sd1718955, 32'sd331272, 32'sd472159, -32'sd167236, -32'sd298229, 32'sd954151, -32'sd360811, 32'sd1481966, 32'sd1260310, -32'sd403563, -32'sd470080, 32'sd2117122, 32'sd1468825, 32'sd9508, 32'sd1584412, -32'sd54434, -32'sd304462, -32'sd395566, -32'sd122535, 32'sd843108, 32'sd652045, 32'sd363752, 32'sd1788881, -32'sd438856, 32'sd1929468, 32'sd2889431, 32'sd1741711, 32'sd2681306, 32'sd2079556, 32'sd2261872, 32'sd964937, -32'sd97333, -32'sd715479, 32'sd1408580, 32'sd1857557, 32'sd2396006, 32'sd302798, -32'sd251242, 32'sd697647, 32'sd0, 32'sd1310228, 32'sd1801042, -32'sd589744, -32'sd1520144, -32'sd215013, -32'sd495550, -32'sd1290387, -32'sd1170284, 32'sd1931911, 32'sd2580205, 32'sd2666122, 32'sd2012841, 32'sd2512131, 32'sd2692996, 32'sd993131, 32'sd2378351, 32'sd2061712, 32'sd1634151, 32'sd211831, 32'sd102993, 32'sd682775, 32'sd600117, -32'sd339818, 32'sd1347048, 32'sd1164668, -32'sd497560, 32'sd0, 32'sd0, 32'sd0, -32'sd206520, 32'sd648173, -32'sd782936, -32'sd175636, -32'sd767466, -32'sd22088, 32'sd1069422, -32'sd934580, -32'sd838222, -32'sd1229, 32'sd2233850, 32'sd2659012, 32'sd239898, 32'sd478403, -32'sd493185, 32'sd375787, -32'sd823055, -32'sd647679, 32'sd589577, 32'sd169440, -32'sd18339, -32'sd5381, 32'sd986292, 32'sd1125877, 32'sd586847, 32'sd0, 32'sd0, 32'sd0, 32'sd176256, 32'sd791122, -32'sd941913, -32'sd656524, -32'sd895606, -32'sd123020, 32'sd816928, -32'sd522223, 32'sd936451, -32'sd1798319, -32'sd2553191, 32'sd816090, -32'sd28523, -32'sd1579290, -32'sd2677836, -32'sd466531, 32'sd2028182, 32'sd729227, -32'sd953076, -32'sd2206844, -32'sd168413, 32'sd1166555, 32'sd525611, 32'sd365578, 32'sd1020985, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1274607, 32'sd958573, -32'sd784642, 32'sd392087, -32'sd315342, 32'sd119318, 32'sd1262852, -32'sd134131, -32'sd1995870, -32'sd2041292, 32'sd361867, -32'sd941544, -32'sd2492223, -32'sd715724, -32'sd3586002, -32'sd1340789, -32'sd666818, -32'sd1978009, -32'sd195223, -32'sd609011, -32'sd34758, 32'sd1071638, 32'sd81039, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1354013, -32'sd592842, 32'sd1113381, 32'sd496114, -32'sd391321, 32'sd652064, 32'sd613292, 32'sd886058, 32'sd1300008, -32'sd79067, 32'sd836524, 32'sd1490214, -32'sd233148, 32'sd356537, 32'sd292654, -32'sd1129941, 32'sd1054251, -32'sd469585, -32'sd532016, 32'sd496083, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd582102, 32'sd154993, -32'sd185552, -32'sd675480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd525045, -32'sd1795200, -32'sd433893, 32'sd88505, -32'sd2059893, 32'sd319536, -32'sd1067953, -32'sd1233874, -32'sd301359, -32'sd678831, 32'sd246554, -32'sd826775, -32'sd1129517, -32'sd1387113, -32'sd319155, -32'sd248828, 32'sd1409320, 32'sd288465, -32'sd887780, 32'sd9007, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd107014, 32'sd514926, -32'sd536689, -32'sd396606, -32'sd689823, -32'sd567939, -32'sd780012, -32'sd289624, -32'sd2087504, -32'sd802422, -32'sd283394, -32'sd514376, -32'sd1741060, -32'sd151422, 32'sd616983, -32'sd607767, -32'sd61860, 32'sd450742, 32'sd190906, 32'sd596330, -32'sd484117, 32'sd1878280, 32'sd1312599, 32'sd209, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd543570, 32'sd145791, -32'sd1151877, -32'sd247128, 32'sd374852, -32'sd1269441, -32'sd1363960, 32'sd732330, -32'sd1215359, -32'sd2362136, -32'sd1572410, -32'sd3203095, -32'sd3036676, -32'sd1810631, 32'sd2677087, 32'sd2390962, 32'sd1255399, 32'sd73995, -32'sd2117911, -32'sd1396520, -32'sd539846, -32'sd483575, -32'sd496677, -32'sd407228, 32'sd353315, 32'sd0, 32'sd0, 32'sd876021, -32'sd495571, 32'sd884125, 32'sd455449, 32'sd654586, -32'sd1250078, -32'sd1420999, -32'sd847999, -32'sd45275, -32'sd474350, -32'sd733707, -32'sd1420713, -32'sd3254133, -32'sd1821332, -32'sd1135177, -32'sd801300, 32'sd878563, 32'sd271860, 32'sd390708, -32'sd1736487, -32'sd1345874, -32'sd2925928, -32'sd3499459, -32'sd2361385, 32'sd904735, -32'sd1767829, 32'sd783504, 32'sd0, -32'sd13167, -32'sd512353, 32'sd19659, 32'sd605554, 32'sd538383, 32'sd695236, -32'sd540339, 32'sd1365243, -32'sd119746, 32'sd1900456, 32'sd1974330, 32'sd646770, 32'sd1521459, -32'sd79041, 32'sd243570, -32'sd1161044, -32'sd1794085, 32'sd241304, 32'sd652769, -32'sd1592801, -32'sd184639, -32'sd1887244, -32'sd519135, -32'sd416593, 32'sd836118, -32'sd24505, 32'sd87412, 32'sd0, -32'sd734315, 32'sd194563, 32'sd114884, -32'sd1624669, -32'sd566720, 32'sd689634, 32'sd236406, -32'sd361506, 32'sd567410, 32'sd254399, 32'sd1263100, 32'sd1310681, 32'sd1311487, -32'sd378401, -32'sd921427, -32'sd1141633, 32'sd532271, 32'sd375932, 32'sd2058309, 32'sd798434, 32'sd2865860, -32'sd1692158, -32'sd297207, -32'sd1252065, -32'sd98160, -32'sd619166, -32'sd361280, -32'sd569941, -32'sd609485, -32'sd547783, 32'sd1070573, 32'sd259535, -32'sd1058980, 32'sd1894104, 32'sd1394491, 32'sd736619, 32'sd1309999, 32'sd354551, -32'sd449247, -32'sd63735, -32'sd1693496, -32'sd1644191, -32'sd843845, 32'sd1748183, 32'sd258967, 32'sd2250597, 32'sd1363329, 32'sd1354804, 32'sd1743340, 32'sd438155, 32'sd677936, -32'sd271472, 32'sd257303, 32'sd912577, -32'sd409312, 32'sd561645, 32'sd1232820, -32'sd344367, -32'sd725078, 32'sd1453023, -32'sd638694, 32'sd148535, -32'sd725626, 32'sd2571438, 32'sd2056404, -32'sd1142920, -32'sd1640403, -32'sd62253, -32'sd738061, 32'sd448541, 32'sd1071777, 32'sd1087687, -32'sd1204703, 32'sd1089752, -32'sd499155, 32'sd580510, 32'sd816682, 32'sd595889, 32'sd118426, -32'sd206503, -32'sd754330, -32'sd16189, 32'sd942260, -32'sd450360, 32'sd239374, -32'sd463030, -32'sd495750, 32'sd2052325, 32'sd895875, 32'sd920464, -32'sd442813, -32'sd266750, -32'sd838677, -32'sd881766, -32'sd695908, -32'sd219892, -32'sd106060, -32'sd140195, -32'sd978796, 32'sd1438765, 32'sd627751, -32'sd312302, -32'sd903314, 32'sd584194, 32'sd304583, -32'sd142355, -32'sd758232, 32'sd542912, 32'sd427415, 32'sd59160, 32'sd84336, 32'sd595835, -32'sd603321, 32'sd98921, -32'sd1537292, -32'sd430464, 32'sd835418, 32'sd1332046, 32'sd842738, 32'sd1716176, 32'sd2118633, -32'sd454798, -32'sd1060544, -32'sd469910, 32'sd104726, 32'sd467314, -32'sd1577127, 32'sd1184063, 32'sd865005, -32'sd1032451, 32'sd139056, -32'sd1581343, 32'sd187538, 32'sd1803324, 32'sd1525082, 32'sd1231647, 32'sd332618, 32'sd783859, -32'sd164188, 32'sd305930, 32'sd393814, 32'sd1093803, 32'sd494458, 32'sd865764, -32'sd549424, -32'sd278366, 32'sd944479, 32'sd586506, 32'sd1683384, 32'sd2987155, -32'sd155142, -32'sd868819, -32'sd1448816, -32'sd5418, -32'sd1120116, -32'sd1017418, -32'sd1478076, -32'sd1034924, -32'sd1351035, -32'sd942191, 32'sd371846, 32'sd2065733, -32'sd758469, 32'sd1606690, -32'sd404474, -32'sd393592, -32'sd2482197, 32'sd743082, 32'sd777341, 32'sd43061, 32'sd1714402, 32'sd6831, -32'sd329514, -32'sd144805, 32'sd276456, -32'sd127140, 32'sd401251, 32'sd1875154, -32'sd704872, 32'sd223839, -32'sd531701, -32'sd2706544, -32'sd905452, -32'sd937494, 32'sd346947, 32'sd590125, -32'sd634236, 32'sd170821, -32'sd166297, 32'sd1994671, 32'sd1089973, 32'sd2493045, -32'sd1646695, -32'sd2029060, -32'sd909889, -32'sd384487, 32'sd1305761, 32'sd705353, 32'sd1663208, 32'sd526979, 32'sd664741, 32'sd1139864, 32'sd860862, 32'sd452463, -32'sd234235, 32'sd781948, -32'sd1206446, -32'sd2105626, -32'sd2383733, -32'sd2137360, -32'sd422137, -32'sd188999, 32'sd992847, -32'sd1522248, 32'sd614904, 32'sd790755, 32'sd2822647, 32'sd3516305, 32'sd899302, -32'sd413331, -32'sd914556, 32'sd279495, -32'sd185955, -32'sd428476, 32'sd105566, -32'sd90758, -32'sd385644, -32'sd853632, 32'sd1244147, 32'sd410770, -32'sd232330, -32'sd928693, 32'sd161780, -32'sd1174862, -32'sd587209, 32'sd824435, -32'sd697124, -32'sd641905, 32'sd711509, -32'sd768806, 32'sd2754063, 32'sd2546314, 32'sd1900906, 32'sd1637338, 32'sd2701503, 32'sd847563, -32'sd135428, 32'sd216328, 32'sd573019, 32'sd1899326, 32'sd579948, -32'sd531934, 32'sd606274, 32'sd989061, 32'sd1751744, -32'sd1434449, 32'sd990795, 32'sd72642, 32'sd845368, -32'sd926206, -32'sd637602, -32'sd2063467, 32'sd654436, -32'sd803216, 32'sd535975, 32'sd1143349, 32'sd2469239, -32'sd1283, 32'sd3264342, 32'sd887621, 32'sd121290, 32'sd1153867, 32'sd717983, -32'sd270634, 32'sd399489, 32'sd1969528, 32'sd1623363, 32'sd1701774, 32'sd882637, 32'sd228311, -32'sd1064618, -32'sd334184, 32'sd63717, 32'sd1229992, 32'sd1660718, 32'sd187394, -32'sd5271, -32'sd286636, -32'sd4409598, -32'sd1912706, 32'sd52322, 32'sd934080, 32'sd98245, 32'sd498839, 32'sd170677, 32'sd2167125, 32'sd1507687, 32'sd956916, 32'sd39258, 32'sd1348230, 32'sd2138137, -32'sd958131, 32'sd715287, -32'sd209985, -32'sd1159622, 32'sd304081, -32'sd999427, 32'sd0, -32'sd222679, -32'sd34061, 32'sd668286, 32'sd1434518, 32'sd708031, -32'sd491315, -32'sd2399389, -32'sd2346970, -32'sd4662772, -32'sd2512485, 32'sd2621100, 32'sd2374427, 32'sd507826, 32'sd782315, 32'sd1580674, 32'sd1112417, -32'sd609960, -32'sd519828, 32'sd1809493, 32'sd622471, 32'sd778281, 32'sd1910404, 32'sd403219, 32'sd208770, 32'sd1102151, 32'sd2358200, 32'sd1962605, -32'sd489835, 32'sd500549, -32'sd1106985, 32'sd576478, -32'sd1381257, -32'sd513057, -32'sd710171, -32'sd2329414, -32'sd3507490, -32'sd2452070, -32'sd603851, 32'sd2187343, 32'sd2698548, 32'sd2251066, 32'sd523794, -32'sd52109, -32'sd820096, -32'sd118209, -32'sd852921, -32'sd745959, 32'sd543600, 32'sd1410400, -32'sd13707, -32'sd1268157, -32'sd253930, -32'sd1037598, 32'sd1284934, 32'sd1678287, -32'sd213192, 32'sd1000511, 32'sd143885, -32'sd367506, -32'sd1998758, -32'sd1470201, -32'sd3665328, -32'sd2727347, -32'sd2672703, 32'sd1342796, 32'sd4297474, 32'sd1624773, 32'sd427238, 32'sd224377, -32'sd715924, -32'sd240503, -32'sd71253, -32'sd2071234, -32'sd1892760, -32'sd927585, -32'sd1784597, 32'sd52088, -32'sd2211410, -32'sd2941736, -32'sd169383, -32'sd1308600, 32'sd702069, 32'sd1622284, 32'sd0, 32'sd425108, 32'sd1007781, -32'sd876894, -32'sd2407818, -32'sd1065959, -32'sd2719996, -32'sd2511439, 32'sd611030, 32'sd760412, 32'sd3602928, 32'sd2515766, 32'sd43440, -32'sd967737, -32'sd14387, -32'sd788041, -32'sd1224070, -32'sd2714280, -32'sd889913, -32'sd1988726, -32'sd2369653, -32'sd884275, -32'sd1416291, -32'sd2365845, 32'sd1253856, 32'sd586538, -32'sd807636, -32'sd68342, 32'sd260528, -32'sd633178, -32'sd1756961, 32'sd735072, -32'sd723641, -32'sd2206630, -32'sd3136297, -32'sd3802041, -32'sd71917, 32'sd477879, 32'sd826127, 32'sd1066876, 32'sd1488130, 32'sd1186975, -32'sd1790514, -32'sd2113603, -32'sd997498, -32'sd2493956, -32'sd3101246, -32'sd1652762, -32'sd1457820, -32'sd1968905, -32'sd1829156, -32'sd1343793, 32'sd1437650, -32'sd1791891, -32'sd1317708, -32'sd652167, -32'sd518441, -32'sd447924, 32'sd292693, -32'sd970820, -32'sd1685950, -32'sd2483200, -32'sd2791298, -32'sd1673741, -32'sd2137243, -32'sd183495, -32'sd280818, 32'sd1094528, 32'sd4055705, 32'sd3772655, 32'sd928066, -32'sd453732, -32'sd1775405, -32'sd2246668, -32'sd2149138, -32'sd1780129, -32'sd1192212, -32'sd253566, -32'sd284186, 32'sd609099, -32'sd93916, 32'sd224734, 32'sd838923, 32'sd386963, 32'sd0, -32'sd105540, 32'sd48558, -32'sd1886674, 32'sd733390, -32'sd1786058, -32'sd1813506, -32'sd692908, -32'sd671540, -32'sd429687, -32'sd1689698, 32'sd291022, 32'sd3463631, 32'sd4752236, 32'sd1320846, 32'sd282914, -32'sd1170712, -32'sd2061736, -32'sd1824651, -32'sd3455740, -32'sd1794186, 32'sd988652, 32'sd629709, 32'sd465825, -32'sd524540, -32'sd1264451, -32'sd409327, 32'sd0, 32'sd0, 32'sd0, 32'sd863744, 32'sd501458, 32'sd1239242, -32'sd477633, -32'sd1017752, -32'sd418316, -32'sd1279530, -32'sd1536610, 32'sd538967, 32'sd493496, 32'sd1010005, 32'sd464743, 32'sd1071732, 32'sd3213518, 32'sd2458237, -32'sd578974, -32'sd1612088, 32'sd741219, -32'sd27019, -32'sd286558, 32'sd1006913, 32'sd813559, -32'sd1956530, -32'sd1067375, -32'sd479787, 32'sd0, 32'sd0, 32'sd0, -32'sd527027, -32'sd661514, -32'sd1772147, -32'sd2114044, -32'sd497028, -32'sd490317, 32'sd277152, 32'sd1237718, 32'sd453919, 32'sd18576, -32'sd281204, -32'sd851715, 32'sd2319024, 32'sd658113, 32'sd1824632, -32'sd1290568, 32'sd335404, -32'sd886267, -32'sd734110, -32'sd2224487, -32'sd1184232, 32'sd228654, 32'sd660072, 32'sd340603, -32'sd565992, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd462693, 32'sd588218, 32'sd754813, -32'sd511260, 32'sd115574, -32'sd1685089, 32'sd869332, 32'sd634530, -32'sd1071543, -32'sd1021534, 32'sd1395231, 32'sd1113640, 32'sd342836, 32'sd505699, 32'sd653473, 32'sd477066, -32'sd386474, 32'sd539905, 32'sd2322, -32'sd572638, 32'sd636331, 32'sd935801, 32'sd399031, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd381379, -32'sd875110, -32'sd269280, 32'sd1141181, -32'sd279461, 32'sd14505, 32'sd434687, 32'sd799048, -32'sd792382, -32'sd378243, 32'sd123262, -32'sd809522, -32'sd179272, 32'sd2041836, 32'sd1355920, -32'sd553205, 32'sd2186, -32'sd675673, -32'sd1784978, 32'sd355263, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd202967, -32'sd981040, 32'sd31609, -32'sd157225, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd294640, -32'sd563333, 32'sd661801, -32'sd707624, -32'sd638646, 32'sd748916, 32'sd26395, -32'sd1233708, -32'sd1777205, -32'sd2022309, -32'sd1595322, 32'sd338943, 32'sd1000424, 32'sd299461, 32'sd1650336, 32'sd453928, -32'sd1114251, -32'sd613833, -32'sd298642, 32'sd1038540, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd870966, 32'sd411453, -32'sd851990, -32'sd913160, 32'sd370625, -32'sd1275301, 32'sd1039655, 32'sd2045930, -32'sd510636, 32'sd2039998, 32'sd245193, 32'sd1209152, 32'sd1738262, 32'sd2408723, -32'sd263282, 32'sd1287555, 32'sd233005, 32'sd948844, 32'sd1190768, 32'sd2004225, 32'sd372187, -32'sd154755, -32'sd768817, -32'sd1077651, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd624249, 32'sd552706, -32'sd65763, 32'sd562940, 32'sd128254, -32'sd1421484, 32'sd1334379, -32'sd860209, 32'sd910608, 32'sd1778437, 32'sd1624687, 32'sd1346133, -32'sd378925, 32'sd781966, -32'sd276023, -32'sd419692, 32'sd1398902, -32'sd154059, 32'sd430217, -32'sd2055562, -32'sd2748114, 32'sd525664, 32'sd800188, 32'sd109156, -32'sd994553, 32'sd0, 32'sd0, 32'sd1252412, -32'sd797210, 32'sd158821, 32'sd357151, -32'sd1881411, -32'sd1553142, -32'sd317423, 32'sd2000988, 32'sd544192, 32'sd1490556, 32'sd995818, 32'sd1437925, 32'sd2248650, 32'sd1182558, 32'sd500503, 32'sd2970842, -32'sd394115, -32'sd207508, 32'sd359599, -32'sd1005575, 32'sd160783, -32'sd908658, -32'sd288666, -32'sd192482, -32'sd2304350, 32'sd638987, -32'sd387177, 32'sd0, -32'sd715496, -32'sd482301, -32'sd1099938, -32'sd1263445, -32'sd1603033, 32'sd291448, 32'sd1194204, 32'sd845463, 32'sd749417, 32'sd1430469, 32'sd812641, 32'sd4832, 32'sd1890428, 32'sd391456, -32'sd144662, 32'sd1349057, -32'sd987160, -32'sd674776, 32'sd1102106, -32'sd408497, -32'sd1342373, 32'sd66600, 32'sd1102840, -32'sd914002, -32'sd1481522, -32'sd77052, -32'sd980755, 32'sd0, -32'sd995140, 32'sd799204, 32'sd1158333, 32'sd1194581, 32'sd797750, -32'sd239201, 32'sd444426, -32'sd822681, 32'sd1477290, 32'sd2227523, -32'sd566616, -32'sd208586, 32'sd445225, -32'sd1670898, 32'sd587978, -32'sd1863362, -32'sd207402, 32'sd343882, -32'sd843000, 32'sd49170, 32'sd1084677, 32'sd342810, -32'sd783224, -32'sd1142949, -32'sd1274993, -32'sd207006, -32'sd986844, -32'sd288257, -32'sd253393, -32'sd454364, 32'sd2370530, 32'sd1905704, -32'sd1017147, 32'sd1177094, 32'sd1974546, 32'sd780811, -32'sd323147, 32'sd2162225, -32'sd746914, -32'sd538693, -32'sd1778141, -32'sd993595, -32'sd2226134, 32'sd41227, 32'sd333162, -32'sd1345875, -32'sd1041801, -32'sd946388, -32'sd1009664, -32'sd658325, -32'sd1342226, -32'sd1400308, 32'sd198953, 32'sd255637, 32'sd425781, -32'sd21094, -32'sd361454, -32'sd1491911, -32'sd1443729, -32'sd829659, 32'sd425901, 32'sd651570, -32'sd138915, -32'sd1215358, -32'sd301001, -32'sd1921602, -32'sd1486617, -32'sd282424, -32'sd576446, -32'sd319809, 32'sd1091872, 32'sd1510333, 32'sd481361, -32'sd2334647, -32'sd852204, -32'sd195689, 32'sd291878, 32'sd1358729, -32'sd101002, -32'sd1116783, -32'sd631940, 32'sd23206, -32'sd244320, -32'sd729581, 32'sd856550, 32'sd696976, -32'sd931385, 32'sd516723, 32'sd605336, -32'sd1899687, 32'sd193566, -32'sd2096065, -32'sd2199678, -32'sd2350280, -32'sd1849805, 32'sd808804, 32'sd1556365, 32'sd2180257, 32'sd1397169, -32'sd218095, 32'sd153891, -32'sd1585698, -32'sd665675, 32'sd2125202, -32'sd553078, 32'sd2344974, 32'sd2862605, -32'sd9477, 32'sd1378873, -32'sd1937733, -32'sd575093, 32'sd108734, -32'sd1220381, 32'sd94073, 32'sd296302, -32'sd1192759, -32'sd1136228, -32'sd989777, -32'sd2198899, -32'sd1352705, 32'sd271733, 32'sd29868, 32'sd798263, 32'sd672407, 32'sd4436683, 32'sd319704, -32'sd1087399, -32'sd204826, -32'sd695504, 32'sd642078, -32'sd1631912, 32'sd1479938, 32'sd2090959, 32'sd2494586, 32'sd2623998, 32'sd1046267, -32'sd486323, -32'sd1234992, -32'sd524099, -32'sd706206, 32'sd2270105, -32'sd1025917, -32'sd1262387, -32'sd1584913, -32'sd2072372, -32'sd1382892, -32'sd990157, 32'sd473876, 32'sd1391194, 32'sd3131514, 32'sd2305914, 32'sd3429463, 32'sd275832, -32'sd2399909, -32'sd2242253, -32'sd3252664, -32'sd2179658, 32'sd72707, 32'sd842805, 32'sd1758583, -32'sd100948, 32'sd353256, 32'sd473895, 32'sd1668412, -32'sd890900, -32'sd244106, -32'sd544081, -32'sd186842, -32'sd612078, -32'sd876327, -32'sd202652, -32'sd1318464, 32'sd57580, -32'sd60116, 32'sd3729378, 32'sd2927230, 32'sd4159543, 32'sd4563784, 32'sd2521171, 32'sd1456078, -32'sd3284568, -32'sd2445044, -32'sd3639905, -32'sd57465, -32'sd786159, -32'sd1402919, -32'sd2150906, -32'sd1834110, -32'sd250287, 32'sd799526, -32'sd440702, -32'sd631446, -32'sd43221, -32'sd909122, -32'sd135811, 32'sd932025, 32'sd533092, -32'sd1388376, -32'sd510424, 32'sd86619, -32'sd1811028, 32'sd305992, 32'sd3430938, 32'sd5078183, 32'sd4682091, 32'sd1269514, 32'sd6328, -32'sd3062829, -32'sd3724639, -32'sd1387369, -32'sd2905985, -32'sd512648, 32'sd298233, -32'sd2500808, -32'sd4550788, -32'sd763874, -32'sd957054, -32'sd17429, 32'sd1045687, -32'sd534086, 32'sd42995, 32'sd1111627, 32'sd641444, -32'sd671306, -32'sd219986, -32'sd1243593, -32'sd552114, -32'sd739112, 32'sd678732, -32'sd250083, -32'sd54710, 32'sd1818847, -32'sd757133, -32'sd2622446, -32'sd3884205, -32'sd4132229, -32'sd2145905, -32'sd2266972, -32'sd1509706, -32'sd970837, -32'sd942728, -32'sd945036, -32'sd3054145, -32'sd1353548, 32'sd1044764, 32'sd454598, -32'sd178501, 32'sd411259, 32'sd1302784, 32'sd974651, 32'sd1863592, -32'sd896180, 32'sd45410, -32'sd957109, 32'sd414647, -32'sd636167, 32'sd999759, -32'sd1557998, 32'sd1334629, 32'sd322604, -32'sd1660116, -32'sd4963243, -32'sd4829057, -32'sd5969778, -32'sd2230303, -32'sd1879900, -32'sd1595168, 32'sd586094, -32'sd1792913, -32'sd1774182, -32'sd2633193, -32'sd499616, 32'sd119890, 32'sd996702, -32'sd1239707, 32'sd867688, 32'sd517870, 32'sd497567, -32'sd1212943, -32'sd390253, 32'sd1251852, -32'sd243195, 32'sd851708, -32'sd1567795, -32'sd1015076, -32'sd1953981, -32'sd1465252, -32'sd1965727, -32'sd1670368, -32'sd2734805, -32'sd3411868, -32'sd4230623, -32'sd3849578, -32'sd689419, -32'sd422805, 32'sd970804, -32'sd2699777, -32'sd2517460, -32'sd2887505, -32'sd932897, 32'sd485238, -32'sd243138, 32'sd919262, 32'sd1968960, 32'sd512678, -32'sd739539, -32'sd234734, 32'sd0, -32'sd504836, 32'sd1761729, -32'sd405011, 32'sd1640998, 32'sd893574, -32'sd2116885, -32'sd58283, -32'sd2345773, -32'sd1911835, -32'sd2396431, -32'sd4073589, -32'sd2101624, -32'sd1028525, -32'sd2383101, -32'sd1305586, 32'sd1962126, -32'sd1335454, -32'sd1744240, -32'sd919690, 32'sd548420, -32'sd22643, 32'sd412251, 32'sd1831510, 32'sd2341882, 32'sd805396, -32'sd928100, 32'sd880961, -32'sd399078, 32'sd283802, -32'sd542488, 32'sd521354, -32'sd130947, 32'sd1758186, 32'sd370772, 32'sd48910, -32'sd723061, 32'sd262476, -32'sd1189223, -32'sd3225668, -32'sd1197184, -32'sd276012, -32'sd3499031, -32'sd2037415, 32'sd1583560, -32'sd1313810, 32'sd146513, -32'sd752811, -32'sd734518, 32'sd1364903, 32'sd391348, 32'sd1684359, 32'sd286400, -32'sd2712331, -32'sd54561, -32'sd985697, -32'sd703338, -32'sd762446, -32'sd17354, 32'sd462303, -32'sd694683, 32'sd1420174, 32'sd1114516, 32'sd1838268, 32'sd113403, 32'sd151453, -32'sd1013721, 32'sd830392, -32'sd1661006, 32'sd146177, 32'sd320804, -32'sd2691, 32'sd462256, -32'sd302247, 32'sd1120511, 32'sd781972, 32'sd1241592, 32'sd482548, -32'sd477983, 32'sd16078, 32'sd399219, -32'sd1947984, 32'sd116474, -32'sd585971, 32'sd0, 32'sd364133, -32'sd1551871, -32'sd90151, 32'sd824308, 32'sd351450, 32'sd1356652, 32'sd2463707, 32'sd1770874, 32'sd1618701, 32'sd1704785, 32'sd1723378, -32'sd1345114, -32'sd296793, 32'sd1228632, 32'sd1823481, 32'sd1781850, 32'sd864921, 32'sd1471790, 32'sd573326, 32'sd1239736, 32'sd1601102, -32'sd117494, 32'sd173022, 32'sd97626, -32'sd151296, 32'sd332373, -32'sd480173, -32'sd564629, -32'sd339539, -32'sd105113, -32'sd382044, 32'sd791017, -32'sd740528, -32'sd163282, 32'sd963654, 32'sd978465, -32'sd452412, 32'sd1126793, 32'sd2192222, -32'sd1424111, 32'sd135240, 32'sd3001203, 32'sd575303, 32'sd2214743, 32'sd2336175, 32'sd1489297, 32'sd942105, -32'sd1031622, -32'sd1383299, 32'sd636169, 32'sd1048259, -32'sd1756424, 32'sd728066, -32'sd1013199, 32'sd709910, 32'sd216023, -32'sd796373, -32'sd544051, -32'sd23390, -32'sd510919, 32'sd885323, 32'sd260527, -32'sd570409, 32'sd498281, -32'sd323625, 32'sd1027331, 32'sd982957, 32'sd2188487, 32'sd153138, 32'sd89775, 32'sd1927641, -32'sd685312, 32'sd1300540, 32'sd401916, 32'sd252916, 32'sd565207, -32'sd332624, 32'sd1993604, 32'sd1275563, 32'sd16176, -32'sd1095489, 32'sd44311, 32'sd666306, 32'sd0, -32'sd519764, 32'sd160947, -32'sd2288415, -32'sd30850, 32'sd93520, 32'sd346618, 32'sd1284299, -32'sd319684, 32'sd1073866, 32'sd1051555, 32'sd1900388, 32'sd842543, 32'sd641067, -32'sd1864934, 32'sd2836886, 32'sd1542021, 32'sd36417, 32'sd209798, -32'sd2525539, -32'sd652451, -32'sd771615, -32'sd1516436, 32'sd1526995, 32'sd1358829, -32'sd172783, -32'sd350657, 32'sd0, 32'sd0, 32'sd0, -32'sd29629, 32'sd44476, 32'sd831469, -32'sd209780, -32'sd243314, 32'sd2567045, 32'sd675402, 32'sd2032179, 32'sd191579, 32'sd502274, -32'sd21962, -32'sd1333219, 32'sd463496, 32'sd1955328, -32'sd271872, 32'sd851262, 32'sd901862, -32'sd739320, -32'sd2659495, -32'sd17032, -32'sd343343, 32'sd149333, 32'sd279658, -32'sd1299252, 32'sd1126243, 32'sd0, 32'sd0, 32'sd0, -32'sd206954, -32'sd16724, -32'sd1116713, 32'sd202712, -32'sd698399, 32'sd911065, 32'sd366162, 32'sd2709373, 32'sd542809, 32'sd2175179, 32'sd2618434, 32'sd1405501, 32'sd988253, 32'sd1659962, 32'sd196280, 32'sd367376, 32'sd813461, 32'sd2181970, 32'sd1387164, 32'sd1621704, 32'sd433742, 32'sd625747, 32'sd1341062, -32'sd89450, -32'sd195766, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd252385, 32'sd490321, -32'sd454475, 32'sd909993, 32'sd741301, -32'sd281343, -32'sd1470980, 32'sd1001562, 32'sd591224, 32'sd1602388, 32'sd715385, 32'sd279744, 32'sd1669854, 32'sd2208978, 32'sd1179368, 32'sd311621, 32'sd1490022, 32'sd293076, 32'sd550393, 32'sd695893, 32'sd596234, -32'sd1471921, 32'sd1028163, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd293923, -32'sd1021666, -32'sd377345, -32'sd247756, 32'sd1816156, 32'sd842391, 32'sd1403411, -32'sd1157667, 32'sd970420, 32'sd586361, -32'sd713730, -32'sd1492913, -32'sd1139718, -32'sd146771, 32'sd545933, 32'sd1203604, 32'sd28759, 32'sd443989, 32'sd1060512, 32'sd259518, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1023125, -32'sd35134, 32'sd255376, -32'sd54238, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd540954, 32'sd294005, -32'sd335819, -32'sd757827, -32'sd1323168, 32'sd81040, 32'sd478580, 32'sd1770273, 32'sd323732, 32'sd289647, 32'sd416818, 32'sd890654, -32'sd361379, 32'sd1484344, -32'sd5231, 32'sd1336190, 32'sd1072825, 32'sd832805, 32'sd1231746, 32'sd100017, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd379910, 32'sd155428, 32'sd1336603, -32'sd399121, 32'sd547600, -32'sd933410, -32'sd412468, -32'sd915607, -32'sd470423, 32'sd487955, 32'sd633491, 32'sd2968971, 32'sd647802, 32'sd1878857, 32'sd417421, 32'sd1723155, -32'sd531332, 32'sd405637, -32'sd85356, 32'sd903841, 32'sd1464624, 32'sd862276, 32'sd730571, 32'sd63587, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd267162, -32'sd944033, 32'sd1111572, 32'sd27968, 32'sd732243, 32'sd575726, -32'sd1930458, 32'sd417004, -32'sd1463310, -32'sd1177938, 32'sd2039990, 32'sd611384, 32'sd1893084, 32'sd600262, -32'sd476150, -32'sd114201, -32'sd799602, -32'sd2881353, -32'sd2198053, -32'sd1729386, -32'sd1600576, -32'sd2588459, -32'sd399484, -32'sd926381, 32'sd275556, 32'sd0, 32'sd0, -32'sd12140, 32'sd940952, 32'sd471019, -32'sd1764395, 32'sd13714, -32'sd30015, -32'sd1808425, -32'sd1155580, -32'sd1701529, -32'sd2767628, 32'sd2654310, 32'sd1709960, 32'sd1571797, -32'sd1322046, 32'sd1528819, -32'sd1688338, -32'sd207814, -32'sd158628, -32'sd1664466, -32'sd889266, -32'sd355881, 32'sd669728, 32'sd184690, 32'sd116472, -32'sd1193515, 32'sd477919, 32'sd374479, 32'sd0, 32'sd572495, 32'sd1009320, -32'sd635938, -32'sd1162561, -32'sd766175, -32'sd2582494, -32'sd2611742, -32'sd913463, -32'sd393324, 32'sd603264, 32'sd2022451, 32'sd1695066, 32'sd671477, 32'sd1706052, 32'sd1488678, -32'sd872994, -32'sd2422903, 32'sd146379, -32'sd917403, -32'sd2255195, 32'sd538489, 32'sd883713, -32'sd867009, 32'sd1750635, -32'sd1226924, 32'sd807846, -32'sd303876, 32'sd0, -32'sd163969, 32'sd53774, 32'sd135855, -32'sd661803, -32'sd431401, -32'sd3590398, -32'sd2260409, -32'sd791709, -32'sd1862061, -32'sd2316110, 32'sd1277135, -32'sd102887, 32'sd2594414, 32'sd1318811, -32'sd1420725, -32'sd2156925, -32'sd2347707, -32'sd72906, 32'sd78805, -32'sd230234, 32'sd1614058, 32'sd2239802, 32'sd1347033, 32'sd2867818, 32'sd2231639, 32'sd1985360, 32'sd1339617, 32'sd185399, 32'sd490283, 32'sd45948, 32'sd161, -32'sd64123, -32'sd99536, -32'sd1509330, -32'sd1014960, -32'sd4298615, -32'sd3663648, -32'sd106827, 32'sd3236452, 32'sd2119841, 32'sd2241789, -32'sd1689788, -32'sd103271, 32'sd1030039, 32'sd216309, 32'sd2511065, 32'sd1961784, 32'sd2324614, 32'sd2207282, 32'sd2221349, 32'sd2185376, 32'sd1971718, 32'sd2397353, 32'sd256457, -32'sd509790, 32'sd827620, -32'sd147435, -32'sd1659220, 32'sd357511, -32'sd820318, 32'sd1510168, -32'sd1009702, -32'sd1134831, -32'sd4381765, -32'sd195890, -32'sd310615, 32'sd2365082, 32'sd2989483, 32'sd322385, 32'sd250749, 32'sd1204071, -32'sd384195, 32'sd2158994, 32'sd2407347, 32'sd1013312, -32'sd620808, 32'sd933481, 32'sd1021149, -32'sd1065061, 32'sd737522, -32'sd1247926, -32'sd562920, -32'sd974784, 32'sd1778242, -32'sd475809, -32'sd684778, -32'sd431484, 32'sd769854, 32'sd1267348, -32'sd1222868, -32'sd3145199, -32'sd2869193, 32'sd844466, -32'sd1008962, 32'sd1953057, 32'sd1946718, 32'sd575413, -32'sd2415026, -32'sd470873, -32'sd122738, -32'sd2580025, -32'sd951810, -32'sd2307801, -32'sd1493827, -32'sd1776109, -32'sd701216, -32'sd875693, -32'sd1340777, -32'sd2144471, -32'sd767672, 32'sd402907, -32'sd189962, 32'sd885905, 32'sd69149, -32'sd465351, -32'sd778889, 32'sd1209045, 32'sd334049, -32'sd1618087, -32'sd3278710, -32'sd546024, 32'sd1262891, 32'sd3157659, 32'sd1200685, -32'sd485661, -32'sd939572, -32'sd2119486, -32'sd3017310, -32'sd1601385, -32'sd1506239, -32'sd2922957, -32'sd4219682, -32'sd1235544, -32'sd268464, -32'sd1501598, -32'sd511499, -32'sd250264, -32'sd1174823, -32'sd1326981, 32'sd275869, -32'sd1445210, -32'sd1445043, -32'sd825426, -32'sd200865, 32'sd13271, -32'sd857845, -32'sd124940, -32'sd3057572, -32'sd1510153, 32'sd133723, 32'sd502633, -32'sd147794, -32'sd1026449, -32'sd530970, -32'sd4220424, -32'sd499644, -32'sd122224, -32'sd1321514, -32'sd1114928, -32'sd2799480, -32'sd61525, 32'sd780409, 32'sd1217479, 32'sd1938677, -32'sd1493413, 32'sd1052473, -32'sd841189, 32'sd705284, -32'sd795326, 32'sd817437, -32'sd1535330, 32'sd303388, 32'sd201416, 32'sd546422, -32'sd1723816, -32'sd667308, 32'sd36842, -32'sd231476, 32'sd1759008, -32'sd678728, -32'sd677777, -32'sd595855, -32'sd1111666, -32'sd3189699, 32'sd229948, 32'sd1545023, 32'sd308897, -32'sd1851931, -32'sd1130464, -32'sd1052649, 32'sd1119695, 32'sd446356, 32'sd1486982, 32'sd1628369, 32'sd586731, 32'sd723151, -32'sd99259, -32'sd751513, -32'sd587937, 32'sd773996, 32'sd2127064, -32'sd682639, 32'sd864434, -32'sd1676271, -32'sd1702114, 32'sd387807, -32'sd1073940, -32'sd777562, -32'sd1205913, 32'sd647047, -32'sd160519, -32'sd1342886, -32'sd1386411, -32'sd923675, 32'sd1573715, 32'sd1010206, 32'sd407589, 32'sd180071, 32'sd676847, -32'sd724384, 32'sd790170, 32'sd712153, -32'sd827150, 32'sd577455, 32'sd1338145, 32'sd771492, -32'sd220322, 32'sd524893, 32'sd490262, -32'sd867756, 32'sd1457399, -32'sd603011, 32'sd1007303, -32'sd159416, -32'sd1631302, -32'sd1020292, -32'sd628408, 32'sd236997, 32'sd1979812, 32'sd659511, 32'sd777393, -32'sd286886, -32'sd133669, -32'sd447472, 32'sd591697, 32'sd1902916, 32'sd1599570, -32'sd544382, 32'sd1512900, 32'sd209142, 32'sd502498, 32'sd1870810, -32'sd1117713, -32'sd1508061, 32'sd670238, -32'sd364576, 32'sd1560247, -32'sd1524745, -32'sd1725163, -32'sd1362619, 32'sd490909, 32'sd1276815, 32'sd854858, 32'sd1745426, -32'sd1678473, -32'sd1181886, 32'sd1220419, -32'sd901558, 32'sd1518271, 32'sd559143, -32'sd2594024, -32'sd800739, 32'sd931166, 32'sd2344900, 32'sd698153, 32'sd633163, 32'sd407713, -32'sd112522, 32'sd411614, 32'sd299240, -32'sd280427, 32'sd1098139, 32'sd684992, 32'sd1046183, 32'sd1264799, -32'sd404974, 32'sd718417, -32'sd952747, -32'sd1458569, -32'sd153440, 32'sd1506617, 32'sd18891, -32'sd1340324, -32'sd1084270, -32'sd1403940, -32'sd700692, -32'sd744964, -32'sd252431, -32'sd1880580, -32'sd848962, 32'sd801289, 32'sd1836876, 32'sd282212, -32'sd616528, -32'sd424401, -32'sd1185897, 32'sd206956, 32'sd0, -32'sd74897, 32'sd1057726, -32'sd26436, 32'sd342741, 32'sd559423, -32'sd1065587, -32'sd1364136, -32'sd385724, -32'sd1963181, -32'sd86779, 32'sd475960, -32'sd629993, -32'sd146731, -32'sd590446, -32'sd2557615, 32'sd489623, 32'sd609417, -32'sd662844, -32'sd2794797, -32'sd165661, 32'sd177134, 32'sd1253914, -32'sd176744, -32'sd456329, -32'sd730491, -32'sd203845, 32'sd1436346, 32'sd945372, -32'sd513590, -32'sd272389, 32'sd518200, 32'sd1084853, 32'sd913902, 32'sd294351, 32'sd636677, -32'sd798250, -32'sd1564888, -32'sd2799273, -32'sd2352422, -32'sd1108681, -32'sd2832726, -32'sd1715784, -32'sd738053, 32'sd1040916, 32'sd904851, -32'sd1736030, 32'sd134172, 32'sd433775, 32'sd884732, -32'sd577995, 32'sd365408, -32'sd1837265, -32'sd116124, -32'sd881174, -32'sd587518, 32'sd949019, 32'sd399884, -32'sd816621, -32'sd1196475, -32'sd499258, -32'sd82918, 32'sd264577, 32'sd448537, 32'sd1056172, -32'sd1149951, -32'sd2556100, -32'sd2518639, -32'sd1490664, -32'sd1520919, 32'sd1769918, 32'sd2162027, 32'sd2432231, 32'sd360734, 32'sd1520990, -32'sd1304446, 32'sd545894, -32'sd1745295, 32'sd117060, -32'sd569227, -32'sd1206807, 32'sd2123731, -32'sd1953535, 32'sd10443, 32'sd0, 32'sd649441, 32'sd315112, -32'sd674640, -32'sd1909955, -32'sd579573, 32'sd577534, -32'sd925221, 32'sd1292820, 32'sd188861, 32'sd244987, -32'sd846707, 32'sd548140, -32'sd507108, 32'sd1943684, 32'sd1153099, -32'sd74022, 32'sd948369, 32'sd1337586, -32'sd226522, -32'sd863022, -32'sd2160763, 32'sd840177, -32'sd341583, -32'sd99314, 32'sd795801, -32'sd1566919, 32'sd747437, 32'sd1585509, -32'sd1266730, 32'sd548577, -32'sd273852, -32'sd2051918, -32'sd755311, 32'sd671084, 32'sd1538157, -32'sd76397, -32'sd886387, -32'sd188660, 32'sd719618, 32'sd1113545, 32'sd827614, 32'sd676048, -32'sd1341753, 32'sd551783, -32'sd393988, 32'sd71947, -32'sd1039879, -32'sd74044, 32'sd507504, 32'sd132120, -32'sd1704743, 32'sd589316, 32'sd71370, -32'sd2074088, 32'sd1260618, 32'sd1248765, 32'sd1455829, -32'sd179195, -32'sd187357, 32'sd419723, -32'sd2311933, 32'sd983879, -32'sd1164802, 32'sd839927, 32'sd228194, 32'sd1180357, 32'sd1542611, 32'sd74237, 32'sd881498, 32'sd474105, 32'sd725223, 32'sd1337236, -32'sd298068, -32'sd1157089, 32'sd717123, -32'sd487440, -32'sd625023, -32'sd599177, 32'sd1033009, 32'sd42478, -32'sd51663, 32'sd123094, 32'sd477257, 32'sd0, -32'sd22891, 32'sd207521, -32'sd900879, 32'sd191420, -32'sd1449101, -32'sd1042084, -32'sd625034, -32'sd2815775, -32'sd181782, -32'sd926668, 32'sd1175597, 32'sd2296617, 32'sd1519728, 32'sd2048696, 32'sd840997, 32'sd124005, 32'sd205881, -32'sd68596, 32'sd250914, 32'sd790170, 32'sd1915237, 32'sd1415487, -32'sd50958, 32'sd1157567, 32'sd626952, 32'sd797900, 32'sd0, 32'sd0, 32'sd0, 32'sd542427, -32'sd1452526, 32'sd767552, 32'sd57692, 32'sd457065, -32'sd1065645, -32'sd1477405, 32'sd532397, -32'sd3312869, -32'sd978245, 32'sd918081, 32'sd1076915, 32'sd1312464, -32'sd1588357, 32'sd1049621, -32'sd741965, 32'sd552498, 32'sd892020, 32'sd2605787, 32'sd1190713, -32'sd70706, -32'sd1341589, -32'sd961811, 32'sd668387, 32'sd482568, 32'sd0, 32'sd0, 32'sd0, 32'sd1077247, -32'sd1704775, 32'sd553578, -32'sd2069821, 32'sd672790, -32'sd1272317, 32'sd1041507, 32'sd457082, 32'sd1264948, -32'sd423512, -32'sd225451, 32'sd1626279, 32'sd599630, -32'sd2409059, -32'sd921005, -32'sd2582645, 32'sd1048533, 32'sd2484219, -32'sd59487, -32'sd781726, -32'sd808202, -32'sd963686, -32'sd718444, -32'sd1136290, -32'sd18148, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd241125, 32'sd120420, -32'sd943674, -32'sd1590398, -32'sd1479492, 32'sd2499255, 32'sd1109944, -32'sd994403, 32'sd2953276, 32'sd2060384, -32'sd2217251, -32'sd1799072, 32'sd566414, 32'sd399133, -32'sd691081, 32'sd1224700, 32'sd1547308, 32'sd1305039, 32'sd792666, 32'sd2256398, -32'sd1452026, -32'sd117753, 32'sd24873, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd12187, 32'sd155325, 32'sd414847, 32'sd586791, -32'sd250392, 32'sd43666, 32'sd604464, -32'sd332297, -32'sd1409629, 32'sd1773866, -32'sd345392, 32'sd446277, 32'sd366431, 32'sd1160308, 32'sd333151, -32'sd45947, -32'sd292890, -32'sd922026, -32'sd1948635, 32'sd109958, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd828969, 32'sd531998, 32'sd367609, 32'sd317837, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd227751, -32'sd480100, -32'sd1753946, -32'sd123373, 32'sd502838, -32'sd1384940, -32'sd312537, -32'sd626149, -32'sd844300, -32'sd99082, 32'sd1370029, 32'sd1707003, 32'sd243103, -32'sd733635, 32'sd185831, 32'sd13111, -32'sd1468989, -32'sd504192, -32'sd225316, -32'sd110230, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd198830, 32'sd467266, -32'sd751971, 32'sd1069338, -32'sd338081, 32'sd856184, 32'sd371100, -32'sd285419, 32'sd1625731, -32'sd1250679, 32'sd545695, 32'sd636611, 32'sd1193894, 32'sd2475391, 32'sd3155470, 32'sd1036938, 32'sd1635000, 32'sd438876, -32'sd475980, 32'sd596042, -32'sd1434044, -32'sd168438, -32'sd1022402, 32'sd144469, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd853855, -32'sd350196, -32'sd390677, -32'sd406800, 32'sd1601491, -32'sd728641, -32'sd821561, -32'sd127502, 32'sd1113748, -32'sd153421, 32'sd1995924, 32'sd1141855, 32'sd1774702, -32'sd33875, -32'sd276719, 32'sd1959354, 32'sd1052406, 32'sd2633375, -32'sd424663, -32'sd939296, 32'sd14336, -32'sd1861631, 32'sd349827, -32'sd949810, 32'sd462888, 32'sd0, 32'sd0, 32'sd1138130, 32'sd1108030, -32'sd293202, -32'sd1077838, 32'sd759391, 32'sd826728, -32'sd927931, -32'sd1206326, -32'sd1113835, -32'sd2029799, 32'sd299719, -32'sd1979243, -32'sd56494, -32'sd95090, -32'sd384519, -32'sd249932, -32'sd1226895, 32'sd314942, -32'sd58122, 32'sd777219, 32'sd695352, 32'sd357062, 32'sd65711, -32'sd644843, -32'sd1727684, -32'sd1309601, 32'sd363679, 32'sd0, 32'sd316952, 32'sd309968, 32'sd117826, -32'sd649751, -32'sd2248638, -32'sd2667612, -32'sd134524, -32'sd2359494, -32'sd1394179, -32'sd2936117, -32'sd4352992, -32'sd1880067, -32'sd2298015, 32'sd438264, -32'sd374817, 32'sd1062713, -32'sd136483, 32'sd847416, 32'sd979697, 32'sd370313, 32'sd1319510, 32'sd2358836, 32'sd2961423, -32'sd166312, -32'sd2442472, -32'sd1852856, -32'sd939908, 32'sd0, -32'sd794363, -32'sd49429, -32'sd151909, 32'sd298196, -32'sd3239479, 32'sd410941, 32'sd854499, -32'sd2123230, 32'sd1419390, 32'sd1989308, -32'sd774613, -32'sd417648, 32'sd6417, 32'sd956054, 32'sd2098825, 32'sd1397888, 32'sd754817, 32'sd163717, 32'sd1091456, -32'sd1140438, -32'sd764289, -32'sd1262511, -32'sd247450, -32'sd838661, -32'sd1517168, -32'sd1465618, 32'sd581352, 32'sd219713, 32'sd839412, 32'sd1060163, 32'sd1062132, 32'sd258243, -32'sd1717183, -32'sd503022, 32'sd101169, -32'sd1197773, -32'sd190702, 32'sd772375, 32'sd1725507, 32'sd1438290, 32'sd1351303, 32'sd3314640, 32'sd2454423, 32'sd1095006, 32'sd1550349, -32'sd1162969, 32'sd355138, -32'sd919705, 32'sd1073503, 32'sd870180, -32'sd309581, -32'sd912076, -32'sd2423486, -32'sd680633, 32'sd407507, 32'sd210830, -32'sd1885424, 32'sd1065949, 32'sd33984, -32'sd209405, -32'sd1009317, -32'sd1724217, 32'sd1260509, 32'sd1619232, 32'sd474748, 32'sd2278202, 32'sd3611028, 32'sd2675507, 32'sd2319293, 32'sd2329133, 32'sd1774181, 32'sd1599912, 32'sd1210959, 32'sd1693706, 32'sd1714105, 32'sd636690, 32'sd1549700, 32'sd466535, -32'sd439973, -32'sd3298521, -32'sd1277151, -32'sd345130, -32'sd844081, -32'sd291143, 32'sd1329783, -32'sd763264, -32'sd1175370, -32'sd1230810, -32'sd395260, 32'sd3288420, 32'sd1180155, 32'sd3025544, 32'sd2529334, 32'sd2958933, 32'sd329896, 32'sd1359609, -32'sd632812, -32'sd1445503, -32'sd303728, 32'sd1397111, 32'sd274030, 32'sd1405785, 32'sd2173918, 32'sd99303, -32'sd535460, 32'sd589139, 32'sd182765, -32'sd890577, -32'sd1167512, -32'sd835270, -32'sd547553, -32'sd85342, -32'sd521194, -32'sd342155, 32'sd1593978, 32'sd51010, 32'sd66321, 32'sd2745520, 32'sd1815161, 32'sd2527370, -32'sd249122, -32'sd1331119, -32'sd1217511, -32'sd1394011, -32'sd2790490, -32'sd6201663, -32'sd1581700, 32'sd521520, 32'sd993632, 32'sd2351630, 32'sd2144300, 32'sd360959, 32'sd1319307, 32'sd167369, -32'sd973457, -32'sd1629450, -32'sd25173, 32'sd222434, -32'sd433368, -32'sd332067, -32'sd397337, 32'sd971576, 32'sd1516582, 32'sd718613, -32'sd384157, 32'sd1137198, -32'sd475113, -32'sd2407664, -32'sd833472, -32'sd2902602, -32'sd4296885, -32'sd5588164, -32'sd5019255, -32'sd4107943, -32'sd1021482, -32'sd628566, 32'sd2118410, 32'sd3865743, 32'sd1527181, 32'sd669836, 32'sd1931179, 32'sd1199109, -32'sd2745436, -32'sd4036, 32'sd145359, -32'sd652616, -32'sd1067021, 32'sd536679, 32'sd541464, -32'sd1421466, -32'sd120498, 32'sd1349373, -32'sd2552682, -32'sd2100612, -32'sd1951238, -32'sd2497668, -32'sd3357653, -32'sd4138742, -32'sd6034428, -32'sd2853437, -32'sd5479683, 32'sd850868, 32'sd3428740, 32'sd1598753, 32'sd1905497, 32'sd546983, 32'sd1249866, -32'sd1170636, -32'sd1011652, -32'sd1797715, 32'sd94756, -32'sd1965034, -32'sd2667228, -32'sd583766, 32'sd884227, 32'sd243018, -32'sd1307008, -32'sd717225, 32'sd875992, -32'sd2959654, -32'sd2947016, -32'sd3637438, -32'sd1156593, -32'sd374046, -32'sd3921903, -32'sd2024081, -32'sd1634580, -32'sd776316, -32'sd614801, 32'sd1050214, 32'sd182685, 32'sd1032767, 32'sd1648357, 32'sd648763, 32'sd125056, -32'sd1426091, -32'sd1188490, -32'sd2637460, -32'sd1914697, -32'sd1611885, -32'sd1393060, -32'sd1219271, -32'sd874219, 32'sd265496, -32'sd352938, 32'sd286886, 32'sd248132, -32'sd2074982, -32'sd2514256, -32'sd332391, 32'sd810418, 32'sd393900, -32'sd2833465, -32'sd650463, 32'sd2202138, 32'sd1029598, 32'sd2060681, 32'sd1454562, 32'sd3053073, 32'sd1981161, 32'sd141758, 32'sd941719, -32'sd917663, 32'sd1159655, 32'sd356766, -32'sd2155788, -32'sd1306329, 32'sd467945, -32'sd114367, 32'sd697050, -32'sd360112, -32'sd813848, -32'sd583645, -32'sd531934, -32'sd566859, -32'sd986353, -32'sd6593, 32'sd1856744, 32'sd1695443, 32'sd1627802, 32'sd197364, 32'sd1181434, 32'sd1135348, 32'sd1647371, -32'sd103482, 32'sd1013892, 32'sd634731, 32'sd858107, -32'sd603529, -32'sd371749, 32'sd713721, -32'sd1715597, -32'sd1521158, -32'sd2446559, 32'sd850044, -32'sd1713260, -32'sd378995, 32'sd807843, -32'sd1038725, 32'sd463153, 32'sd1655388, 32'sd1555276, -32'sd145322, -32'sd359389, -32'sd165058, 32'sd1136403, 32'sd847422, -32'sd535403, -32'sd627805, -32'sd256817, -32'sd226482, -32'sd347658, 32'sd44033, 32'sd210842, 32'sd1796299, -32'sd582331, -32'sd1105490, 32'sd920434, -32'sd503584, -32'sd2267091, -32'sd1237128, -32'sd2639511, -32'sd650777, 32'sd724932, -32'sd496308, -32'sd2047523, -32'sd968806, 32'sd0, 32'sd408022, 32'sd1248227, -32'sd822906, 32'sd1080645, 32'sd586616, -32'sd405893, 32'sd193957, -32'sd407820, -32'sd1739033, 32'sd747590, -32'sd172872, 32'sd857444, 32'sd723524, 32'sd4248507, 32'sd3325608, 32'sd493324, -32'sd830450, -32'sd508891, 32'sd1515213, -32'sd389715, -32'sd2526272, -32'sd2335988, -32'sd181718, 32'sd436773, 32'sd558560, -32'sd614947, -32'sd383034, 32'sd184362, 32'sd552774, 32'sd1483986, 32'sd172100, -32'sd135042, -32'sd429027, -32'sd3946, -32'sd1786094, -32'sd829803, 32'sd858932, 32'sd720933, 32'sd1376207, 32'sd228631, 32'sd644952, 32'sd539544, 32'sd634004, 32'sd1966899, 32'sd1496464, 32'sd287105, 32'sd1348969, -32'sd467696, -32'sd941891, 32'sd198460, -32'sd1560994, 32'sd973434, -32'sd1268767, -32'sd596948, 32'sd1122676, 32'sd279166, -32'sd797376, -32'sd898007, -32'sd34240, 32'sd1497052, 32'sd31059, 32'sd2083227, 32'sd640150, 32'sd802954, -32'sd508376, 32'sd1147290, -32'sd56385, 32'sd714565, 32'sd2648130, -32'sd535264, 32'sd349393, 32'sd1415215, 32'sd8079, -32'sd69300, 32'sd1695863, -32'sd254961, -32'sd399800, -32'sd565902, -32'sd1124264, 32'sd154139, -32'sd523859, 32'sd1295306, 32'sd600676, 32'sd0, -32'sd436125, -32'sd33611, -32'sd940883, 32'sd1150358, -32'sd570718, -32'sd227872, 32'sd2210592, 32'sd1386844, 32'sd1063541, 32'sd2120718, 32'sd35584, 32'sd1319306, -32'sd463853, 32'sd1207517, -32'sd232648, -32'sd446758, -32'sd570616, 32'sd1803961, 32'sd2049778, -32'sd956139, 32'sd335352, 32'sd574047, -32'sd158113, -32'sd1121951, -32'sd883295, -32'sd148105, 32'sd295436, 32'sd1462707, -32'sd575041, -32'sd466694, 32'sd1117365, 32'sd2177845, -32'sd127140, 32'sd54918, -32'sd291803, -32'sd965731, 32'sd142622, 32'sd274993, 32'sd249105, 32'sd336458, -32'sd347565, 32'sd52074, -32'sd481873, -32'sd59987, -32'sd395979, 32'sd527988, 32'sd492100, 32'sd1875043, 32'sd1895776, -32'sd1173, -32'sd2587067, -32'sd427177, -32'sd1116943, -32'sd324526, -32'sd370321, -32'sd51247, -32'sd1097602, -32'sd312360, -32'sd946983, 32'sd337494, -32'sd450295, 32'sd47550, 32'sd128686, -32'sd1272522, -32'sd1478097, -32'sd1994153, -32'sd1001858, -32'sd1786431, -32'sd1897611, -32'sd1212669, -32'sd636482, 32'sd1937527, 32'sd134172, 32'sd899365, 32'sd2242163, 32'sd363530, 32'sd1204672, -32'sd660756, 32'sd9343, -32'sd257044, -32'sd1371187, 32'sd54904, 32'sd461526, 32'sd0, -32'sd124481, -32'sd31567, -32'sd1651825, -32'sd1458955, 32'sd747464, -32'sd548838, 32'sd1355365, 32'sd353689, -32'sd416045, 32'sd679435, -32'sd739272, -32'sd2159464, 32'sd1192923, -32'sd1531782, 32'sd414351, -32'sd415027, -32'sd1405564, 32'sd30106, 32'sd1294853, -32'sd1354883, 32'sd728698, -32'sd145860, 32'sd485849, 32'sd88859, -32'sd488649, 32'sd847643, 32'sd0, 32'sd0, 32'sd0, 32'sd101246, 32'sd480155, -32'sd153053, 32'sd740516, -32'sd683484, -32'sd1539594, -32'sd842030, -32'sd906931, 32'sd825725, 32'sd770564, -32'sd1760504, -32'sd529862, 32'sd726577, -32'sd927470, -32'sd52221, 32'sd505729, -32'sd356636, 32'sd585794, 32'sd694243, 32'sd271416, -32'sd85380, -32'sd393359, 32'sd629905, -32'sd1031514, 32'sd45563, 32'sd0, 32'sd0, 32'sd0, -32'sd306989, -32'sd463704, 32'sd801093, 32'sd601746, -32'sd351543, 32'sd618333, 32'sd311376, 32'sd1047388, -32'sd998013, -32'sd1406624, 32'sd1196982, -32'sd686594, -32'sd673444, -32'sd1054707, -32'sd138804, -32'sd1438263, -32'sd149825, -32'sd413367, 32'sd691316, 32'sd689012, -32'sd1085055, 32'sd184013, 32'sd618117, -32'sd227520, 32'sd306917, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd136573, -32'sd599204, -32'sd482390, -32'sd899038, -32'sd528507, -32'sd1628411, -32'sd342759, 32'sd44458, -32'sd200016, -32'sd966604, -32'sd1074235, -32'sd1916479, -32'sd318984, -32'sd833019, -32'sd1106530, -32'sd2456947, -32'sd54730, 32'sd817414, 32'sd1505085, 32'sd835235, -32'sd1347717, 32'sd317667, 32'sd802168, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd97073, 32'sd972641, 32'sd1289774, 32'sd475656, 32'sd454302, -32'sd79549, 32'sd1520767, -32'sd13536, -32'sd353714, 32'sd1512039, -32'sd724665, 32'sd1008666, 32'sd1521426, -32'sd438737, -32'sd99942, 32'sd338827, 32'sd2009915, 32'sd105004, 32'sd137433, -32'sd643672, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd177173, 32'sd850602, 32'sd1563741, 32'sd927146, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd63339, 32'sd29916, -32'sd852574, 32'sd591701, -32'sd181629, 32'sd169676, 32'sd377772, 32'sd1120429, -32'sd1390438, 32'sd1079458, 32'sd1962565, 32'sd1812517, -32'sd557413, -32'sd670504, 32'sd790181, -32'sd373167, 32'sd1136829, 32'sd747169, -32'sd259533, 32'sd212754, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd26467, 32'sd1108589, 32'sd5769, -32'sd784962, 32'sd284821, -32'sd1573092, 32'sd1466802, 32'sd988604, 32'sd1818494, -32'sd276871, 32'sd234264, -32'sd790714, 32'sd258454, 32'sd688141, -32'sd1134659, 32'sd1406032, -32'sd334581, -32'sd23040, 32'sd1211402, 32'sd898728, 32'sd257650, 32'sd1541470, -32'sd1291526, 32'sd514897, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd173342, -32'sd300164, 32'sd8382, 32'sd1891629, 32'sd1038605, 32'sd1042067, 32'sd1522773, 32'sd717206, -32'sd221332, -32'sd1597178, -32'sd1458026, -32'sd640383, -32'sd1819586, -32'sd2847028, -32'sd3052999, -32'sd2074393, 32'sd1176567, -32'sd352171, -32'sd1250063, -32'sd1965084, -32'sd616880, -32'sd324764, -32'sd69902, -32'sd1655164, -32'sd86065, 32'sd0, 32'sd0, 32'sd749156, -32'sd360314, -32'sd56786, -32'sd2961154, -32'sd1502723, -32'sd2527568, -32'sd26326, -32'sd2083121, -32'sd2107888, -32'sd1877524, -32'sd3878147, -32'sd2800111, -32'sd3091041, -32'sd1459568, -32'sd2484241, -32'sd406945, 32'sd99361, -32'sd961789, -32'sd816958, -32'sd1223205, 32'sd2885347, 32'sd952075, 32'sd619516, 32'sd1403491, 32'sd588468, -32'sd166855, 32'sd28253, 32'sd0, 32'sd350588, -32'sd436477, -32'sd1339626, 32'sd970063, -32'sd1421768, -32'sd1018001, -32'sd2146761, -32'sd1041686, -32'sd2118181, -32'sd1622376, -32'sd1388162, -32'sd1796389, -32'sd3777902, -32'sd934770, 32'sd368823, -32'sd1036936, -32'sd1094775, -32'sd1124555, -32'sd1025349, 32'sd56500, 32'sd2222393, 32'sd216426, 32'sd935931, 32'sd696848, -32'sd361676, 32'sd1324932, 32'sd1102159, 32'sd0, 32'sd312324, -32'sd1867317, 32'sd687905, -32'sd683704, -32'sd833549, -32'sd2206493, -32'sd1801714, -32'sd2533076, -32'sd712409, 32'sd487979, -32'sd76815, 32'sd1150119, 32'sd278632, 32'sd1469557, 32'sd249768, -32'sd1646080, 32'sd611690, -32'sd3096358, -32'sd3392651, -32'sd2009355, -32'sd895827, -32'sd452201, 32'sd835117, 32'sd952954, 32'sd2106665, 32'sd2218047, -32'sd779247, 32'sd144615, 32'sd1333452, 32'sd45373, -32'sd402656, -32'sd51367, -32'sd752582, 32'sd231447, -32'sd1219546, -32'sd75434, 32'sd1638006, 32'sd1590385, 32'sd132079, 32'sd222982, 32'sd2148634, 32'sd1245441, -32'sd16698, -32'sd143633, -32'sd1681466, -32'sd2064103, -32'sd2908428, -32'sd3035525, -32'sd2828949, -32'sd919351, -32'sd1479026, 32'sd888444, 32'sd2488654, -32'sd31692, -32'sd656453, 32'sd29577, -32'sd928148, 32'sd1555455, 32'sd679707, 32'sd837013, 32'sd218459, -32'sd196012, 32'sd278734, 32'sd1336725, 32'sd2310984, 32'sd4728804, 32'sd2620577, 32'sd2669708, 32'sd1110928, 32'sd893859, 32'sd1154867, 32'sd503353, 32'sd695605, 32'sd1332124, 32'sd712785, -32'sd1614077, -32'sd1550003, -32'sd2460814, -32'sd817009, 32'sd840538, -32'sd203090, 32'sd528811, 32'sd358671, 32'sd1036726, -32'sd1168396, -32'sd112876, 32'sd297569, -32'sd313092, 32'sd1871433, 32'sd2538876, 32'sd1278541, 32'sd1640897, 32'sd4259313, 32'sd3973813, 32'sd2390056, 32'sd3851835, 32'sd2357115, 32'sd3444620, 32'sd1453953, 32'sd2533877, 32'sd942355, -32'sd150449, -32'sd598562, 32'sd344484, -32'sd1625158, -32'sd713901, 32'sd1879168, -32'sd672914, 32'sd1030684, 32'sd640144, -32'sd735570, 32'sd625171, -32'sd890384, 32'sd643487, -32'sd1322592, -32'sd101947, 32'sd229699, 32'sd2518963, 32'sd369558, 32'sd2605257, 32'sd3954417, 32'sd2144826, 32'sd2812270, 32'sd1377844, 32'sd1555717, 32'sd2027358, 32'sd2139299, 32'sd2638886, 32'sd1836176, -32'sd1157263, 32'sd693906, 32'sd368188, 32'sd726954, -32'sd1499584, -32'sd155203, 32'sd600103, 32'sd205202, -32'sd116646, 32'sd470004, -32'sd285560, -32'sd4218, 32'sd617038, 32'sd876202, 32'sd350421, 32'sd1063493, -32'sd548993, -32'sd241359, -32'sd1428896, -32'sd481180, 32'sd831732, -32'sd54359, 32'sd559434, 32'sd2632468, 32'sd3592370, 32'sd2627143, 32'sd1742884, 32'sd2162274, 32'sd519327, -32'sd2146974, -32'sd1422216, -32'sd1339623, -32'sd252229, 32'sd189313, -32'sd259737, 32'sd1236634, -32'sd1393793, -32'sd187411, 32'sd940881, 32'sd1046092, -32'sd1051207, 32'sd462221, 32'sd1132873, -32'sd1029472, -32'sd1019446, 32'sd33414, -32'sd1842203, -32'sd1804082, -32'sd3621148, -32'sd1444576, -32'sd846127, 32'sd606960, 32'sd1670468, 32'sd377594, 32'sd578475, -32'sd967775, -32'sd1136409, -32'sd1239598, -32'sd768309, -32'sd757234, -32'sd1697295, 32'sd452092, -32'sd1429824, -32'sd10466, 32'sd933447, 32'sd716480, 32'sd303675, 32'sd1011253, 32'sd240683, -32'sd802975, 32'sd384384, -32'sd1132519, -32'sd707996, -32'sd1293006, -32'sd156191, -32'sd3299853, -32'sd1917601, 32'sd1048091, 32'sd1134027, 32'sd1980298, 32'sd1943678, 32'sd82939, 32'sd822857, -32'sd1096206, 32'sd340556, -32'sd3004643, -32'sd1530301, -32'sd2035341, 32'sd280282, -32'sd894214, 32'sd1632720, 32'sd703570, -32'sd999289, -32'sd825770, -32'sd1360678, -32'sd713638, 32'sd840819, -32'sd911945, 32'sd992117, -32'sd2348188, -32'sd1232909, -32'sd2093309, 32'sd32888, -32'sd1739997, -32'sd745856, -32'sd450376, -32'sd901944, 32'sd312587, -32'sd1265383, -32'sd1154740, -32'sd2842370, -32'sd1023496, -32'sd1189488, -32'sd1696798, 32'sd391509, -32'sd232406, -32'sd1067668, 32'sd2021733, 32'sd1730308, -32'sd33023, 32'sd973743, 32'sd172389, 32'sd510906, -32'sd2207975, -32'sd1754974, -32'sd1284175, -32'sd607114, -32'sd1694926, -32'sd733917, -32'sd1605648, -32'sd580216, -32'sd67601, 32'sd196635, -32'sd478291, -32'sd2473048, -32'sd2535410, -32'sd1187043, -32'sd2165663, -32'sd920038, -32'sd589771, 32'sd625219, 32'sd827144, 32'sd858286, 32'sd680859, -32'sd317905, 32'sd310298, 32'sd1445557, 32'sd163656, 32'sd1125152, 32'sd82883, 32'sd554252, 32'sd736232, -32'sd966866, -32'sd1109910, -32'sd1156220, 32'sd598934, 32'sd1625671, -32'sd335926, 32'sd1661897, 32'sd1968638, 32'sd364654, -32'sd24735, -32'sd156002, -32'sd932099, -32'sd1239208, -32'sd1148716, -32'sd1401193, -32'sd167705, -32'sd606822, 32'sd708073, 32'sd1455814, 32'sd1440497, 32'sd2876926, 32'sd1198107, 32'sd2188305, -32'sd153745, 32'sd1309693, -32'sd333498, 32'sd0, -32'sd97400, -32'sd225360, -32'sd1290061, -32'sd726656, -32'sd1275719, 32'sd217713, 32'sd125063, -32'sd440845, -32'sd867209, -32'sd891743, -32'sd502317, 32'sd965545, 32'sd951413, -32'sd972143, -32'sd974420, -32'sd1118814, -32'sd521217, -32'sd780481, 32'sd2107068, 32'sd609339, 32'sd1642835, 32'sd2306687, 32'sd707046, 32'sd400405, 32'sd1914679, 32'sd1775934, -32'sd521966, -32'sd490227, -32'sd1311616, 32'sd401421, -32'sd289886, -32'sd202330, -32'sd1240764, -32'sd1501393, -32'sd408326, -32'sd1923041, 32'sd500263, 32'sd329635, 32'sd865891, -32'sd62675, -32'sd1389117, -32'sd1726818, -32'sd2521086, -32'sd1980055, 32'sd2112855, 32'sd1523640, 32'sd989328, 32'sd1064543, 32'sd335751, -32'sd168070, 32'sd193210, -32'sd874800, 32'sd226258, 32'sd1748442, 32'sd1450176, 32'sd612503, 32'sd595315, -32'sd148381, -32'sd618036, 32'sd384278, -32'sd135120, -32'sd3076741, -32'sd1598119, -32'sd273918, -32'sd1202522, -32'sd1140585, -32'sd1095613, -32'sd2402829, -32'sd3642383, -32'sd1280204, -32'sd1280607, -32'sd1054291, 32'sd975014, 32'sd2151329, 32'sd2583791, 32'sd2063322, 32'sd1073343, 32'sd310064, -32'sd1588289, -32'sd795682, -32'sd741916, 32'sd98264, 32'sd761565, 32'sd0, -32'sd623523, -32'sd1255352, -32'sd1607313, 32'sd317535, -32'sd200322, -32'sd2208172, -32'sd1385315, -32'sd2110862, -32'sd3561278, -32'sd2504439, -32'sd826516, -32'sd3374856, -32'sd3785390, -32'sd2419976, -32'sd2685632, -32'sd1014528, 32'sd1128517, 32'sd387454, 32'sd986886, 32'sd715526, 32'sd191071, 32'sd914941, 32'sd515087, 32'sd1090857, 32'sd2764905, 32'sd1201190, -32'sd189759, 32'sd141448, 32'sd36271, -32'sd1075320, -32'sd514519, 32'sd166390, 32'sd679395, -32'sd889265, -32'sd698189, -32'sd1148343, -32'sd889011, -32'sd381247, -32'sd988582, -32'sd420523, -32'sd1685163, -32'sd2868022, -32'sd2413665, 32'sd360602, 32'sd229266, 32'sd958095, 32'sd1424493, 32'sd860459, 32'sd124341, 32'sd497974, 32'sd1194421, 32'sd257029, 32'sd647789, -32'sd431729, 32'sd101504, 32'sd507009, 32'sd32037, -32'sd1465911, -32'sd968518, -32'sd130727, -32'sd615410, 32'sd429448, -32'sd392679, -32'sd2348716, -32'sd280233, -32'sd1778900, -32'sd1216088, -32'sd672426, 32'sd1148264, 32'sd1346321, -32'sd848339, 32'sd149544, -32'sd224675, -32'sd325757, 32'sd2139698, 32'sd928630, -32'sd399816, 32'sd1635157, -32'sd248214, -32'sd264170, 32'sd902542, -32'sd1386840, 32'sd945739, 32'sd0, 32'sd1024201, -32'sd266683, -32'sd518841, -32'sd1003006, 32'sd1868217, 32'sd1232799, -32'sd669106, -32'sd538713, -32'sd881515, -32'sd1682306, 32'sd1007916, -32'sd2051057, 32'sd423875, 32'sd836196, 32'sd1771300, -32'sd561665, -32'sd1049970, 32'sd1552019, -32'sd955003, 32'sd1046414, -32'sd912751, 32'sd1257484, 32'sd400124, 32'sd1132119, 32'sd227365, -32'sd246998, 32'sd0, 32'sd0, 32'sd0, -32'sd150459, -32'sd1114334, -32'sd1024195, 32'sd1194663, -32'sd1296276, -32'sd1096277, -32'sd440401, 32'sd480792, -32'sd806388, -32'sd1934044, -32'sd3302410, 32'sd984987, -32'sd325623, -32'sd1606980, -32'sd3144, -32'sd348483, 32'sd98265, 32'sd270319, 32'sd657813, -32'sd1470856, 32'sd1138117, 32'sd498421, -32'sd951745, -32'sd326853, 32'sd176254, 32'sd0, 32'sd0, 32'sd0, 32'sd238174, -32'sd223811, -32'sd1016920, 32'sd248151, 32'sd1573871, 32'sd998547, 32'sd2368234, -32'sd652243, 32'sd1430162, -32'sd899999, 32'sd2291636, -32'sd397759, 32'sd984171, 32'sd596265, 32'sd499509, 32'sd1686940, 32'sd919985, 32'sd1586157, 32'sd714133, 32'sd544713, 32'sd924882, -32'sd526283, -32'sd984986, 32'sd126530, 32'sd266497, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1143929, -32'sd1441626, 32'sd1619039, 32'sd1262440, -32'sd269913, -32'sd94829, 32'sd525329, 32'sd1562722, 32'sd539448, 32'sd2522940, 32'sd1040596, 32'sd894888, 32'sd2017166, 32'sd1425091, 32'sd1361814, 32'sd70424, -32'sd126696, 32'sd1691697, 32'sd350228, 32'sd152146, 32'sd451872, -32'sd824914, 32'sd293959, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd880490, 32'sd409744, -32'sd58813, 32'sd561968, 32'sd992962, -32'sd1454332, -32'sd314519, 32'sd220708, 32'sd1106557, 32'sd1681595, 32'sd1419705, 32'sd921313, 32'sd1810606, 32'sd2313328, 32'sd496601, 32'sd230509, -32'sd121262, 32'sd1432926, -32'sd1244025, 32'sd1422050, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd897749, 32'sd1153446, 32'sd758536, 32'sd275352, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd54167, -32'sd396313, -32'sd197942, -32'sd2193469, 32'sd303329, 32'sd222127, 32'sd257521, -32'sd78598, 32'sd741410, 32'sd1019600, -32'sd677048, 32'sd641974, 32'sd344802, 32'sd1002145, 32'sd762091, -32'sd372404, 32'sd140541, 32'sd450164, 32'sd1042485, 32'sd650108, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd866354, 32'sd433760, 32'sd998106, -32'sd1173223, -32'sd986899, -32'sd444558, -32'sd337719, 32'sd532808, 32'sd2459098, -32'sd765815, 32'sd1223828, -32'sd1884905, 32'sd1916214, 32'sd1326667, -32'sd1002295, 32'sd2186075, 32'sd1487902, -32'sd644831, 32'sd1426964, 32'sd1780608, 32'sd209842, 32'sd400683, -32'sd96975, 32'sd816530, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd387577, -32'sd1369370, -32'sd204716, 32'sd1599522, 32'sd560158, -32'sd829094, 32'sd3134305, -32'sd271838, -32'sd536887, 32'sd3260925, 32'sd686527, 32'sd817071, 32'sd3071279, 32'sd2815367, 32'sd451456, -32'sd2304376, -32'sd331268, 32'sd368908, 32'sd1160632, 32'sd701951, -32'sd874521, -32'sd801724, -32'sd1908445, 32'sd846540, -32'sd194672, 32'sd0, 32'sd0, 32'sd508253, 32'sd177712, -32'sd78366, -32'sd1898891, 32'sd208296, 32'sd489616, -32'sd37502, 32'sd1525333, 32'sd558761, 32'sd3299634, 32'sd2633887, -32'sd1032352, -32'sd321434, 32'sd647218, -32'sd1070077, 32'sd176414, 32'sd827119, -32'sd1113161, -32'sd577322, -32'sd1723683, -32'sd1421231, -32'sd1708704, 32'sd271967, -32'sd357748, 32'sd534806, -32'sd7251, 32'sd156572, 32'sd0, 32'sd733336, -32'sd409533, -32'sd142850, 32'sd1198756, -32'sd1002863, 32'sd1579396, 32'sd913306, 32'sd1111345, 32'sd1955643, -32'sd334164, -32'sd1513922, -32'sd486913, -32'sd887703, -32'sd1456207, -32'sd1378092, -32'sd434859, 32'sd592631, -32'sd2621692, -32'sd1458548, -32'sd1342913, -32'sd1547293, -32'sd3367620, -32'sd2060371, 32'sd152476, -32'sd230981, -32'sd2122602, 32'sd429161, 32'sd0, 32'sd930587, 32'sd614692, 32'sd1420107, 32'sd927419, -32'sd961841, 32'sd946028, -32'sd416774, -32'sd591739, 32'sd1619846, -32'sd480972, -32'sd411318, -32'sd1630662, -32'sd2030148, -32'sd2545387, -32'sd284882, 32'sd1288362, -32'sd1823300, -32'sd3389228, -32'sd2541441, -32'sd3164853, -32'sd4354480, -32'sd2384793, -32'sd3282637, -32'sd2866499, 32'sd1566927, -32'sd1185892, 32'sd1190878, 32'sd1013739, -32'sd389055, 32'sd597589, 32'sd928549, -32'sd418398, -32'sd151423, 32'sd1050109, -32'sd1218404, -32'sd825427, -32'sd1999068, -32'sd1176243, -32'sd2036592, -32'sd1354772, -32'sd982250, -32'sd2957721, 32'sd435443, 32'sd51949, -32'sd1948289, -32'sd1426729, -32'sd2306890, -32'sd2461816, -32'sd3092599, -32'sd3968727, -32'sd4555802, -32'sd1116821, -32'sd47981, -32'sd1938858, 32'sd824112, -32'sd152067, 32'sd960475, -32'sd1439945, -32'sd2699648, -32'sd1232963, 32'sd1259977, -32'sd987509, -32'sd1652832, 32'sd1236029, -32'sd1430632, -32'sd972477, -32'sd2218373, 32'sd426598, -32'sd1581644, -32'sd1571389, 32'sd989421, 32'sd2970907, -32'sd1063124, -32'sd583723, -32'sd1837956, -32'sd556231, -32'sd2106846, -32'sd2032272, -32'sd3343286, -32'sd1787574, -32'sd1370808, -32'sd475973, 32'sd1404765, -32'sd168452, 32'sd537156, -32'sd229534, -32'sd537440, 32'sd691813, -32'sd1260737, -32'sd625830, -32'sd1637726, 32'sd270727, -32'sd265912, 32'sd306380, 32'sd786536, 32'sd782333, -32'sd1117388, 32'sd516289, -32'sd253404, 32'sd1212561, 32'sd362947, -32'sd1615910, -32'sd368558, 32'sd1277323, -32'sd928327, -32'sd1436576, -32'sd553086, 32'sd274815, -32'sd649431, -32'sd13543, 32'sd413520, 32'sd731556, -32'sd287662, 32'sd804803, 32'sd2714182, 32'sd758682, 32'sd164884, -32'sd419424, -32'sd1256651, -32'sd716796, 32'sd78761, 32'sd1025133, 32'sd629433, -32'sd22177, -32'sd764348, 32'sd717391, -32'sd3432765, -32'sd1543456, -32'sd1595333, -32'sd463297, -32'sd490621, -32'sd64225, -32'sd913255, -32'sd2634563, 32'sd30725, 32'sd1219292, -32'sd2176362, 32'sd793808, -32'sd1052618, -32'sd659716, -32'sd768642, 32'sd524602, 32'sd857866, 32'sd757816, 32'sd1382257, -32'sd1132176, -32'sd1432146, 32'sd982929, 32'sd1795695, -32'sd365907, -32'sd334493, 32'sd789670, -32'sd1152151, 32'sd166170, -32'sd2242916, -32'sd2501565, -32'sd2095529, -32'sd1725332, 32'sd405597, -32'sd1231896, 32'sd1037055, 32'sd650515, 32'sd639511, -32'sd156616, 32'sd1017606, -32'sd485134, -32'sd1195281, 32'sd820742, -32'sd139600, 32'sd156566, 32'sd195397, 32'sd1124827, 32'sd66276, -32'sd2548289, -32'sd677745, 32'sd1421110, 32'sd1029352, 32'sd3207067, 32'sd966076, 32'sd555024, -32'sd32415, -32'sd1875291, -32'sd3302281, 32'sd1944336, -32'sd1447657, 32'sd416555, -32'sd2025834, 32'sd1565819, 32'sd1839253, 32'sd1374849, 32'sd1507035, -32'sd66705, 32'sd713254, -32'sd641319, 32'sd43840, -32'sd113175, -32'sd114593, 32'sd267563, -32'sd621405, 32'sd657122, 32'sd402344, -32'sd1644977, 32'sd512989, 32'sd2366169, 32'sd2188259, 32'sd1985211, 32'sd1098928, 32'sd506433, 32'sd3041763, 32'sd860178, -32'sd677300, 32'sd2973288, 32'sd1901616, 32'sd2574784, -32'sd519324, -32'sd1228858, 32'sd1564745, 32'sd2791962, 32'sd2922935, 32'sd1616234, -32'sd257475, 32'sd419527, 32'sd1417013, 32'sd347525, -32'sd112061, -32'sd46762, -32'sd1656481, 32'sd659427, 32'sd1464593, 32'sd893991, 32'sd1005959, 32'sd1278026, 32'sd2761661, 32'sd1012081, -32'sd801050, 32'sd2100912, 32'sd1941614, 32'sd1082362, 32'sd1047131, 32'sd2993065, 32'sd468341, 32'sd2037130, 32'sd786250, 32'sd598865, 32'sd516132, 32'sd1084021, 32'sd1997576, 32'sd1445417, -32'sd347572, -32'sd463547, 32'sd952980, -32'sd668278, -32'sd945602, -32'sd913721, 32'sd914775, 32'sd199198, -32'sd1481000, 32'sd1743407, 32'sd1599928, -32'sd347447, -32'sd955183, -32'sd1464268, -32'sd2510717, 32'sd1256707, 32'sd2125099, 32'sd1116840, 32'sd1011114, 32'sd3284532, 32'sd743039, 32'sd1999386, 32'sd1428163, 32'sd1171920, -32'sd530064, 32'sd123817, 32'sd219832, -32'sd145436, 32'sd659235, -32'sd774104, -32'sd1004604, 32'sd147148, 32'sd575487, 32'sd725285, 32'sd1390310, 32'sd191359, 32'sd140506, 32'sd1946856, -32'sd1137784, -32'sd1897928, 32'sd227581, 32'sd735099, 32'sd827855, 32'sd1235181, 32'sd609800, 32'sd2743236, 32'sd2461910, 32'sd634369, 32'sd1573796, 32'sd3141514, 32'sd2007571, 32'sd1361373, 32'sd1562452, 32'sd1129274, -32'sd57563, -32'sd247352, 32'sd178168, 32'sd129278, 32'sd760686, 32'sd0, -32'sd378623, -32'sd375815, 32'sd771322, -32'sd1961392, 32'sd303259, 32'sd2151263, -32'sd2112855, -32'sd402200, 32'sd31795, -32'sd1663853, 32'sd71438, -32'sd688666, 32'sd976320, 32'sd884495, 32'sd276078, 32'sd994907, 32'sd904105, 32'sd724684, 32'sd889942, 32'sd1866835, 32'sd1398595, 32'sd855051, 32'sd1228026, -32'sd1077271, 32'sd627691, -32'sd198591, 32'sd176720, 32'sd44641, -32'sd490241, -32'sd9677, 32'sd1069565, 32'sd697368, 32'sd1697857, 32'sd1429179, -32'sd396823, -32'sd436756, -32'sd178079, -32'sd11078, -32'sd627908, 32'sd706094, 32'sd23170, -32'sd1026692, 32'sd1147704, 32'sd1430937, 32'sd1712321, 32'sd545666, 32'sd2226979, 32'sd1367486, -32'sd850929, 32'sd1646827, 32'sd2521295, -32'sd1065917, 32'sd1710934, -32'sd831714, -32'sd653430, -32'sd89948, 32'sd660437, 32'sd390322, -32'sd1119222, -32'sd955725, 32'sd1273471, 32'sd862132, 32'sd296656, 32'sd175132, -32'sd1033750, 32'sd699803, -32'sd204312, -32'sd1110551, -32'sd1597700, 32'sd106061, -32'sd812077, 32'sd1344545, 32'sd1643286, -32'sd846991, 32'sd893188, -32'sd1499622, -32'sd269112, 32'sd2656654, 32'sd1059871, -32'sd2154686, 32'sd1087654, -32'sd840413, -32'sd249043, 32'sd0, -32'sd1434006, -32'sd1038793, 32'sd1654250, -32'sd1877599, 32'sd789237, 32'sd2004881, 32'sd3583782, 32'sd2651602, 32'sd639134, 32'sd1312392, 32'sd430148, -32'sd913975, -32'sd211705, 32'sd371936, -32'sd503173, -32'sd126414, -32'sd1445634, -32'sd894745, -32'sd1795580, -32'sd1957946, -32'sd1613120, -32'sd1529464, -32'sd2246031, -32'sd838361, -32'sd1177071, -32'sd251961, -32'sd263494, -32'sd640175, 32'sd132400, 32'sd518110, 32'sd2362432, -32'sd474648, -32'sd1309120, 32'sd1048856, 32'sd2183810, 32'sd984273, 32'sd2352593, 32'sd1613509, -32'sd857302, -32'sd1219590, 32'sd2574857, 32'sd1447042, -32'sd437335, -32'sd634767, 32'sd204433, -32'sd941472, -32'sd1867977, -32'sd636216, -32'sd911725, -32'sd1622973, -32'sd188235, -32'sd1561080, -32'sd212653, 32'sd752224, -32'sd306669, 32'sd813350, 32'sd469674, 32'sd320717, 32'sd346710, -32'sd3164348, 32'sd1101708, -32'sd1361461, -32'sd369753, 32'sd1532953, 32'sd1964514, 32'sd1999213, -32'sd673850, -32'sd395080, 32'sd1068305, -32'sd909506, -32'sd1465457, -32'sd2475664, -32'sd2797510, -32'sd3824297, -32'sd2090738, -32'sd3941583, -32'sd1058505, -32'sd1145954, -32'sd1458116, -32'sd815423, -32'sd778053, -32'sd1515203, 32'sd669995, 32'sd0, 32'sd68441, 32'sd1756051, 32'sd1415754, -32'sd1461302, -32'sd1607323, -32'sd2734674, -32'sd2693414, -32'sd1567668, -32'sd701888, 32'sd639234, 32'sd511852, 32'sd192069, -32'sd2320404, -32'sd853316, -32'sd1455298, -32'sd3858418, -32'sd4189961, -32'sd5158896, -32'sd3803407, -32'sd1663972, -32'sd2460857, -32'sd2173901, -32'sd1937653, 32'sd330427, -32'sd436278, -32'sd1034325, 32'sd0, 32'sd0, 32'sd0, 32'sd852558, 32'sd903406, -32'sd1337104, -32'sd1783333, -32'sd1318798, -32'sd2818977, -32'sd3376809, -32'sd309164, 32'sd237946, 32'sd399469, -32'sd3359032, -32'sd2555001, -32'sd1382948, -32'sd2946112, -32'sd2039834, 32'sd227351, -32'sd2592937, -32'sd2253521, -32'sd762900, -32'sd369598, 32'sd52019, -32'sd742812, -32'sd321305, -32'sd861006, 32'sd837909, 32'sd0, 32'sd0, 32'sd0, -32'sd790585, 32'sd96482, -32'sd588348, 32'sd333725, -32'sd238953, -32'sd1351068, -32'sd2867412, -32'sd1129082, -32'sd1688115, -32'sd2177239, -32'sd1895406, -32'sd1475496, -32'sd933682, 32'sd228179, -32'sd655219, 32'sd387237, -32'sd1427205, 32'sd909546, 32'sd708309, -32'sd189283, -32'sd886406, -32'sd1913395, -32'sd1744160, 32'sd18572, 32'sd223462, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd653485, 32'sd616524, -32'sd450384, -32'sd13782, 32'sd883364, -32'sd364636, -32'sd2319061, -32'sd1084649, -32'sd1090497, -32'sd128094, -32'sd1934221, 32'sd1125087, 32'sd1524254, -32'sd2178284, -32'sd2515942, 32'sd1260980, -32'sd130486, 32'sd406827, -32'sd696763, -32'sd932921, -32'sd1441077, 32'sd200812, 32'sd197777, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd531087, -32'sd199558, 32'sd850056, 32'sd223936, -32'sd294179, 32'sd1347834, 32'sd446919, -32'sd985474, 32'sd1901688, -32'sd1279896, -32'sd1063289, 32'sd614192, 32'sd745276, -32'sd481966, -32'sd2912, 32'sd509255, -32'sd760978, -32'sd582847, 32'sd456798, 32'sd44722, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1866340, 32'sd2169257, 32'sd1327336, 32'sd1047303, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2202038, 32'sd1289689, 32'sd101323, -32'sd197674, 32'sd1504037, -32'sd902240, 32'sd1340553, -32'sd181046, -32'sd21267, -32'sd23474, -32'sd51518, 32'sd1383398, 32'sd218613, 32'sd1772971, 32'sd1362287, 32'sd745747, 32'sd635035, -32'sd88065, -32'sd134372, 32'sd282031, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd112097, -32'sd240135, 32'sd1373599, -32'sd949310, -32'sd191552, -32'sd494006, 32'sd1421080, 32'sd1284792, 32'sd1190874, 32'sd682507, -32'sd610346, -32'sd2000227, 32'sd1699714, 32'sd1331587, 32'sd453543, -32'sd2003832, -32'sd623177, -32'sd366156, 32'sd649154, -32'sd39712, 32'sd1356535, -32'sd17852, 32'sd572915, 32'sd311303, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd494186, 32'sd282885, -32'sd46452, -32'sd201728, -32'sd2440988, -32'sd1959625, 32'sd2434801, 32'sd855468, -32'sd1541743, -32'sd353478, -32'sd508683, -32'sd71553, -32'sd1837019, -32'sd2408610, -32'sd1216527, -32'sd1350302, -32'sd307259, 32'sd913013, -32'sd1873426, 32'sd653753, 32'sd1219921, 32'sd688850, 32'sd977317, 32'sd292037, 32'sd1509198, 32'sd0, 32'sd0, 32'sd642595, 32'sd1455658, 32'sd736548, -32'sd416111, -32'sd1405656, 32'sd878827, 32'sd226468, 32'sd1380199, 32'sd294160, 32'sd2016254, -32'sd1366354, 32'sd1059770, -32'sd1668427, -32'sd2953138, -32'sd2700207, -32'sd3085907, -32'sd3387751, -32'sd3521639, -32'sd1521305, -32'sd1097076, 32'sd203422, -32'sd737185, 32'sd50600, 32'sd230786, 32'sd559845, 32'sd691669, -32'sd274218, 32'sd0, 32'sd194013, -32'sd414989, -32'sd870689, 32'sd255329, -32'sd1375802, 32'sd1295516, 32'sd1353489, -32'sd1359498, -32'sd726801, -32'sd2655799, -32'sd1924220, -32'sd3064785, -32'sd1886909, -32'sd1228764, -32'sd987976, -32'sd1199099, -32'sd2378558, 32'sd55223, 32'sd488198, -32'sd2208091, -32'sd1398391, -32'sd239146, -32'sd1966743, 32'sd1283522, 32'sd2148487, 32'sd841581, 32'sd1321154, 32'sd0, 32'sd1823128, 32'sd250799, 32'sd1145732, -32'sd296209, -32'sd1768016, -32'sd357288, -32'sd79205, -32'sd686649, 32'sd533225, -32'sd34196, -32'sd779462, -32'sd839476, -32'sd792196, 32'sd353462, -32'sd137200, 32'sd529848, -32'sd139255, -32'sd2025442, 32'sd1122417, -32'sd2018320, -32'sd3000894, -32'sd3267872, -32'sd645598, -32'sd2139874, 32'sd1542437, 32'sd1451619, -32'sd415937, 32'sd826083, 32'sd1090558, -32'sd722757, -32'sd806698, -32'sd1866163, -32'sd285808, -32'sd144196, -32'sd915067, -32'sd1392037, 32'sd1201498, 32'sd514907, 32'sd356015, 32'sd503444, 32'sd1897655, 32'sd426190, -32'sd2764959, -32'sd4047621, -32'sd2830739, -32'sd3255527, -32'sd2556807, -32'sd838923, 32'sd443339, -32'sd1464428, -32'sd1527741, -32'sd781724, 32'sd1725128, 32'sd1154919, 32'sd711831, 32'sd842175, 32'sd1667492, -32'sd465923, -32'sd735483, -32'sd1141110, -32'sd957501, -32'sd776807, -32'sd1889737, 32'sd926588, 32'sd1890619, 32'sd3542642, 32'sd2411015, 32'sd1860485, 32'sd3227999, -32'sd24727, -32'sd728299, -32'sd2264504, -32'sd2849225, -32'sd1288184, 32'sd1098196, -32'sd592549, 32'sd98253, -32'sd777221, 32'sd141099, -32'sd1925810, -32'sd345427, 32'sd62703, 32'sd63492, 32'sd2030045, 32'sd1333389, 32'sd2082120, 32'sd251732, 32'sd494254, -32'sd1233373, 32'sd1192405, -32'sd517333, 32'sd467875, 32'sd290640, 32'sd2715930, 32'sd426013, 32'sd1100225, 32'sd1253329, 32'sd1641982, -32'sd217946, -32'sd2127997, -32'sd91740, -32'sd974713, 32'sd2305875, 32'sd2218669, 32'sd2947460, 32'sd1469279, 32'sd269419, 32'sd847817, -32'sd322698, 32'sd1292065, 32'sd1282373, 32'sd30118, -32'sd970885, -32'sd328725, 32'sd569040, 32'sd1553993, 32'sd891865, 32'sd500897, 32'sd447681, 32'sd1862002, 32'sd2849997, 32'sd878868, 32'sd946847, -32'sd773643, -32'sd994302, -32'sd2305695, -32'sd2193946, -32'sd419094, -32'sd797344, 32'sd423384, 32'sd2272572, 32'sd2210867, 32'sd1262729, 32'sd1394175, 32'sd1240306, -32'sd929445, -32'sd563774, 32'sd1040277, 32'sd1288009, 32'sd908608, 32'sd592881, 32'sd1032064, 32'sd803326, 32'sd1127251, 32'sd1933550, 32'sd478582, -32'sd228741, 32'sd1485731, 32'sd1330562, -32'sd688150, -32'sd1575593, -32'sd4880506, -32'sd3251079, -32'sd1043835, -32'sd1447534, -32'sd994388, -32'sd829493, -32'sd2090159, 32'sd1564879, 32'sd1654246, 32'sd1669461, 32'sd2420652, 32'sd1477238, -32'sd1565960, 32'sd536641, 32'sd1569063, 32'sd950572, 32'sd66936, 32'sd688105, 32'sd51191, 32'sd515090, 32'sd1638464, 32'sd1411691, -32'sd1158754, -32'sd184998, 32'sd88721, 32'sd32882, -32'sd1908755, -32'sd4733454, -32'sd3226756, -32'sd2086435, -32'sd53208, 32'sd3046452, 32'sd2906428, -32'sd542502, -32'sd1393408, -32'sd1080519, -32'sd913586, 32'sd123038, 32'sd2205902, 32'sd1427954, 32'sd551297, 32'sd477077, 32'sd378152, 32'sd275882, -32'sd99916, -32'sd1158297, -32'sd1057520, 32'sd657257, 32'sd478940, 32'sd862695, -32'sd1358650, -32'sd483396, -32'sd1939223, -32'sd4560208, -32'sd4308289, -32'sd2356327, -32'sd1086187, -32'sd144032, -32'sd161904, 32'sd412865, 32'sd2884976, -32'sd79797, 32'sd1040713, 32'sd130987, 32'sd611517, 32'sd1456682, 32'sd802143, 32'sd84415, 32'sd2483099, 32'sd129532, 32'sd83133, 32'sd171808, -32'sd1329099, 32'sd405281, -32'sd89488, -32'sd75308, -32'sd562043, -32'sd98241, 32'sd1222501, -32'sd984122, -32'sd726970, -32'sd4268004, -32'sd1996742, -32'sd1287793, 32'sd1677346, 32'sd2578253, -32'sd441138, 32'sd157108, -32'sd1935165, 32'sd239070, 32'sd1312657, 32'sd1605297, -32'sd615477, 32'sd825977, -32'sd124838, -32'sd1666447, -32'sd458772, -32'sd827402, 32'sd1761062, -32'sd775972, 32'sd478221, 32'sd1041944, -32'sd1185753, 32'sd206769, -32'sd1417251, 32'sd723752, 32'sd508727, -32'sd1685321, -32'sd3223181, -32'sd1471694, -32'sd1161781, 32'sd1119075, 32'sd615362, 32'sd1952134, 32'sd2696650, 32'sd2138934, 32'sd869029, 32'sd475156, 32'sd681464, 32'sd1910850, 32'sd2156513, 32'sd83387, 32'sd427697, 32'sd420251, -32'sd1329271, -32'sd403862, 32'sd1531910, 32'sd935815, 32'sd113910, -32'sd261341, 32'sd404831, 32'sd539018, -32'sd837684, -32'sd535099, 32'sd1225485, -32'sd67297, -32'sd1279711, -32'sd230390, 32'sd49916, -32'sd1051184, 32'sd1058723, 32'sd2971927, 32'sd4028280, 32'sd1607003, 32'sd1052055, 32'sd646359, 32'sd2906561, 32'sd3245826, 32'sd1386922, -32'sd432123, -32'sd468117, -32'sd1833632, 32'sd98723, 32'sd441007, 32'sd1437324, -32'sd1722880, 32'sd0, 32'sd341748, -32'sd1875619, 32'sd1268637, 32'sd320631, -32'sd457651, 32'sd51392, -32'sd1456309, -32'sd230988, 32'sd1394759, -32'sd501295, 32'sd606781, 32'sd2544294, 32'sd2802539, 32'sd2224703, -32'sd4318, -32'sd387433, 32'sd169043, 32'sd2294790, 32'sd1592743, 32'sd612042, -32'sd2120813, -32'sd1045519, -32'sd2308208, -32'sd2348876, -32'sd1740939, -32'sd1114112, -32'sd351615, 32'sd1075708, -32'sd1064110, 32'sd360326, 32'sd669398, -32'sd649176, 32'sd231628, 32'sd254773, 32'sd3404156, 32'sd729118, -32'sd594550, 32'sd620504, 32'sd1400196, -32'sd625264, 32'sd1522279, 32'sd1839030, -32'sd710728, 32'sd305336, 32'sd3599940, 32'sd1684435, 32'sd3272715, 32'sd81819, -32'sd1052778, -32'sd652395, -32'sd1173112, -32'sd874112, -32'sd1850627, -32'sd627335, 32'sd1447199, 32'sd57414, 32'sd979492, -32'sd2273118, -32'sd1324347, 32'sd3176602, 32'sd2309845, 32'sd850483, 32'sd2284770, 32'sd2313960, -32'sd902295, -32'sd700051, 32'sd772823, -32'sd1051271, -32'sd2396583, -32'sd359691, 32'sd583921, 32'sd2886419, 32'sd253360, 32'sd29968, 32'sd1064649, -32'sd1743225, 32'sd702886, 32'sd702928, -32'sd326275, -32'sd783989, -32'sd3912206, 32'sd1646405, -32'sd260915, 32'sd0, -32'sd257715, -32'sd852644, 32'sd717239, 32'sd3035380, 32'sd1691939, 32'sd373521, 32'sd1242719, 32'sd1084732, -32'sd226232, 32'sd1011897, -32'sd2302450, -32'sd2751828, -32'sd2639052, 32'sd99574, 32'sd263740, 32'sd848008, -32'sd2476246, 32'sd20322, -32'sd416026, -32'sd1044268, -32'sd1694300, -32'sd1315045, -32'sd1006516, -32'sd104634, -32'sd2601018, 32'sd1542144, 32'sd658852, -32'sd540327, 32'sd66881, 32'sd276495, 32'sd2679054, 32'sd375592, 32'sd1455257, 32'sd112772, 32'sd1008081, 32'sd359643, -32'sd2110913, 32'sd205770, -32'sd2116994, -32'sd1547820, -32'sd2545195, 32'sd340951, -32'sd2230695, -32'sd317613, -32'sd1152507, 32'sd313987, -32'sd1800823, -32'sd2826778, -32'sd1510714, -32'sd1069713, 32'sd603216, 32'sd560632, -32'sd113407, 32'sd929109, 32'sd1366372, -32'sd431352, -32'sd81326, 32'sd1066488, 32'sd300811, 32'sd111510, -32'sd690327, -32'sd2449883, -32'sd2056093, -32'sd586868, -32'sd2038733, -32'sd888779, -32'sd2602972, -32'sd591795, -32'sd2493718, -32'sd2612585, 32'sd274760, 32'sd565238, 32'sd333134, 32'sd659499, 32'sd328202, -32'sd1007785, -32'sd1747044, -32'sd1792999, 32'sd797237, 32'sd178759, -32'sd108436, -32'sd1506827, 32'sd164049, 32'sd0, -32'sd5558, 32'sd361321, -32'sd448719, -32'sd708449, -32'sd725931, -32'sd435474, -32'sd2101497, -32'sd1737783, -32'sd506874, -32'sd1040970, -32'sd57937, -32'sd165193, -32'sd89091, -32'sd329148, -32'sd276534, 32'sd83063, -32'sd12792, 32'sd843265, -32'sd152107, -32'sd342599, -32'sd1343561, -32'sd906843, 32'sd918366, 32'sd1704829, -32'sd250999, -32'sd1399622, 32'sd0, 32'sd0, 32'sd0, 32'sd1424268, -32'sd339217, 32'sd744337, -32'sd400451, -32'sd971469, -32'sd1148226, -32'sd208667, 32'sd235205, -32'sd133735, 32'sd241485, 32'sd5429, -32'sd1272055, -32'sd16332, -32'sd1025966, -32'sd1316689, 32'sd765218, -32'sd1190956, -32'sd384492, 32'sd2003737, 32'sd1108120, -32'sd602579, -32'sd880707, 32'sd1254267, -32'sd924172, 32'sd915322, 32'sd0, 32'sd0, 32'sd0, -32'sd677725, 32'sd297065, -32'sd902440, -32'sd216306, -32'sd2079179, -32'sd276702, -32'sd755429, 32'sd1983041, -32'sd148700, -32'sd2073231, 32'sd277095, -32'sd783579, -32'sd1311493, -32'sd1832851, 32'sd1503458, -32'sd412307, -32'sd676243, 32'sd1547991, 32'sd336927, -32'sd531321, -32'sd371063, -32'sd239954, -32'sd846265, -32'sd723334, 32'sd762711, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd6269, -32'sd1299332, -32'sd203586, 32'sd288152, 32'sd1126586, 32'sd693690, 32'sd603381, -32'sd801442, -32'sd189898, 32'sd301071, 32'sd39980, 32'sd658717, -32'sd1607730, 32'sd349703, -32'sd208982, -32'sd782538, 32'sd903111, 32'sd1547390, 32'sd1132592, 32'sd45587, -32'sd985241, -32'sd147000, -32'sd34292, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd307606, -32'sd237298, -32'sd9017, 32'sd2052446, 32'sd115893, 32'sd848193, 32'sd488026, 32'sd838206, 32'sd866743, -32'sd149901, 32'sd1879680, 32'sd441200, 32'sd1230808, -32'sd101963, 32'sd361525, 32'sd2222868, 32'sd349472, 32'sd591271, -32'sd1013249, 32'sd359014, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd907446, 32'sd466535, 32'sd1369565, 32'sd2182902, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd636112, 32'sd629422, -32'sd66326, 32'sd1118508, -32'sd1534157, 32'sd233924, 32'sd891294, 32'sd414806, 32'sd162497, -32'sd591241, 32'sd1124654, 32'sd1157149, -32'sd229680, 32'sd335665, 32'sd58784, -32'sd714209, 32'sd584212, 32'sd528556, 32'sd830242, 32'sd1206458, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1245288, 32'sd188860, -32'sd425895, -32'sd143504, -32'sd184317, -32'sd889513, -32'sd1093599, -32'sd969414, -32'sd1635217, 32'sd823430, 32'sd431039, 32'sd2782906, 32'sd403127, 32'sd2127472, 32'sd998563, 32'sd736061, 32'sd1144309, 32'sd2001067, 32'sd1627644, 32'sd606698, -32'sd356183, 32'sd403799, 32'sd1333316, 32'sd1642593, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1581934, -32'sd427621, 32'sd936346, 32'sd1704277, 32'sd76205, 32'sd362649, 32'sd1696711, 32'sd1901209, 32'sd2393810, 32'sd42364, -32'sd546479, 32'sd503477, 32'sd695559, -32'sd652043, 32'sd2518210, 32'sd105497, 32'sd1480549, -32'sd1197483, 32'sd305933, 32'sd844189, -32'sd408785, -32'sd906242, 32'sd1034157, -32'sd5501, -32'sd304377, 32'sd0, 32'sd0, 32'sd758960, 32'sd992461, 32'sd1588314, 32'sd263581, 32'sd596613, 32'sd1778184, 32'sd1764431, -32'sd141899, 32'sd2000706, 32'sd19720, 32'sd1678317, 32'sd2323641, 32'sd972834, -32'sd265460, -32'sd78270, -32'sd193765, -32'sd1501396, 32'sd50931, -32'sd924714, -32'sd1180130, -32'sd648829, 32'sd1419850, 32'sd2074932, 32'sd1380849, -32'sd519888, 32'sd1084388, 32'sd1340964, 32'sd0, 32'sd1848122, 32'sd259621, 32'sd1584059, -32'sd1666106, 32'sd315920, -32'sd1310709, 32'sd1304502, -32'sd1041170, -32'sd1169293, 32'sd420404, -32'sd539018, 32'sd983379, -32'sd1998919, -32'sd640949, -32'sd488599, -32'sd576895, -32'sd1765882, 32'sd1792889, -32'sd146746, -32'sd1855040, 32'sd484879, -32'sd573910, -32'sd114267, -32'sd154572, 32'sd34344, 32'sd1305764, -32'sd311040, 32'sd0, 32'sd1088754, 32'sd64099, 32'sd138877, -32'sd1003871, -32'sd187971, -32'sd1824822, -32'sd1868475, -32'sd60751, -32'sd712237, -32'sd952619, -32'sd113468, 32'sd962290, -32'sd925404, -32'sd93009, 32'sd771478, -32'sd788119, 32'sd450538, -32'sd687102, -32'sd961420, -32'sd2142940, 32'sd407636, -32'sd1088157, -32'sd1510285, 32'sd862105, -32'sd120179, 32'sd932858, -32'sd345465, 32'sd1431765, -32'sd980814, -32'sd397594, 32'sd408083, -32'sd857269, -32'sd1340428, 32'sd266487, -32'sd62053, -32'sd559179, -32'sd316581, 32'sd336325, 32'sd614217, 32'sd62433, 32'sd3040704, 32'sd1240133, 32'sd2083712, 32'sd871801, -32'sd184872, 32'sd701847, -32'sd739440, -32'sd676371, -32'sd2478819, -32'sd2690342, 32'sd62528, 32'sd108861, -32'sd1667248, 32'sd590555, -32'sd19371, 32'sd1361686, 32'sd205251, -32'sd514035, 32'sd305190, -32'sd1803472, -32'sd1325081, -32'sd704929, -32'sd91550, 32'sd613299, 32'sd51220, -32'sd128489, 32'sd353712, 32'sd2282699, 32'sd2648462, 32'sd2422295, 32'sd2605076, 32'sd310230, 32'sd2061964, 32'sd1962275, 32'sd2034304, -32'sd119100, -32'sd289448, 32'sd201931, -32'sd155642, -32'sd642035, 32'sd425921, -32'sd1270730, 32'sd824220, 32'sd45990, 32'sd1140676, 32'sd957778, -32'sd591743, -32'sd2026410, -32'sd1977981, 32'sd1400413, 32'sd136241, -32'sd496327, 32'sd569498, 32'sd110900, 32'sd337870, 32'sd1045593, 32'sd1883885, 32'sd1506821, 32'sd1345253, 32'sd1124940, 32'sd1810574, 32'sd2092369, 32'sd1866562, 32'sd1357821, -32'sd3011073, -32'sd1676013, -32'sd951938, 32'sd534748, 32'sd860960, 32'sd705813, 32'sd102306, 32'sd1332775, -32'sd477356, 32'sd335625, -32'sd1126193, -32'sd2308259, -32'sd378830, 32'sd554921, 32'sd775086, 32'sd1593161, 32'sd952629, 32'sd484052, -32'sd6320, -32'sd202005, 32'sd2305897, 32'sd2543278, 32'sd4875928, 32'sd2496739, 32'sd2182213, 32'sd778753, 32'sd2042476, 32'sd2847699, -32'sd2016144, 32'sd1600459, 32'sd1304358, -32'sd1465825, 32'sd1274091, -32'sd1689916, 32'sd607920, 32'sd1360462, 32'sd1991461, 32'sd345253, 32'sd2685125, 32'sd524018, -32'sd816272, 32'sd1839633, 32'sd651777, 32'sd803933, 32'sd446004, 32'sd372259, 32'sd299643, 32'sd561708, -32'sd1058452, 32'sd807374, 32'sd2443564, -32'sd514450, 32'sd1105249, 32'sd3241571, 32'sd448596, 32'sd3648053, 32'sd592437, 32'sd1357880, -32'sd342797, -32'sd1351376, 32'sd1525755, 32'sd724986, 32'sd398346, 32'sd670961, 32'sd132049, 32'sd511045, 32'sd1261139, 32'sd921092, 32'sd112624, 32'sd178918, -32'sd1301753, -32'sd970754, 32'sd718110, -32'sd1737741, -32'sd1934453, -32'sd1951007, -32'sd1671790, 32'sd373401, 32'sd225118, 32'sd2036511, 32'sd277217, 32'sd2999177, 32'sd1772227, 32'sd2651387, 32'sd71029, -32'sd865897, -32'sd752177, 32'sd111736, -32'sd163443, -32'sd292941, -32'sd796990, 32'sd875923, -32'sd725211, 32'sd174390, 32'sd936479, 32'sd948463, -32'sd1575763, 32'sd944332, -32'sd1346228, 32'sd674468, -32'sd707635, -32'sd2937379, -32'sd1714678, -32'sd2036781, -32'sd2160738, -32'sd77350, 32'sd667665, 32'sd191443, 32'sd959978, 32'sd1650412, 32'sd1891091, 32'sd2445418, 32'sd979636, -32'sd1071771, -32'sd2424635, -32'sd1675503, -32'sd736081, -32'sd11781, -32'sd56124, 32'sd515845, 32'sd1507730, 32'sd1123658, -32'sd105921, -32'sd608142, 32'sd6692, 32'sd1231627, -32'sd1017165, 32'sd505200, -32'sd421807, -32'sd1459201, -32'sd2131350, -32'sd2492239, -32'sd3371832, -32'sd1634065, -32'sd535619, 32'sd805607, -32'sd231957, 32'sd2120416, -32'sd24840, 32'sd2031010, 32'sd642444, -32'sd811860, -32'sd175002, -32'sd691993, 32'sd480644, 32'sd1106588, -32'sd930408, 32'sd398171, -32'sd22852, -32'sd1751423, -32'sd1598165, 32'sd569529, -32'sd441598, -32'sd506220, -32'sd1823052, -32'sd935178, -32'sd781422, -32'sd2450237, -32'sd2460401, -32'sd2267207, -32'sd742688, -32'sd1486669, -32'sd1358918, -32'sd1201159, -32'sd316027, -32'sd502356, 32'sd473285, 32'sd1717271, 32'sd1739077, 32'sd61465, 32'sd1973917, 32'sd895897, 32'sd356088, -32'sd871669, 32'sd816824, 32'sd876619, 32'sd627331, -32'sd1725087, 32'sd347853, 32'sd1194651, 32'sd1624491, -32'sd873766, -32'sd685765, -32'sd849608, -32'sd940787, -32'sd1180780, -32'sd1127564, 32'sd97368, -32'sd2007894, -32'sd615575, -32'sd1212654, 32'sd475519, 32'sd771780, -32'sd213345, -32'sd1342817, -32'sd417766, -32'sd240927, -32'sd1438485, -32'sd237316, 32'sd2009981, -32'sd874752, -32'sd1137096, 32'sd341626, 32'sd0, -32'sd588089, -32'sd422035, 32'sd746431, 32'sd1120447, 32'sd240091, -32'sd341278, -32'sd847919, -32'sd720730, -32'sd662776, 32'sd200183, -32'sd903342, -32'sd110827, -32'sd471422, -32'sd1074306, -32'sd1782887, -32'sd1756745, 32'sd411490, 32'sd2060816, 32'sd1089560, 32'sd92157, 32'sd961383, 32'sd361524, -32'sd1705365, 32'sd486822, 32'sd365369, -32'sd303999, 32'sd284104, -32'sd181040, 32'sd360975, 32'sd60568, 32'sd903325, -32'sd97805, -32'sd144317, 32'sd907848, -32'sd959432, -32'sd1170163, -32'sd2130874, 32'sd882851, -32'sd350940, -32'sd271896, -32'sd749537, -32'sd1770458, -32'sd2007823, -32'sd1636575, 32'sd2098207, 32'sd1266412, 32'sd532609, 32'sd899681, 32'sd824945, 32'sd1289259, -32'sd1902398, -32'sd942189, 32'sd134997, -32'sd946537, 32'sd1528934, 32'sd859782, -32'sd1194444, -32'sd340866, -32'sd122208, 32'sd370479, 32'sd417199, -32'sd1970916, -32'sd202044, -32'sd1514052, -32'sd609983, -32'sd486076, -32'sd958895, 32'sd283857, -32'sd2149230, -32'sd473413, 32'sd44703, -32'sd884604, 32'sd638541, 32'sd2020655, 32'sd2879057, 32'sd2413140, 32'sd109217, -32'sd318720, -32'sd3756193, 32'sd268992, 32'sd160108, -32'sd1303522, 32'sd763817, 32'sd0, 32'sd755531, 32'sd94282, -32'sd1872244, 32'sd95464, -32'sd54222, -32'sd1265467, -32'sd1045411, -32'sd104022, -32'sd1242292, -32'sd1896841, -32'sd197901, -32'sd1590439, -32'sd416235, 32'sd240283, 32'sd385749, 32'sd1035445, 32'sd2005780, 32'sd236102, 32'sd690214, -32'sd323637, -32'sd2114070, -32'sd1353865, -32'sd1348195, -32'sd1916738, 32'sd1283293, 32'sd1442038, 32'sd998175, 32'sd1417115, 32'sd337902, -32'sd303812, 32'sd267688, -32'sd809441, 32'sd362719, -32'sd699681, 32'sd727351, -32'sd1711514, 32'sd402664, -32'sd1193068, -32'sd545234, 32'sd292029, 32'sd900845, -32'sd420007, -32'sd69312, 32'sd1241816, 32'sd356753, 32'sd621062, -32'sd703701, 32'sd664937, -32'sd1461528, -32'sd947661, -32'sd311422, -32'sd1193003, 32'sd1615525, 32'sd445612, 32'sd1397070, 32'sd1965614, -32'sd333759, 32'sd1426910, 32'sd244213, 32'sd1375518, 32'sd1599724, 32'sd803803, 32'sd26964, -32'sd249873, 32'sd435226, -32'sd292356, 32'sd2434321, 32'sd1545766, 32'sd1474093, 32'sd2079118, -32'sd252058, -32'sd193944, 32'sd176685, -32'sd555716, 32'sd1477248, -32'sd1374055, -32'sd1826499, -32'sd1412224, -32'sd645974, -32'sd265711, 32'sd445615, -32'sd196148, 32'sd511597, 32'sd0, 32'sd1255164, -32'sd146155, -32'sd483642, -32'sd988462, 32'sd159341, 32'sd1701392, 32'sd254875, -32'sd302623, -32'sd1732143, -32'sd441031, 32'sd1096812, -32'sd10013, 32'sd341004, 32'sd1284944, 32'sd1927148, 32'sd498236, 32'sd534274, 32'sd1126628, 32'sd897372, -32'sd448150, -32'sd616800, -32'sd1049371, 32'sd1247486, 32'sd645547, -32'sd278288, 32'sd1117232, 32'sd0, 32'sd0, 32'sd0, -32'sd505862, 32'sd1557931, -32'sd352927, -32'sd433439, 32'sd561107, 32'sd179128, 32'sd748912, 32'sd2179661, 32'sd828244, 32'sd165182, 32'sd331883, 32'sd112700, 32'sd608505, -32'sd1130543, -32'sd874344, -32'sd434211, 32'sd334347, -32'sd1320402, -32'sd1446243, -32'sd83929, 32'sd1253578, 32'sd1648240, 32'sd6235, 32'sd488310, -32'sd309588, 32'sd0, 32'sd0, 32'sd0, 32'sd1340548, 32'sd1683395, 32'sd774021, 32'sd319426, -32'sd299127, 32'sd1144039, 32'sd2497577, 32'sd1955665, 32'sd393678, 32'sd1392424, 32'sd1178825, -32'sd1030801, 32'sd2966699, -32'sd915159, 32'sd102113, -32'sd286460, 32'sd839855, -32'sd492900, -32'sd1185830, -32'sd441577, 32'sd1563934, -32'sd903240, 32'sd1347030, 32'sd546807, -32'sd91674, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1948832, 32'sd909423, -32'sd1426923, -32'sd1513502, 32'sd346774, -32'sd68301, 32'sd2112539, 32'sd3011082, 32'sd817600, 32'sd393437, 32'sd609276, 32'sd792288, 32'sd1487635, 32'sd1649476, 32'sd635205, 32'sd1685684, 32'sd2090986, -32'sd622613, -32'sd1302372, 32'sd1106491, -32'sd446766, 32'sd451600, 32'sd991807, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2338521, 32'sd1139119, 32'sd974675, 32'sd1231614, 32'sd922344, -32'sd795383, 32'sd2073170, 32'sd425721, 32'sd1033791, -32'sd118890, 32'sd1197838, 32'sd1903395, 32'sd798928, 32'sd705201, -32'sd507287, 32'sd1171001, 32'sd1390869, 32'sd194626, 32'sd567159, 32'sd1343512, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1683596, 32'sd376109, -32'sd414789, 32'sd157249, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd219869, 32'sd250312, -32'sd875619, 32'sd360025, -32'sd957075, -32'sd727933, -32'sd163679, -32'sd27718, 32'sd1349244, -32'sd1975560, -32'sd2076278, -32'sd1859837, -32'sd1419242, -32'sd1700176, 32'sd257558, -32'sd1541581, -32'sd14008, -32'sd1506154, -32'sd1173443, -32'sd1013636, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd989174, -32'sd1124799, -32'sd1628426, -32'sd1591350, 32'sd709016, -32'sd918138, 32'sd928712, 32'sd334031, 32'sd1410903, -32'sd796623, 32'sd1167828, 32'sd1957246, 32'sd801919, 32'sd221079, 32'sd582464, -32'sd1279420, -32'sd1702423, -32'sd335366, -32'sd991743, -32'sd570408, 32'sd391424, -32'sd995759, -32'sd459536, 32'sd389049, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd869821, 32'sd464022, -32'sd1197581, -32'sd2294940, 32'sd548176, -32'sd663023, 32'sd934868, -32'sd600372, 32'sd1925290, 32'sd379626, 32'sd611681, 32'sd1894591, -32'sd859464, 32'sd2151054, 32'sd2876775, 32'sd1930939, -32'sd62023, 32'sd706614, -32'sd12384, 32'sd690021, -32'sd1651897, -32'sd316350, -32'sd1318221, -32'sd1771731, -32'sd1324170, 32'sd0, 32'sd0, 32'sd431865, -32'sd1205967, -32'sd1485586, -32'sd1324765, 32'sd405855, 32'sd1726436, 32'sd237216, 32'sd975381, 32'sd2801525, -32'sd300512, 32'sd808345, 32'sd2601404, -32'sd506691, 32'sd907399, -32'sd338998, 32'sd2437783, 32'sd2712616, 32'sd1476705, -32'sd327930, 32'sd479249, -32'sd120631, 32'sd345205, -32'sd543789, -32'sd530889, 32'sd361074, -32'sd287088, 32'sd821852, 32'sd0, 32'sd433360, -32'sd1308741, -32'sd907909, -32'sd778215, 32'sd1636127, -32'sd537876, 32'sd2307202, -32'sd756498, 32'sd1184991, -32'sd699746, 32'sd1489376, 32'sd2376474, 32'sd2184772, 32'sd1837260, 32'sd434587, 32'sd393342, 32'sd926612, -32'sd261589, -32'sd697473, 32'sd1017605, 32'sd2976650, -32'sd768201, -32'sd780069, -32'sd3173961, -32'sd526450, 32'sd174605, 32'sd1067117, 32'sd0, -32'sd820264, -32'sd568266, -32'sd484804, 32'sd742318, 32'sd1310347, 32'sd847140, 32'sd1902659, 32'sd982334, 32'sd95115, 32'sd445888, 32'sd690490, 32'sd1817620, 32'sd264949, 32'sd1672617, -32'sd462827, 32'sd1256581, -32'sd354737, 32'sd1094074, 32'sd992080, 32'sd1381577, 32'sd2518950, 32'sd872977, -32'sd91612, 32'sd574213, -32'sd387359, -32'sd633349, 32'sd445765, -32'sd41350, -32'sd1295136, 32'sd161781, -32'sd734520, -32'sd212270, -32'sd1307308, 32'sd521617, -32'sd941158, 32'sd1194, 32'sd1705073, 32'sd1123155, 32'sd2194289, 32'sd2044366, 32'sd1842701, 32'sd1872748, 32'sd636747, -32'sd1616169, -32'sd497293, 32'sd1237536, 32'sd2470303, 32'sd425991, -32'sd88279, 32'sd1647797, 32'sd1000402, 32'sd354930, 32'sd799805, -32'sd1397724, -32'sd1007396, -32'sd516819, 32'sd829644, 32'sd701889, -32'sd658848, -32'sd899383, -32'sd700811, 32'sd1077248, 32'sd1020174, -32'sd551772, 32'sd693717, 32'sd1966823, 32'sd3449685, 32'sd2666989, 32'sd1819622, -32'sd592103, -32'sd804990, -32'sd1044852, 32'sd469400, 32'sd629261, 32'sd207109, -32'sd869593, -32'sd732598, 32'sd1604237, 32'sd2348516, 32'sd970395, 32'sd224939, 32'sd869660, -32'sd671958, 32'sd1609557, 32'sd1878795, -32'sd685065, -32'sd2220719, -32'sd749981, -32'sd1629804, -32'sd799118, -32'sd1870454, -32'sd1119676, -32'sd541281, 32'sd1470921, 32'sd2457510, 32'sd2847011, 32'sd2404045, 32'sd1600549, 32'sd1184536, -32'sd2206420, 32'sd716852, 32'sd684048, 32'sd997711, -32'sd662232, 32'sd39802, -32'sd595855, 32'sd644415, -32'sd259918, 32'sd555192, 32'sd81296, -32'sd1138799, -32'sd141912, 32'sd904474, -32'sd207041, -32'sd1213761, -32'sd1132165, -32'sd1267654, -32'sd2902918, -32'sd1847538, -32'sd3142645, -32'sd2440179, -32'sd376873, 32'sd836766, 32'sd2728462, 32'sd2766900, 32'sd1255202, 32'sd674230, -32'sd866768, 32'sd678068, 32'sd1944559, -32'sd1258800, -32'sd635875, -32'sd2234021, -32'sd2808190, -32'sd460565, -32'sd2185228, -32'sd1144391, 32'sd885487, -32'sd255989, 32'sd422501, 32'sd1503307, 32'sd1655526, 32'sd568789, 32'sd778012, -32'sd1479764, -32'sd1719038, -32'sd3672997, -32'sd2734708, -32'sd3136146, -32'sd1984021, -32'sd471279, 32'sd2762631, 32'sd499671, 32'sd1537801, 32'sd3571331, 32'sd1380583, 32'sd1604700, -32'sd431165, -32'sd1190850, -32'sd1711465, -32'sd2133255, -32'sd953431, -32'sd667172, -32'sd2060566, -32'sd43502, 32'sd191759, -32'sd1485808, -32'sd538572, 32'sd878805, 32'sd185836, 32'sd1131295, -32'sd1932305, -32'sd645416, -32'sd767320, -32'sd2457504, -32'sd1890726, -32'sd4891302, -32'sd6131829, -32'sd3510616, -32'sd860965, 32'sd404632, 32'sd2731323, 32'sd1930380, 32'sd2338443, 32'sd1557600, -32'sd1516147, -32'sd1317496, -32'sd2501852, 32'sd91325, 32'sd654706, 32'sd1001606, -32'sd1116609, -32'sd1485045, -32'sd397711, -32'sd612769, -32'sd645614, 32'sd2113586, 32'sd1578130, -32'sd1707752, -32'sd280118, -32'sd15925, -32'sd1691183, -32'sd2058612, -32'sd2265726, -32'sd4172147, -32'sd5910715, -32'sd4003298, -32'sd2055556, -32'sd1113731, 32'sd2558265, 32'sd2851260, -32'sd409416, -32'sd260432, -32'sd1097281, -32'sd1895586, -32'sd624264, -32'sd1289199, -32'sd1149285, 32'sd412053, -32'sd3055291, -32'sd1505862, -32'sd584903, -32'sd1396951, -32'sd1021385, -32'sd331188, 32'sd251962, -32'sd184989, 32'sd653401, -32'sd732811, -32'sd1703021, -32'sd3600340, -32'sd4026028, -32'sd1800946, -32'sd3099105, -32'sd915236, -32'sd943533, 32'sd501980, 32'sd1898864, 32'sd3907217, 32'sd326224, 32'sd111462, -32'sd353112, -32'sd602588, -32'sd2849667, -32'sd1457802, -32'sd576326, 32'sd1594363, -32'sd2126406, 32'sd1054912, 32'sd2565834, 32'sd156487, -32'sd428377, 32'sd315675, 32'sd1487946, 32'sd119791, 32'sd2176185, -32'sd496811, -32'sd928001, -32'sd1800498, -32'sd1098513, 32'sd896148, -32'sd1073736, -32'sd601835, -32'sd1121886, -32'sd507760, 32'sd498598, -32'sd128469, 32'sd731816, 32'sd822643, 32'sd918579, 32'sd452729, 32'sd231125, -32'sd247206, -32'sd359660, -32'sd1083846, -32'sd1481623, -32'sd1016406, 32'sd901885, -32'sd1483342, -32'sd420062, 32'sd329127, -32'sd171490, -32'sd169100, 32'sd1492817, 32'sd603523, 32'sd716132, -32'sd1727762, 32'sd302103, 32'sd1534774, 32'sd1610868, -32'sd204725, -32'sd1460634, -32'sd74984, 32'sd837015, 32'sd1155919, 32'sd375460, 32'sd1788497, -32'sd339256, 32'sd3267365, 32'sd2072618, 32'sd213685, -32'sd273750, 32'sd1491719, -32'sd675768, -32'sd293679, 32'sd925563, -32'sd610170, 32'sd0, -32'sd433814, 32'sd246491, -32'sd284392, -32'sd707447, -32'sd842558, 32'sd634312, 32'sd2186116, 32'sd693270, 32'sd2593540, 32'sd42129, 32'sd898313, -32'sd2517928, -32'sd2061481, -32'sd337784, 32'sd3181948, 32'sd1848457, 32'sd619497, 32'sd2057492, 32'sd1065741, 32'sd1279546, 32'sd725782, 32'sd450281, 32'sd1417654, -32'sd999899, 32'sd1367518, -32'sd94574, -32'sd837035, 32'sd96007, 32'sd711084, 32'sd54542, 32'sd32950, 32'sd138190, 32'sd842766, 32'sd269021, 32'sd1385511, 32'sd884091, 32'sd1979022, 32'sd425769, -32'sd852349, -32'sd1754175, -32'sd1148056, 32'sd1644317, 32'sd1460339, 32'sd1023147, 32'sd1498842, -32'sd38504, 32'sd1972315, 32'sd4086836, 32'sd953545, -32'sd1242950, -32'sd801859, 32'sd1900231, -32'sd351517, 32'sd2118935, 32'sd1772572, -32'sd794231, 32'sd634832, 32'sd309014, 32'sd1325243, 32'sd2458278, 32'sd660675, 32'sd588973, 32'sd2486170, 32'sd2500209, 32'sd984834, 32'sd75801, -32'sd679478, -32'sd1701474, -32'sd1414432, -32'sd332021, -32'sd638713, 32'sd374821, -32'sd14276, 32'sd1155918, 32'sd1754121, 32'sd2013427, 32'sd323640, -32'sd988684, -32'sd69037, 32'sd1775499, 32'sd1031417, 32'sd612328, 32'sd1131140, 32'sd0, -32'sd279891, -32'sd464067, -32'sd337521, 32'sd242070, -32'sd494583, -32'sd163519, 32'sd1521961, 32'sd723168, -32'sd1640554, -32'sd1283855, -32'sd3696357, -32'sd2046903, -32'sd193849, -32'sd3034445, -32'sd47349, 32'sd609873, 32'sd369853, -32'sd575966, 32'sd2411451, 32'sd563835, -32'sd1715754, -32'sd747564, -32'sd2563433, 32'sd643933, 32'sd1134659, 32'sd1417475, -32'sd241386, 32'sd1558484, -32'sd577217, -32'sd63930, -32'sd14524, 32'sd1297249, -32'sd920453, 32'sd929376, -32'sd64525, 32'sd496181, -32'sd84737, -32'sd1601546, -32'sd2971374, -32'sd776278, -32'sd343973, -32'sd19219, -32'sd1863429, -32'sd1155516, 32'sd52991, -32'sd799008, -32'sd140988, -32'sd227130, -32'sd867806, -32'sd2267253, -32'sd1522327, 32'sd878138, -32'sd186645, 32'sd254348, 32'sd189132, 32'sd791030, 32'sd827108, -32'sd1637207, -32'sd737009, 32'sd1397826, 32'sd461396, -32'sd900294, 32'sd1068674, -32'sd869987, -32'sd1995383, -32'sd961441, 32'sd645957, -32'sd2228419, -32'sd279396, 32'sd233580, 32'sd70530, -32'sd1650565, 32'sd1601900, 32'sd284017, -32'sd1650497, -32'sd2982316, 32'sd894296, -32'sd2097136, -32'sd1957677, -32'sd1376001, -32'sd161228, 32'sd38272, -32'sd958388, 32'sd0, 32'sd237469, -32'sd989705, -32'sd721096, 32'sd496013, 32'sd408979, 32'sd181809, -32'sd258659, 32'sd981541, -32'sd864276, 32'sd776016, -32'sd1100356, -32'sd1328713, -32'sd1401372, 32'sd31236, 32'sd984758, 32'sd1885273, 32'sd2399515, -32'sd2403751, -32'sd1957211, -32'sd179328, -32'sd1319760, -32'sd1503815, 32'sd45315, -32'sd1783626, 32'sd291380, -32'sd971793, 32'sd0, 32'sd0, 32'sd0, -32'sd924018, 32'sd552723, -32'sd1126766, -32'sd1582045, 32'sd158436, -32'sd2241561, 32'sd470939, 32'sd222565, 32'sd791736, 32'sd560145, 32'sd1929705, 32'sd1432002, -32'sd2098216, -32'sd430593, 32'sd1597888, -32'sd1330328, -32'sd1210078, -32'sd3241463, -32'sd662235, 32'sd295173, 32'sd426779, 32'sd240085, -32'sd1391088, 32'sd223267, -32'sd749037, 32'sd0, 32'sd0, 32'sd0, -32'sd571587, 32'sd978575, -32'sd473864, 32'sd783973, 32'sd1414714, 32'sd442067, 32'sd660299, 32'sd535857, 32'sd963659, 32'sd777659, 32'sd2224313, 32'sd588108, 32'sd1569018, 32'sd1062164, -32'sd1847135, -32'sd1288661, -32'sd2081892, -32'sd298528, 32'sd577051, 32'sd324666, 32'sd398753, -32'sd685426, -32'sd624069, 32'sd1194095, 32'sd510832, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd327176, 32'sd133835, -32'sd1006920, -32'sd112049, 32'sd310694, -32'sd1004551, 32'sd15441, 32'sd1090754, -32'sd585690, -32'sd2330605, -32'sd342929, 32'sd623126, -32'sd2498085, -32'sd1767909, -32'sd2798954, -32'sd711819, 32'sd489793, -32'sd525454, -32'sd23065, -32'sd18019, 32'sd173740, 32'sd790578, 32'sd345305, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd489306, 32'sd1505912, -32'sd946669, -32'sd516675, 32'sd1182241, -32'sd550901, -32'sd1194991, -32'sd770041, 32'sd460430, -32'sd1018293, -32'sd1676973, -32'sd1257772, -32'sd383629, 32'sd892745, -32'sd705426, -32'sd432986, -32'sd1121204, 32'sd96238, 32'sd345794, 32'sd457679, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1208395, -32'sd10924, 32'sd2159044, -32'sd79869, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd461536, 32'sd1549323, 32'sd605630, -32'sd506403, 32'sd592965, 32'sd1134320, 32'sd325827, -32'sd480730, 32'sd158295, -32'sd67348, 32'sd813468, 32'sd1183703, 32'sd400862, 32'sd446683, -32'sd213409, 32'sd600443, 32'sd354851, -32'sd916110, 32'sd252246, -32'sd6643, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1169601, 32'sd302015, -32'sd1082533, 32'sd706278, 32'sd987042, -32'sd1194772, -32'sd454551, -32'sd558375, 32'sd2339577, -32'sd802999, 32'sd1816902, 32'sd2505042, 32'sd2144486, 32'sd1425619, 32'sd2915847, 32'sd1776178, 32'sd633290, -32'sd409211, 32'sd280680, -32'sd59943, 32'sd217140, 32'sd653901, 32'sd362151, 32'sd428797, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1385456, 32'sd191147, 32'sd807229, -32'sd2264630, -32'sd132383, -32'sd1451400, 32'sd372892, 32'sd95355, 32'sd304723, -32'sd512374, 32'sd536867, 32'sd1158219, -32'sd690847, 32'sd3037320, 32'sd1983609, 32'sd1864478, -32'sd885957, 32'sd811090, 32'sd230150, -32'sd98866, -32'sd251909, 32'sd981876, -32'sd237248, -32'sd342418, 32'sd465618, 32'sd0, 32'sd0, 32'sd886151, -32'sd876328, 32'sd812240, -32'sd673706, -32'sd841844, -32'sd1035608, -32'sd776601, -32'sd2362941, -32'sd2950453, -32'sd1536526, 32'sd1169947, 32'sd1507500, -32'sd48443, 32'sd2773057, 32'sd1666072, 32'sd2910008, 32'sd211309, 32'sd969920, 32'sd1600315, -32'sd686160, -32'sd1913257, 32'sd25402, -32'sd1012677, -32'sd2578851, -32'sd1219707, -32'sd146255, 32'sd13968, 32'sd0, 32'sd1273695, 32'sd265401, 32'sd416365, 32'sd634595, -32'sd850953, -32'sd1037104, -32'sd1722462, -32'sd1064819, -32'sd1857863, -32'sd2120536, -32'sd1373533, 32'sd352510, 32'sd428459, 32'sd2034408, 32'sd1826396, 32'sd2631710, -32'sd303821, 32'sd2132155, 32'sd1833733, 32'sd46875, -32'sd759457, 32'sd1876253, 32'sd153237, -32'sd1725834, 32'sd696048, -32'sd1333756, -32'sd168586, 32'sd0, -32'sd59354, 32'sd788668, -32'sd74202, 32'sd255423, -32'sd1329872, -32'sd1416395, 32'sd433551, -32'sd1236819, -32'sd1135783, -32'sd744941, -32'sd2412231, -32'sd1375186, -32'sd1455102, -32'sd1474011, 32'sd2811079, 32'sd999542, -32'sd805134, 32'sd2521121, 32'sd491378, 32'sd599046, 32'sd692212, -32'sd1194635, -32'sd191114, 32'sd103235, 32'sd1128320, -32'sd2101722, 32'sd714398, 32'sd191117, -32'sd272369, 32'sd746308, 32'sd1464429, -32'sd426240, -32'sd678340, -32'sd1320237, -32'sd499502, -32'sd1784039, 32'sd864035, -32'sd2178313, -32'sd3271251, -32'sd4553307, -32'sd2755073, -32'sd657290, 32'sd1547766, 32'sd1968129, 32'sd1554308, 32'sd1756293, 32'sd3154421, 32'sd691483, -32'sd67826, 32'sd1171864, -32'sd1090838, -32'sd2209128, 32'sd705010, -32'sd664334, -32'sd476071, 32'sd604267, 32'sd2138719, -32'sd142194, -32'sd381946, -32'sd1010592, 32'sd1080600, 32'sd1115911, -32'sd1115495, -32'sd2051354, -32'sd133592, -32'sd2508250, -32'sd5233357, -32'sd5587137, -32'sd3805086, -32'sd795067, 32'sd442415, 32'sd1300056, 32'sd2585751, -32'sd59092, 32'sd874109, -32'sd159767, -32'sd1099503, -32'sd1362477, 32'sd338792, -32'sd1185507, -32'sd147104, -32'sd383159, 32'sd832384, -32'sd998050, 32'sd1447583, -32'sd474035, 32'sd1739332, 32'sd1191247, 32'sd355930, -32'sd1047077, -32'sd1278849, 32'sd1023015, 32'sd2067811, -32'sd947780, -32'sd3699926, -32'sd3898555, -32'sd1568094, 32'sd1922020, 32'sd2254425, 32'sd1215592, 32'sd1110179, 32'sd3385928, 32'sd1190514, -32'sd485605, -32'sd1698480, -32'sd1063332, -32'sd431643, -32'sd925039, -32'sd840744, -32'sd1219495, 32'sd40477, 32'sd557748, 32'sd301298, 32'sd884250, -32'sd1283882, 32'sd266552, -32'sd1083608, 32'sd1321478, -32'sd901035, 32'sd289641, 32'sd1150478, -32'sd219240, -32'sd237576, -32'sd1721955, -32'sd936677, 32'sd340333, 32'sd2630916, 32'sd2337739, 32'sd2900844, 32'sd172455, -32'sd1070767, -32'sd997544, 32'sd102268, -32'sd2742366, 32'sd829740, -32'sd1339757, 32'sd151715, -32'sd360740, 32'sd533831, 32'sd126131, 32'sd1372596, 32'sd1306839, 32'sd2006937, -32'sd933088, 32'sd1266994, 32'sd1385715, 32'sd1522134, 32'sd1722937, 32'sd2355485, 32'sd470224, -32'sd2074793, -32'sd2241790, -32'sd1540940, 32'sd1846628, 32'sd1222753, 32'sd1949174, 32'sd2142618, -32'sd604100, 32'sd929758, 32'sd1058359, -32'sd835411, -32'sd1213569, 32'sd213435, -32'sd3531112, 32'sd205864, -32'sd609351, 32'sd323908, 32'sd329855, 32'sd266860, 32'sd643651, 32'sd971893, 32'sd832083, 32'sd1557308, 32'sd682813, 32'sd1556269, 32'sd602996, 32'sd3194732, -32'sd42805, -32'sd843836, -32'sd621116, -32'sd443351, 32'sd1067401, 32'sd752293, 32'sd2909488, 32'sd159946, 32'sd352879, 32'sd705312, 32'sd70215, 32'sd340092, -32'sd2137919, 32'sd72908, -32'sd1600235, -32'sd580249, 32'sd416013, 32'sd133536, 32'sd837880, -32'sd1279739, -32'sd517051, 32'sd1060212, 32'sd1497067, -32'sd18692, 32'sd1459728, -32'sd215559, -32'sd1108363, 32'sd2750893, 32'sd563852, -32'sd602293, -32'sd2176847, -32'sd2184032, 32'sd921518, 32'sd38376, 32'sd274656, 32'sd1495595, 32'sd1687612, -32'sd1701418, -32'sd598422, -32'sd545821, -32'sd2534972, -32'sd2358046, -32'sd256424, -32'sd864386, -32'sd920120, -32'sd13440, 32'sd1114954, 32'sd49546, -32'sd549275, 32'sd320030, 32'sd1136119, 32'sd2410207, 32'sd157320, -32'sd5556, 32'sd765038, 32'sd622764, -32'sd1159655, -32'sd1950537, -32'sd759365, -32'sd792160, 32'sd3403849, 32'sd1455645, 32'sd3876094, -32'sd559034, 32'sd238217, -32'sd95246, -32'sd2313531, -32'sd1395169, -32'sd1889130, -32'sd3034073, 32'sd292912, 32'sd1159024, 32'sd1199426, 32'sd1217739, -32'sd696433, 32'sd1072009, -32'sd422838, 32'sd1084247, 32'sd778908, -32'sd478165, 32'sd925207, -32'sd379451, -32'sd782810, -32'sd2850460, -32'sd3825118, 32'sd1163638, 32'sd349308, 32'sd43645, 32'sd2233680, 32'sd1795756, 32'sd1075384, -32'sd1718663, -32'sd1613771, 32'sd324781, -32'sd500765, -32'sd1088141, -32'sd3013451, -32'sd2127804, -32'sd953158, -32'sd1177861, -32'sd937835, 32'sd953293, 32'sd622366, 32'sd563416, 32'sd943701, 32'sd17440, -32'sd505750, -32'sd1876000, 32'sd557633, -32'sd1367967, -32'sd2532922, -32'sd3289838, -32'sd2476785, 32'sd163378, -32'sd1950761, 32'sd1333584, -32'sd267968, -32'sd58697, -32'sd1956524, -32'sd2802076, -32'sd3158, 32'sd124235, -32'sd674806, 32'sd455742, -32'sd2246857, -32'sd1074082, 32'sd2047183, -32'sd1304891, 32'sd804343, -32'sd811311, 32'sd0, 32'sd859408, 32'sd1642494, 32'sd354630, 32'sd1576749, 32'sd1127062, -32'sd710681, -32'sd885349, -32'sd2404085, -32'sd1649366, -32'sd420775, 32'sd520660, 32'sd395083, -32'sd432998, -32'sd193415, 32'sd966939, -32'sd1096744, -32'sd1258285, 32'sd132639, 32'sd264545, -32'sd293060, 32'sd959559, -32'sd148346, 32'sd754674, 32'sd3085914, 32'sd2269683, -32'sd284907, -32'sd781032, 32'sd439726, -32'sd489376, 32'sd1546922, 32'sd459504, 32'sd121966, -32'sd470478, -32'sd456866, 32'sd783745, 32'sd525733, 32'sd459559, 32'sd448709, -32'sd874194, 32'sd473115, 32'sd1430132, 32'sd309336, 32'sd183027, -32'sd534692, -32'sd1588622, -32'sd877143, 32'sd313266, 32'sd1100783, 32'sd861022, 32'sd89393, 32'sd1090998, 32'sd2379247, 32'sd2863134, 32'sd341938, 32'sd874960, 32'sd1664367, -32'sd566169, -32'sd63735, -32'sd902509, 32'sd349539, -32'sd1265048, -32'sd156642, 32'sd532953, -32'sd414081, 32'sd2530788, 32'sd706848, 32'sd352901, -32'sd1369381, 32'sd1893440, -32'sd102757, -32'sd565735, 32'sd431181, -32'sd133408, -32'sd525218, -32'sd163575, 32'sd1881164, 32'sd1131452, -32'sd144188, 32'sd1021505, 32'sd1094309, 32'sd1318555, -32'sd1031920, 32'sd853206, 32'sd0, -32'sd66449, -32'sd635577, 32'sd1852410, 32'sd2020524, -32'sd1087067, 32'sd2520302, 32'sd1739829, 32'sd1192997, 32'sd276034, 32'sd1298428, 32'sd65180, 32'sd172286, -32'sd227082, -32'sd2126802, -32'sd1579400, 32'sd2362279, 32'sd1791828, 32'sd3080802, -32'sd858707, 32'sd412962, -32'sd383952, 32'sd699853, 32'sd182271, 32'sd2338917, 32'sd296284, -32'sd163686, -32'sd83270, 32'sd973570, 32'sd945157, 32'sd780734, 32'sd1275167, -32'sd427936, -32'sd1270723, 32'sd1182131, 32'sd1606426, 32'sd1638928, -32'sd438702, -32'sd212016, -32'sd622055, -32'sd1133431, -32'sd343231, 32'sd211304, -32'sd220226, -32'sd1036994, -32'sd363995, -32'sd346793, -32'sd394286, -32'sd488245, -32'sd937514, -32'sd114025, -32'sd1571428, 32'sd1078535, 32'sd748898, 32'sd1034483, 32'sd9822, 32'sd2066925, 32'sd1058860, 32'sd1461232, -32'sd806050, 32'sd541000, 32'sd2334361, 32'sd1079310, 32'sd1028484, 32'sd657240, 32'sd334040, -32'sd1200416, 32'sd1372901, -32'sd204925, -32'sd1317182, 32'sd1501121, -32'sd548565, 32'sd632165, 32'sd591500, 32'sd729398, -32'sd1347331, -32'sd922963, 32'sd1042245, -32'sd337847, -32'sd567762, -32'sd1552778, -32'sd176984, -32'sd102549, 32'sd77393, 32'sd0, -32'sd918943, -32'sd271190, 32'sd1244855, 32'sd1461496, 32'sd831857, 32'sd840489, -32'sd1640192, -32'sd895926, 32'sd1017892, 32'sd721640, -32'sd143358, 32'sd513459, 32'sd2438670, 32'sd2765677, 32'sd2032144, 32'sd1071901, 32'sd133769, 32'sd59862, -32'sd21438, 32'sd544595, -32'sd282495, -32'sd841723, -32'sd993858, -32'sd1416322, 32'sd423470, 32'sd1299186, 32'sd0, 32'sd0, 32'sd0, -32'sd954999, -32'sd10908, 32'sd1311334, 32'sd913639, -32'sd915489, -32'sd1310534, -32'sd1474914, -32'sd1473648, -32'sd1551993, 32'sd321274, -32'sd721472, 32'sd692548, 32'sd2757033, 32'sd1591458, -32'sd592672, -32'sd1714366, 32'sd1588308, 32'sd1834785, 32'sd998655, -32'sd637923, -32'sd1623534, -32'sd1222325, -32'sd1075203, 32'sd698504, 32'sd1222373, 32'sd0, 32'sd0, 32'sd0, -32'sd188676, 32'sd444666, 32'sd553368, 32'sd170345, -32'sd407862, -32'sd1743077, 32'sd1331620, 32'sd1392561, -32'sd3007845, -32'sd2339750, 32'sd222400, -32'sd1189000, -32'sd890448, -32'sd1923069, -32'sd2007688, 32'sd2567782, 32'sd2365602, 32'sd794183, -32'sd1837965, -32'sd936863, -32'sd421633, -32'sd1316187, -32'sd1088140, 32'sd1053521, -32'sd511412, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd194164, 32'sd312054, -32'sd888679, 32'sd275774, 32'sd868062, 32'sd217181, -32'sd1505733, 32'sd706655, 32'sd1033332, 32'sd921579, -32'sd137874, -32'sd668091, -32'sd909601, 32'sd1420944, -32'sd1995754, -32'sd1552079, -32'sd2064163, -32'sd1835965, -32'sd1153202, -32'sd345092, 32'sd540755, 32'sd777740, 32'sd1673057, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1088444, 32'sd397521, 32'sd1046975, 32'sd503028, -32'sd504284, -32'sd757350, 32'sd5886, -32'sd1450631, -32'sd625525, -32'sd836058, 32'sd83890, 32'sd201644, 32'sd1745673, 32'sd1585338, 32'sd1140166, 32'sd69405, -32'sd645090, 32'sd868911, -32'sd1034620, -32'sd303680, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1085978, 32'sd1243733, -32'sd766512, 32'sd379868, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd417868, 32'sd1009097, -32'sd555284, 32'sd1289878, 32'sd1303138, 32'sd1358466, 32'sd1051576, 32'sd1542991, 32'sd1609420, -32'sd296898, -32'sd703151, 32'sd1007107, 32'sd1286186, -32'sd429316, 32'sd582786, -32'sd598087, -32'sd1284343, -32'sd975922, -32'sd724648, 32'sd785743, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd465145, -32'sd751193, -32'sd369304, 32'sd1805360, -32'sd132152, -32'sd814787, 32'sd1032944, 32'sd1416320, -32'sd504585, 32'sd1888493, 32'sd753723, 32'sd2267490, 32'sd1610269, 32'sd758537, 32'sd461602, -32'sd1291648, -32'sd2087177, 32'sd734778, 32'sd1291342, -32'sd894196, -32'sd8917, 32'sd489256, 32'sd1080749, 32'sd430235, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd348801, 32'sd47539, -32'sd681074, 32'sd525630, 32'sd1432801, -32'sd385875, 32'sd1495001, 32'sd3121103, 32'sd1631495, -32'sd1428605, -32'sd401560, 32'sd727525, 32'sd1585682, -32'sd87145, -32'sd1148110, -32'sd604405, -32'sd50770, 32'sd20920, -32'sd1455910, -32'sd1139578, 32'sd160825, -32'sd1300045, 32'sd278123, 32'sd993090, -32'sd397556, 32'sd0, 32'sd0, -32'sd255890, 32'sd126947, 32'sd367610, -32'sd1707701, 32'sd424208, 32'sd1872771, 32'sd1301213, 32'sd395141, -32'sd1445806, -32'sd341785, -32'sd527243, 32'sd1680941, 32'sd239462, 32'sd1137058, -32'sd100115, -32'sd2310494, -32'sd1395052, -32'sd2560962, -32'sd2652738, -32'sd1948330, -32'sd1709963, -32'sd2244177, -32'sd2080261, 32'sd362548, -32'sd22101, -32'sd1504718, -32'sd703798, 32'sd0, 32'sd606760, -32'sd512209, -32'sd957964, 32'sd6548, 32'sd135960, 32'sd1476646, -32'sd1868509, -32'sd1627901, -32'sd247347, -32'sd43122, 32'sd660620, 32'sd2722744, 32'sd2344679, -32'sd571870, 32'sd155114, -32'sd238460, -32'sd1230502, -32'sd809318, -32'sd2044931, -32'sd470502, -32'sd1660469, -32'sd1918634, 32'sd399605, 32'sd657843, 32'sd135913, -32'sd858581, -32'sd242098, 32'sd0, -32'sd776079, 32'sd65244, 32'sd418494, -32'sd397011, -32'sd778899, -32'sd1517591, -32'sd1295868, -32'sd826691, 32'sd1413289, -32'sd256331, -32'sd416691, 32'sd2251105, 32'sd1192100, 32'sd1292845, -32'sd440245, -32'sd656057, 32'sd83467, 32'sd126103, -32'sd1392650, -32'sd1425400, 32'sd781291, -32'sd1617399, -32'sd416853, -32'sd2151411, -32'sd1973058, 32'sd1669936, -32'sd673532, -32'sd287816, 32'sd1537991, -32'sd1102779, 32'sd1049129, 32'sd920323, -32'sd1383138, -32'sd1848560, -32'sd1674582, 32'sd1939153, 32'sd1551641, -32'sd461592, -32'sd451759, 32'sd35603, 32'sd166014, -32'sd462804, -32'sd625436, -32'sd495413, -32'sd133413, 32'sd2037967, 32'sd146083, -32'sd1086158, -32'sd304808, -32'sd1095954, -32'sd1555229, -32'sd1113076, -32'sd938851, -32'sd723159, 32'sd429532, -32'sd758108, -32'sd546191, 32'sd212639, -32'sd138586, -32'sd90310, 32'sd520432, -32'sd1436969, 32'sd304747, 32'sd3044647, -32'sd261346, -32'sd532086, -32'sd3160775, -32'sd1998711, -32'sd2561171, 32'sd413024, 32'sd553893, -32'sd665284, 32'sd935018, -32'sd66423, -32'sd1462454, -32'sd1451606, -32'sd952971, -32'sd771107, -32'sd565063, -32'sd590205, -32'sd923836, -32'sd1781102, -32'sd884466, 32'sd1573267, 32'sd277398, -32'sd3536375, -32'sd270850, -32'sd99499, 32'sd1602959, 32'sd2100805, -32'sd496836, 32'sd3516156, -32'sd7102, -32'sd1523316, -32'sd2010680, -32'sd3582134, -32'sd1426762, 32'sd2174127, 32'sd1333520, 32'sd1206999, 32'sd2059028, 32'sd902996, -32'sd1144404, -32'sd1132133, 32'sd424418, -32'sd877358, 32'sd512413, -32'sd701307, -32'sd95468, -32'sd2056339, -32'sd157050, 32'sd502403, 32'sd211240, -32'sd1466025, -32'sd3256125, 32'sd551005, 32'sd2256194, 32'sd1046598, 32'sd2638421, 32'sd3101237, 32'sd1671242, -32'sd546840, -32'sd1120809, -32'sd3023021, -32'sd1131561, 32'sd821172, -32'sd81806, 32'sd1478620, -32'sd1448902, 32'sd1580428, 32'sd2273976, 32'sd1581738, -32'sd882554, 32'sd1443787, -32'sd320646, 32'sd1249292, -32'sd516006, -32'sd1359262, -32'sd497067, 32'sd137543, -32'sd1417030, -32'sd364051, -32'sd1198633, -32'sd374776, 32'sd178684, 32'sd2184305, 32'sd975335, 32'sd357550, -32'sd752, 32'sd1133105, 32'sd1144431, 32'sd864386, 32'sd28668, -32'sd759520, 32'sd126428, 32'sd1099336, 32'sd1790493, 32'sd2177346, 32'sd2202179, 32'sd3281286, 32'sd287367, 32'sd1603711, 32'sd1127703, -32'sd2331292, 32'sd120068, 32'sd426834, -32'sd485561, 32'sd644657, -32'sd551402, 32'sd46267, 32'sd444118, -32'sd1887133, 32'sd918681, -32'sd1131724, 32'sd687988, 32'sd1286495, 32'sd559026, 32'sd1850384, 32'sd1484672, 32'sd519943, 32'sd41103, -32'sd128526, 32'sd1793144, -32'sd204477, 32'sd1060838, 32'sd2917482, 32'sd1663636, 32'sd538761, -32'sd61883, 32'sd1024336, -32'sd627004, 32'sd2374005, -32'sd198548, -32'sd848210, -32'sd1053232, 32'sd696235, -32'sd1393412, 32'sd635156, -32'sd595353, -32'sd1844670, -32'sd113501, -32'sd538109, 32'sd1945979, 32'sd1281228, -32'sd38277, 32'sd2002664, -32'sd1707102, -32'sd2703725, -32'sd3130495, -32'sd1043621, -32'sd43738, 32'sd1964306, 32'sd1215601, -32'sd12706, 32'sd961256, -32'sd1697450, -32'sd233626, -32'sd960723, -32'sd1052051, 32'sd274430, -32'sd2006403, -32'sd1369782, -32'sd630436, -32'sd205908, -32'sd543019, 32'sd1660742, -32'sd2143596, -32'sd3269693, -32'sd1970064, -32'sd286131, 32'sd453136, 32'sd697485, -32'sd205957, 32'sd1747121, 32'sd451596, -32'sd1241244, -32'sd3164505, 32'sd807291, 32'sd2916194, 32'sd4089903, 32'sd1102610, 32'sd1792686, -32'sd70896, -32'sd1256078, -32'sd603589, 32'sd190607, 32'sd1729737, -32'sd1073748, -32'sd1396896, -32'sd123636, 32'sd118465, 32'sd277644, -32'sd785326, -32'sd756511, -32'sd606912, -32'sd2543706, -32'sd1128531, 32'sd338196, -32'sd1167798, -32'sd1022086, -32'sd2586379, -32'sd173000, -32'sd1970533, -32'sd3227775, -32'sd2586275, -32'sd1037216, 32'sd425701, 32'sd1704649, 32'sd1923709, -32'sd386408, -32'sd86122, 32'sd1253274, -32'sd1474241, 32'sd355121, 32'sd1350008, 32'sd289251, -32'sd1198073, 32'sd1188516, -32'sd796707, 32'sd267742, 32'sd1235143, 32'sd1736022, 32'sd481955, 32'sd381620, -32'sd308347, 32'sd42176, -32'sd1121590, -32'sd584628, -32'sd1519511, -32'sd1343244, -32'sd458149, -32'sd722387, -32'sd1902908, -32'sd429054, 32'sd1077809, 32'sd3363612, 32'sd2124795, -32'sd1256060, -32'sd356036, -32'sd926114, -32'sd2733705, -32'sd522358, 32'sd933248, 32'sd1060561, 32'sd1216029, 32'sd67913, 32'sd699624, 32'sd0, -32'sd471118, 32'sd244368, -32'sd1915477, -32'sd1037360, 32'sd724014, -32'sd490803, -32'sd2361883, -32'sd1662371, -32'sd3151617, -32'sd2152646, 32'sd381705, -32'sd1339487, -32'sd965411, -32'sd1086742, 32'sd1445691, 32'sd1769631, 32'sd1279645, 32'sd2482334, -32'sd1990702, -32'sd1880822, -32'sd518140, -32'sd2238005, -32'sd1217132, -32'sd203605, 32'sd918220, -32'sd460537, 32'sd256927, -32'sd955030, 32'sd892046, -32'sd1358425, 32'sd351254, -32'sd2816978, -32'sd318299, 32'sd1132903, 32'sd551342, 32'sd422801, -32'sd2202453, -32'sd1604130, -32'sd881356, -32'sd2100762, -32'sd1529148, -32'sd121418, 32'sd2065072, 32'sd1130132, 32'sd2015007, 32'sd1491927, -32'sd992664, -32'sd1625486, -32'sd537712, -32'sd1302059, -32'sd3260442, -32'sd135729, 32'sd1845476, 32'sd730237, -32'sd730100, -32'sd66660, 32'sd564313, -32'sd904869, 32'sd618298, -32'sd3807838, 32'sd509500, -32'sd820293, 32'sd930229, -32'sd1740771, -32'sd2019319, -32'sd256958, -32'sd41256, -32'sd1094203, 32'sd1080491, 32'sd1231322, -32'sd209724, 32'sd942528, -32'sd297113, 32'sd257077, 32'sd198811, -32'sd2274462, -32'sd198480, -32'sd561014, -32'sd556675, -32'sd1030601, -32'sd282384, -32'sd1046482, -32'sd99945, 32'sd0, -32'sd184764, 32'sd528377, -32'sd593155, -32'sd3312309, -32'sd2057483, -32'sd692654, 32'sd901815, -32'sd1287864, -32'sd350336, -32'sd679732, 32'sd706172, -32'sd525632, -32'sd2158091, -32'sd1383171, 32'sd223792, 32'sd252321, -32'sd342096, -32'sd892914, -32'sd1357022, -32'sd60971, -32'sd1048855, -32'sd882756, -32'sd972529, 32'sd1711102, 32'sd1531604, 32'sd605126, -32'sd157430, -32'sd775527, -32'sd211742, -32'sd1864363, 32'sd573862, 32'sd62202, -32'sd9987, -32'sd981373, -32'sd1640124, 32'sd342873, 32'sd1209773, 32'sd496019, 32'sd1539456, 32'sd759661, -32'sd1414209, -32'sd329937, -32'sd2171340, 32'sd873476, -32'sd314605, -32'sd1445569, 32'sd468001, 32'sd13799, -32'sd340883, -32'sd936317, 32'sd565477, 32'sd1319685, 32'sd498968, -32'sd1103214, -32'sd676563, -32'sd92627, -32'sd154201, -32'sd740666, 32'sd268183, 32'sd563410, -32'sd1326481, -32'sd1684754, -32'sd319950, -32'sd211398, -32'sd4072, 32'sd2034330, 32'sd1142799, 32'sd1627810, -32'sd921170, 32'sd179168, -32'sd2293392, -32'sd1265115, -32'sd871891, -32'sd341096, 32'sd170815, -32'sd695505, 32'sd659723, 32'sd491038, -32'sd1100513, 32'sd724298, -32'sd2347642, -32'sd396794, -32'sd22430, 32'sd0, -32'sd393747, -32'sd951221, -32'sd964478, -32'sd1373871, -32'sd736098, -32'sd394289, -32'sd407400, -32'sd475649, 32'sd594272, 32'sd1447773, 32'sd1357090, -32'sd247333, 32'sd376982, -32'sd1127834, 32'sd114191, -32'sd1468054, 32'sd349858, -32'sd1058608, 32'sd754655, 32'sd1066690, 32'sd1238471, 32'sd1170897, 32'sd606761, 32'sd683481, 32'sd445967, -32'sd576506, 32'sd0, 32'sd0, 32'sd0, 32'sd344042, -32'sd105114, -32'sd45301, 32'sd381023, -32'sd355614, -32'sd371736, -32'sd463221, -32'sd302465, 32'sd1755655, 32'sd13239, 32'sd834957, -32'sd2573011, 32'sd265525, 32'sd769633, 32'sd77416, -32'sd1110944, -32'sd1623346, 32'sd1513415, 32'sd1502902, -32'sd1289698, 32'sd421219, -32'sd586667, 32'sd26637, 32'sd625953, -32'sd415251, 32'sd0, 32'sd0, 32'sd0, 32'sd1251221, 32'sd164107, 32'sd936930, 32'sd114480, 32'sd216473, -32'sd1410543, 32'sd1301852, 32'sd1428157, -32'sd202589, 32'sd1289006, 32'sd1162729, -32'sd1795618, 32'sd1548421, -32'sd2225997, -32'sd91938, -32'sd1123552, 32'sd367372, -32'sd1431882, -32'sd211691, -32'sd838987, -32'sd998301, 32'sd379240, -32'sd487976, 32'sd217584, -32'sd423323, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd442729, 32'sd1126298, -32'sd1874259, -32'sd2363875, 32'sd167555, 32'sd851809, 32'sd1601244, 32'sd1396991, -32'sd704800, 32'sd838302, -32'sd270998, 32'sd517850, -32'sd660601, 32'sd587247, 32'sd1906620, -32'sd117769, -32'sd640388, 32'sd191863, -32'sd1491224, 32'sd347593, 32'sd84867, -32'sd1394599, 32'sd751110, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd851984, 32'sd87665, -32'sd612986, -32'sd333253, -32'sd668399, -32'sd189633, -32'sd1121183, -32'sd779706, -32'sd814272, 32'sd720133, 32'sd867775, -32'sd636253, -32'sd569633, 32'sd363650, 32'sd1448278, 32'sd1906685, -32'sd472770, 32'sd365625, 32'sd1275250, 32'sd700449, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd44622, 32'sd1020349, 32'sd441010, 32'sd720637, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1743352, 32'sd507, -32'sd578489, -32'sd185276, 32'sd1096603, -32'sd192093, -32'sd421184, 32'sd94250, 32'sd387410, 32'sd433418, -32'sd804112, -32'sd985086, 32'sd2330851, 32'sd1223742, 32'sd1694179, 32'sd2622395, 32'sd1785402, 32'sd1915137, 32'sd2503954, 32'sd1077518, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2196942, 32'sd1591636, 32'sd467721, 32'sd1116664, 32'sd804254, -32'sd1603197, 32'sd276509, -32'sd1137206, -32'sd1771502, 32'sd1825824, 32'sd687063, -32'sd735871, 32'sd158161, -32'sd1250087, -32'sd1281764, 32'sd36281, 32'sd1467407, 32'sd631354, 32'sd88431, 32'sd1990131, 32'sd2342440, 32'sd1843929, -32'sd380251, 32'sd1915314, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1889375, -32'sd565165, 32'sd397044, -32'sd300476, -32'sd135560, -32'sd442863, 32'sd815248, -32'sd120986, -32'sd810399, 32'sd891991, 32'sd659058, -32'sd378892, -32'sd907457, -32'sd1991957, -32'sd600149, -32'sd88509, 32'sd559722, 32'sd333934, 32'sd933331, 32'sd31172, 32'sd1012383, 32'sd864476, 32'sd387409, 32'sd987819, 32'sd658145, 32'sd0, 32'sd0, 32'sd1020767, 32'sd1100103, -32'sd179214, 32'sd1559944, 32'sd1167051, -32'sd603937, -32'sd151864, 32'sd763748, -32'sd569719, -32'sd1979512, 32'sd1907139, -32'sd44367, 32'sd1256076, -32'sd1047790, -32'sd1432150, 32'sd539118, 32'sd305710, 32'sd235276, 32'sd1243694, 32'sd1511609, 32'sd1358687, -32'sd1592045, 32'sd194801, 32'sd1344447, -32'sd145695, -32'sd840744, 32'sd479525, 32'sd0, 32'sd539432, 32'sd265651, -32'sd1559815, -32'sd209219, -32'sd1000475, 32'sd174530, 32'sd717757, 32'sd901154, -32'sd154352, -32'sd803731, 32'sd2635435, 32'sd2126020, 32'sd1775700, -32'sd551849, 32'sd321581, 32'sd1541237, 32'sd2761660, 32'sd890497, 32'sd1797053, -32'sd291807, 32'sd255872, -32'sd279381, -32'sd572789, 32'sd1655449, -32'sd1108785, 32'sd786244, 32'sd1237303, 32'sd0, 32'sd428324, 32'sd271987, 32'sd1753716, -32'sd808976, -32'sd513341, -32'sd694778, -32'sd6212, -32'sd269877, 32'sd832323, -32'sd135260, 32'sd1765856, 32'sd1532032, 32'sd813036, -32'sd620267, 32'sd88600, -32'sd121484, 32'sd1031201, 32'sd1388830, 32'sd2173633, 32'sd166065, 32'sd364617, 32'sd339, -32'sd102750, 32'sd496616, 32'sd1211646, 32'sd21819, -32'sd139559, 32'sd1685616, 32'sd1612019, 32'sd100450, -32'sd1235733, 32'sd1069690, 32'sd1300934, 32'sd1555650, 32'sd751218, 32'sd728066, -32'sd1422923, -32'sd1109685, -32'sd1669269, -32'sd2280172, 32'sd247680, 32'sd129070, -32'sd119827, -32'sd1304765, 32'sd571302, 32'sd1908937, 32'sd586338, 32'sd794234, 32'sd322144, 32'sd1642803, 32'sd1364924, 32'sd1982183, 32'sd962752, 32'sd1935832, 32'sd1366715, 32'sd1142725, 32'sd1065872, -32'sd1454414, 32'sd1608105, 32'sd418993, 32'sd710252, 32'sd800009, -32'sd496638, -32'sd142739, -32'sd503930, -32'sd1196777, -32'sd2095591, -32'sd1004187, 32'sd280853, -32'sd998057, 32'sd1009768, 32'sd245888, 32'sd791139, 32'sd698506, 32'sd3040217, 32'sd1723974, 32'sd507206, 32'sd3036441, 32'sd2421976, 32'sd2696440, 32'sd654705, 32'sd344022, -32'sd590268, -32'sd302949, 32'sd841185, 32'sd1657539, 32'sd2135280, -32'sd303003, -32'sd77028, -32'sd1237756, -32'sd1676671, -32'sd3456391, -32'sd811688, -32'sd430330, -32'sd57123, -32'sd2124974, -32'sd1266727, -32'sd1085652, 32'sd592177, -32'sd2782506, 32'sd1350002, 32'sd302393, 32'sd1203571, -32'sd565482, 32'sd1709402, 32'sd1032039, 32'sd2228951, -32'sd595085, 32'sd1104610, 32'sd140212, -32'sd162025, 32'sd1085338, 32'sd186429, 32'sd1631250, 32'sd1923375, -32'sd784070, -32'sd1885882, -32'sd260208, -32'sd1666781, -32'sd3176222, 32'sd112539, -32'sd1069013, -32'sd1386730, 32'sd290036, -32'sd3010207, -32'sd3176834, -32'sd2231012, -32'sd1047894, -32'sd2080241, -32'sd1667975, -32'sd2188473, -32'sd724518, -32'sd2864166, -32'sd1239014, -32'sd1768831, -32'sd292549, -32'sd104254, 32'sd1222020, 32'sd1183363, 32'sd34184, 32'sd1091643, 32'sd1560363, 32'sd599415, -32'sd2074683, -32'sd1695824, -32'sd1908381, -32'sd3635262, -32'sd2288975, -32'sd1312308, -32'sd252638, -32'sd622166, -32'sd861023, -32'sd1393531, -32'sd2986340, -32'sd1313464, -32'sd4832123, -32'sd5374091, -32'sd4484574, -32'sd4506365, -32'sd2503215, -32'sd4804054, -32'sd1766789, -32'sd2614958, -32'sd1555379, -32'sd108112, -32'sd631945, -32'sd1004267, 32'sd367555, 32'sd685251, 32'sd1312826, 32'sd516294, -32'sd1761747, -32'sd1720157, -32'sd1866970, -32'sd837102, -32'sd1575305, 32'sd354588, -32'sd577568, 32'sd1545329, 32'sd228812, -32'sd851235, -32'sd2354229, -32'sd1211411, -32'sd2924660, -32'sd5192798, -32'sd1967770, -32'sd2289897, -32'sd4502031, -32'sd4089621, -32'sd3729539, -32'sd1072186, -32'sd805390, -32'sd399174, 32'sd337063, -32'sd49360, 32'sd612420, 32'sd550920, 32'sd1036402, 32'sd258964, -32'sd3425502, -32'sd1544931, -32'sd303955, 32'sd1167230, -32'sd147886, 32'sd362592, 32'sd384231, -32'sd705384, 32'sd2073746, 32'sd2778800, 32'sd1073785, 32'sd2570903, -32'sd278545, -32'sd432250, -32'sd1344147, -32'sd1162850, -32'sd2452401, -32'sd2707390, -32'sd2715766, -32'sd2182883, 32'sd370255, -32'sd777768, -32'sd607587, 32'sd2106992, 32'sd1618170, -32'sd316150, 32'sd1390570, -32'sd803172, 32'sd1314597, -32'sd124028, 32'sd1049465, 32'sd860936, 32'sd830625, -32'sd559811, 32'sd1233727, -32'sd1004106, -32'sd660627, 32'sd1068321, 32'sd292925, 32'sd3368812, 32'sd795463, 32'sd1120776, 32'sd468804, -32'sd1674259, 32'sd332135, -32'sd1303996, -32'sd1561281, -32'sd2423373, -32'sd517670, 32'sd2045312, 32'sd422132, 32'sd1895067, 32'sd1075691, 32'sd1272574, -32'sd448264, 32'sd710812, 32'sd3000657, 32'sd3112550, 32'sd489845, 32'sd898121, 32'sd1352132, -32'sd621264, -32'sd1583277, -32'sd1329812, -32'sd476192, 32'sd269890, 32'sd1744390, 32'sd240260, 32'sd2695000, 32'sd1829245, 32'sd2085353, -32'sd1139118, -32'sd622529, 32'sd216044, -32'sd2224353, -32'sd420586, -32'sd164728, 32'sd845311, 32'sd1539071, 32'sd742981, 32'sd1105959, -32'sd844263, -32'sd993443, -32'sd21874, 32'sd2834482, 32'sd1374620, -32'sd76097, 32'sd2283032, -32'sd1622363, -32'sd1358191, 32'sd254580, -32'sd744849, 32'sd2907563, 32'sd329823, 32'sd626434, 32'sd273087, -32'sd131327, 32'sd916508, 32'sd175703, 32'sd604862, 32'sd166177, 32'sd1035213, 32'sd1694542, 32'sd246559, 32'sd906018, 32'sd209973, -32'sd1427046, -32'sd124329, 32'sd0, 32'sd549328, -32'sd3027084, 32'sd850692, 32'sd2651561, 32'sd1365669, 32'sd843874, 32'sd1636987, -32'sd203326, 32'sd391224, -32'sd1159699, -32'sd622900, 32'sd702157, -32'sd158357, -32'sd2740647, -32'sd982190, -32'sd125186, 32'sd1367944, 32'sd1436250, 32'sd1334646, 32'sd1629184, 32'sd2000566, 32'sd1147287, -32'sd1016139, -32'sd1309819, -32'sd3181129, -32'sd27883, 32'sd979981, -32'sd214083, 32'sd1289842, -32'sd412909, 32'sd1260329, -32'sd939999, 32'sd1333171, 32'sd2083940, 32'sd820337, 32'sd570232, -32'sd520820, -32'sd1155731, -32'sd622736, 32'sd897249, -32'sd3358273, -32'sd1767294, 32'sd386170, 32'sd725596, 32'sd678522, 32'sd1150526, 32'sd2395034, 32'sd2814018, 32'sd2359944, -32'sd967569, -32'sd1141193, -32'sd1039286, -32'sd671018, 32'sd879002, 32'sd1419483, 32'sd269244, -32'sd1124920, -32'sd906337, 32'sd429391, -32'sd44619, -32'sd2641739, -32'sd298190, -32'sd587822, -32'sd212544, -32'sd689027, -32'sd527519, 32'sd536556, 32'sd111291, -32'sd695548, 32'sd212654, 32'sd203965, 32'sd144000, 32'sd2433565, 32'sd2848901, 32'sd1846668, 32'sd1463430, 32'sd797411, 32'sd319985, 32'sd1879058, 32'sd311783, 32'sd913454, 32'sd1921245, 32'sd452582, 32'sd0, -32'sd717216, 32'sd1158657, 32'sd287770, 32'sd543462, -32'sd1971182, -32'sd1074026, -32'sd728407, -32'sd502445, -32'sd634746, 32'sd1379161, 32'sd525674, -32'sd1507406, 32'sd2005462, -32'sd1043128, -32'sd590392, -32'sd933051, 32'sd2753107, -32'sd612334, 32'sd1060464, -32'sd16585, 32'sd93252, 32'sd1139759, -32'sd2897594, -32'sd627191, -32'sd1738526, 32'sd824507, 32'sd330498, 32'sd190059, -32'sd166715, 32'sd1166125, 32'sd1288898, 32'sd78556, -32'sd445861, 32'sd282, -32'sd882550, -32'sd497120, -32'sd375789, 32'sd2559915, 32'sd722883, -32'sd716071, 32'sd677411, 32'sd382401, -32'sd19263, 32'sd1910545, 32'sd2962241, 32'sd997688, -32'sd1071357, -32'sd442466, -32'sd316977, -32'sd2621516, -32'sd3752402, -32'sd735459, -32'sd982513, 32'sd1159706, 32'sd799123, -32'sd537890, -32'sd1682599, -32'sd130326, -32'sd238917, 32'sd1151662, 32'sd47656, -32'sd1119240, -32'sd464773, 32'sd200909, 32'sd935483, 32'sd1261521, 32'sd1880617, 32'sd1662377, 32'sd2128307, 32'sd1882594, 32'sd3188861, 32'sd1719962, 32'sd2033945, -32'sd3255550, 32'sd550606, -32'sd1626160, 32'sd348557, -32'sd2387769, -32'sd1416587, -32'sd1714861, -32'sd1545128, -32'sd1200536, 32'sd1141667, 32'sd0, 32'sd732021, -32'sd892050, 32'sd139924, 32'sd1460195, 32'sd616831, -32'sd811936, -32'sd897510, 32'sd1082536, 32'sd80774, 32'sd738233, 32'sd453236, 32'sd1482465, 32'sd923257, 32'sd2869292, 32'sd2205484, -32'sd648754, -32'sd1683038, -32'sd365961, -32'sd836273, -32'sd946209, -32'sd1906938, -32'sd634880, 32'sd144706, -32'sd565207, -32'sd677056, 32'sd372959, 32'sd0, 32'sd0, 32'sd0, -32'sd1575472, 32'sd1764431, 32'sd987525, -32'sd1044249, -32'sd775779, 32'sd424868, -32'sd133617, -32'sd416615, 32'sd215026, 32'sd1245877, -32'sd649201, -32'sd467216, 32'sd277845, -32'sd391117, -32'sd3512883, -32'sd1481162, -32'sd2994194, -32'sd1026589, -32'sd590010, 32'sd526772, -32'sd1033499, 32'sd1522362, 32'sd696623, 32'sd548965, -32'sd689333, 32'sd0, 32'sd0, 32'sd0, 32'sd189800, 32'sd542556, -32'sd1024892, 32'sd559855, -32'sd1021872, -32'sd59640, -32'sd791244, 32'sd1471164, -32'sd2093847, -32'sd2664216, -32'sd918511, -32'sd1811390, 32'sd587409, 32'sd621658, -32'sd2238625, -32'sd1937450, -32'sd847276, 32'sd1487338, 32'sd96700, -32'sd768036, 32'sd1173858, 32'sd728742, 32'sd29682, -32'sd210177, 32'sd289578, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1527651, -32'sd746044, 32'sd334053, 32'sd355465, -32'sd318900, -32'sd897415, 32'sd502895, 32'sd1160416, -32'sd401024, 32'sd398740, 32'sd1386326, 32'sd176554, -32'sd767902, -32'sd1243496, 32'sd669407, 32'sd362859, -32'sd544767, 32'sd509031, 32'sd1400321, -32'sd220431, -32'sd479806, 32'sd1219118, 32'sd1082996, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1660488, 32'sd701012, -32'sd595181, 32'sd956501, 32'sd1628013, 32'sd232205, 32'sd1658153, 32'sd108169, 32'sd146611, 32'sd2224988, 32'sd3291922, 32'sd658280, 32'sd680751, -32'sd30340, -32'sd5666, -32'sd298261, 32'sd97604, -32'sd40291, -32'sd33154, 32'sd310253, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd823362, 32'sd1417012, -32'sd1199528, 32'sd252192, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd308443, 32'sd877466, -32'sd482647, -32'sd1529905, -32'sd1062724, 32'sd771804, -32'sd692122, 32'sd246329, 32'sd1752784, 32'sd148076, 32'sd1033382, -32'sd852719, -32'sd911988, 32'sd1350346, -32'sd158621, 32'sd1102925, 32'sd963132, 32'sd1006853, -32'sd853507, 32'sd768442, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1403296, 32'sd1177575, 32'sd757605, -32'sd256065, -32'sd337395, -32'sd1919080, 32'sd399614, -32'sd623106, -32'sd620990, -32'sd279284, 32'sd1509568, 32'sd2320546, 32'sd707001, 32'sd1006043, -32'sd254235, 32'sd164404, -32'sd2739641, -32'sd1079833, 32'sd77792, 32'sd3494, -32'sd175282, 32'sd1415066, 32'sd1825785, 32'sd1091627, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd104605, -32'sd91164, 32'sd634201, -32'sd1231604, -32'sd440436, 32'sd583064, -32'sd239490, 32'sd1010034, 32'sd816108, 32'sd693138, 32'sd780937, 32'sd409076, 32'sd572942, -32'sd753438, -32'sd1189641, -32'sd2857199, -32'sd3721391, -32'sd517889, 32'sd1048775, -32'sd1085181, -32'sd618855, 32'sd1544426, -32'sd595195, 32'sd1484134, 32'sd1867501, 32'sd0, 32'sd0, 32'sd728472, -32'sd114392, 32'sd763944, -32'sd204440, -32'sd612007, -32'sd1608716, 32'sd135395, 32'sd724168, 32'sd1695944, 32'sd1008204, -32'sd846036, 32'sd1309775, 32'sd1593016, -32'sd215877, -32'sd748364, -32'sd717142, -32'sd201091, -32'sd90412, 32'sd484374, 32'sd181035, 32'sd1008918, 32'sd99666, 32'sd1010099, -32'sd123640, 32'sd489013, -32'sd1017374, -32'sd788849, 32'sd0, 32'sd90531, -32'sd442118, 32'sd16803, 32'sd113568, -32'sd719270, -32'sd387604, 32'sd1186804, 32'sd1280427, 32'sd1765974, 32'sd1529716, -32'sd901293, -32'sd749464, -32'sd2392997, 32'sd490039, 32'sd26834, 32'sd912917, -32'sd673133, -32'sd2255200, -32'sd122678, -32'sd450828, -32'sd422587, 32'sd1047061, 32'sd1389654, 32'sd765689, 32'sd1391846, -32'sd483424, 32'sd1046252, 32'sd0, 32'sd18904, -32'sd529366, -32'sd951396, -32'sd1274864, 32'sd1371104, 32'sd596439, -32'sd249969, 32'sd1337112, -32'sd648147, 32'sd204334, -32'sd1472120, -32'sd2851851, -32'sd2245334, -32'sd1197927, 32'sd177044, -32'sd3051352, -32'sd1227376, -32'sd2035957, -32'sd3022626, 32'sd780190, -32'sd1459479, 32'sd1826299, 32'sd3060300, 32'sd2969043, 32'sd1316936, 32'sd1705820, 32'sd615714, 32'sd1268964, -32'sd292634, -32'sd489889, -32'sd141254, -32'sd1844029, 32'sd1259920, 32'sd542131, 32'sd1340907, 32'sd415141, 32'sd1113684, 32'sd533578, 32'sd324995, -32'sd2052568, -32'sd1177033, 32'sd423298, -32'sd420066, -32'sd2603483, 32'sd833607, -32'sd1927637, -32'sd317752, 32'sd336509, 32'sd1474229, -32'sd541198, -32'sd633555, 32'sd1293367, 32'sd980303, 32'sd397660, -32'sd108256, 32'sd583003, -32'sd1569193, -32'sd1332056, 32'sd135897, -32'sd1271447, -32'sd370100, 32'sd302429, 32'sd2884863, 32'sd1504157, 32'sd2979818, -32'sd672315, -32'sd1308309, 32'sd217957, -32'sd437969, -32'sd187116, 32'sd524634, -32'sd2322517, -32'sd1932975, -32'sd1176263, -32'sd616261, 32'sd1880606, 32'sd2611090, 32'sd1400681, -32'sd577267, -32'sd383050, 32'sd251324, 32'sd193173, 32'sd741757, 32'sd23790, -32'sd94128, -32'sd377395, -32'sd1716890, -32'sd397948, -32'sd831300, -32'sd1463950, 32'sd2839769, 32'sd751815, -32'sd777221, 32'sd126758, -32'sd991008, -32'sd2092005, -32'sd1516344, -32'sd1843459, 32'sd608882, -32'sd1142636, -32'sd2092985, -32'sd1215721, 32'sd1182507, 32'sd2635091, 32'sd2766922, 32'sd1016539, 32'sd712592, 32'sd545084, 32'sd376941, 32'sd983089, -32'sd146691, 32'sd440198, -32'sd855088, -32'sd1142353, 32'sd761993, -32'sd728156, -32'sd4332326, 32'sd399198, 32'sd873042, 32'sd2069346, 32'sd2796962, 32'sd2493281, -32'sd1014881, -32'sd259590, -32'sd24123, -32'sd1998741, -32'sd273503, -32'sd2017957, -32'sd2069817, -32'sd194057, 32'sd2397207, 32'sd1270291, -32'sd68911, 32'sd1384793, 32'sd3136887, 32'sd1036437, -32'sd1127977, -32'sd912992, -32'sd1122211, 32'sd53977, -32'sd467069, 32'sd1107562, -32'sd278325, -32'sd1540081, -32'sd2256991, -32'sd901118, -32'sd2042137, -32'sd343690, 32'sd1935414, 32'sd1529270, -32'sd1150745, -32'sd98030, 32'sd1204966, -32'sd302981, 32'sd425536, 32'sd18162, -32'sd2123387, -32'sd2075066, 32'sd1724638, 32'sd746787, 32'sd2520323, 32'sd754851, -32'sd606789, -32'sd539767, -32'sd1422986, -32'sd841985, -32'sd448946, 32'sd1103121, 32'sd729873, 32'sd434439, -32'sd125266, -32'sd876140, -32'sd2557104, 32'sd276724, 32'sd1758135, 32'sd1726167, 32'sd1396018, 32'sd61985, -32'sd1188844, -32'sd665888, 32'sd2751498, 32'sd1260896, 32'sd2028472, 32'sd447770, -32'sd1221898, 32'sd121274, -32'sd658665, 32'sd2143223, 32'sd42879, 32'sd698845, -32'sd14203, 32'sd781530, 32'sd201341, -32'sd1683890, 32'sd1199433, 32'sd250636, -32'sd373854, -32'sd10544, -32'sd2054660, -32'sd1977626, -32'sd1930240, 32'sd827532, 32'sd332463, -32'sd585088, 32'sd1240486, 32'sd432146, -32'sd564318, -32'sd804120, 32'sd225815, 32'sd1290239, 32'sd2928645, -32'sd1849587, -32'sd1724399, 32'sd103863, -32'sd206331, 32'sd314463, -32'sd115304, 32'sd776034, 32'sd1783694, -32'sd715719, -32'sd393032, -32'sd756426, -32'sd86509, 32'sd52019, 32'sd332582, 32'sd893484, -32'sd1520193, -32'sd1010493, -32'sd1043667, -32'sd1612879, 32'sd955670, 32'sd90296, -32'sd717781, -32'sd2961813, -32'sd2554943, -32'sd648143, 32'sd298563, 32'sd1706925, 32'sd2565845, 32'sd734530, -32'sd463175, 32'sd231431, 32'sd1132631, -32'sd3194854, -32'sd2088194, 32'sd484639, 32'sd558334, -32'sd495720, -32'sd2325820, -32'sd301298, 32'sd122389, -32'sd1244607, 32'sd541172, -32'sd573483, -32'sd716613, -32'sd498689, -32'sd405314, -32'sd954749, 32'sd173643, -32'sd525244, -32'sd1158625, -32'sd799323, -32'sd2179981, -32'sd1146450, -32'sd182078, 32'sd1212607, 32'sd1675519, -32'sd376056, 32'sd1203438, -32'sd153682, -32'sd2847383, -32'sd1296266, -32'sd2718382, 32'sd687514, -32'sd512081, -32'sd2007032, 32'sd690761, -32'sd1341298, 32'sd305609, 32'sd937957, -32'sd376789, -32'sd1183550, -32'sd581602, -32'sd374216, 32'sd495782, -32'sd1807551, -32'sd1619386, 32'sd91434, -32'sd786497, -32'sd2593099, 32'sd247174, -32'sd558475, 32'sd1571371, -32'sd532363, -32'sd630531, 32'sd1141745, -32'sd1112676, 32'sd194643, -32'sd885566, -32'sd3222798, -32'sd1761433, -32'sd637687, 32'sd6946, 32'sd342808, 32'sd1745791, 32'sd420382, 32'sd756437, 32'sd0, -32'sd1279059, 32'sd394837, -32'sd260908, -32'sd20421, -32'sd142662, 32'sd124595, -32'sd715756, -32'sd1646544, -32'sd1297293, -32'sd790148, 32'sd1683336, 32'sd2792202, 32'sd1704075, 32'sd1079829, 32'sd817330, 32'sd1503486, 32'sd654267, 32'sd805146, 32'sd716076, -32'sd556468, -32'sd148411, -32'sd768555, -32'sd291691, -32'sd271263, 32'sd209864, -32'sd1132098, -32'sd840600, -32'sd239186, 32'sd1311439, -32'sd525072, -32'sd40883, -32'sd685559, -32'sd668543, -32'sd6627, -32'sd1372326, -32'sd1847287, -32'sd2945132, -32'sd882320, 32'sd917955, 32'sd3886286, 32'sd4082053, 32'sd1392347, 32'sd1508035, 32'sd1259054, 32'sd462784, 32'sd2025510, -32'sd1325166, -32'sd370820, -32'sd1249453, -32'sd1472172, -32'sd469364, 32'sd58657, 32'sd484296, -32'sd1233420, -32'sd721749, 32'sd1425250, -32'sd1012073, -32'sd473462, 32'sd424065, -32'sd67071, -32'sd889691, -32'sd2399576, -32'sd1566643, -32'sd1387246, -32'sd682590, -32'sd596107, 32'sd2491010, 32'sd1670975, 32'sd1812535, 32'sd931677, -32'sd53040, 32'sd95952, -32'sd337737, 32'sd1120315, 32'sd5401, -32'sd1146977, -32'sd1185486, -32'sd184197, -32'sd1092007, -32'sd92296, -32'sd554606, -32'sd1586821, 32'sd999712, 32'sd0, -32'sd1429946, 32'sd793397, -32'sd71007, -32'sd2313974, -32'sd2326063, -32'sd572900, -32'sd2452332, -32'sd2574969, -32'sd1397666, -32'sd383332, 32'sd2721811, 32'sd3131102, 32'sd197868, 32'sd147320, 32'sd1358520, 32'sd1879674, 32'sd1240371, -32'sd14438, 32'sd466383, 32'sd1427823, 32'sd385841, -32'sd2357965, -32'sd1233731, 32'sd900943, 32'sd1012627, 32'sd680434, 32'sd482549, 32'sd20585, 32'sd784541, 32'sd124200, 32'sd538494, -32'sd1308706, -32'sd1584220, 32'sd320628, -32'sd2100288, -32'sd1282487, 32'sd326301, 32'sd618414, -32'sd442766, 32'sd175680, -32'sd48073, -32'sd251871, -32'sd370712, 32'sd1033617, 32'sd534325, -32'sd425750, -32'sd159246, -32'sd1024664, 32'sd325266, -32'sd225015, 32'sd1513297, 32'sd220865, -32'sd56171, -32'sd696845, -32'sd431074, 32'sd1316382, 32'sd1485445, 32'sd196671, -32'sd421947, -32'sd189179, -32'sd306380, -32'sd2770001, -32'sd1617450, -32'sd1845678, 32'sd1534107, 32'sd73218, 32'sd541211, 32'sd1325551, 32'sd1043525, 32'sd563755, -32'sd275618, 32'sd230238, -32'sd830653, -32'sd170738, 32'sd844834, -32'sd103360, -32'sd455565, -32'sd325693, 32'sd56558, -32'sd505859, 32'sd2036901, -32'sd632681, 32'sd882463, 32'sd0, 32'sd468489, -32'sd1246559, -32'sd131672, 32'sd1194127, -32'sd52518, -32'sd1974092, -32'sd2523992, 32'sd1152625, 32'sd1666806, 32'sd1004263, -32'sd297168, 32'sd1523017, 32'sd8699, 32'sd2924855, 32'sd463022, 32'sd1052039, 32'sd270603, 32'sd201502, 32'sd181760, -32'sd159714, 32'sd634195, -32'sd800446, -32'sd896553, 32'sd576147, 32'sd1372465, 32'sd1090400, 32'sd0, 32'sd0, 32'sd0, -32'sd1259795, 32'sd695655, -32'sd268763, -32'sd1448648, -32'sd981984, -32'sd2732163, -32'sd3135743, -32'sd917378, -32'sd899875, 32'sd2071545, 32'sd250444, -32'sd211581, 32'sd1585192, -32'sd290034, -32'sd1099943, -32'sd918690, -32'sd612107, -32'sd1073525, -32'sd1618525, 32'sd931429, 32'sd2618800, 32'sd627097, 32'sd423281, 32'sd853814, 32'sd362174, 32'sd0, 32'sd0, 32'sd0, 32'sd844827, 32'sd1049375, -32'sd1134819, 32'sd607962, 32'sd120244, -32'sd719715, -32'sd2043339, -32'sd1238417, -32'sd1538419, -32'sd1061217, -32'sd2565799, -32'sd459375, -32'sd634552, -32'sd176368, -32'sd526245, -32'sd1488823, 32'sd524471, 32'sd549194, 32'sd1385612, 32'sd682393, 32'sd321494, 32'sd213633, -32'sd1737638, 32'sd292081, 32'sd851338, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1179822, -32'sd272336, 32'sd2106114, 32'sd1751011, 32'sd767850, -32'sd611761, -32'sd845449, -32'sd499368, -32'sd1059222, 32'sd378101, -32'sd206557, -32'sd1574342, -32'sd1218269, 32'sd1259044, -32'sd66661, -32'sd370788, -32'sd311210, -32'sd51401, -32'sd338187, 32'sd302236, 32'sd119539, 32'sd425751, 32'sd171195, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1446829, 32'sd458173, 32'sd351954, 32'sd1026532, -32'sd407385, 32'sd272127, -32'sd612201, 32'sd424510, -32'sd651023, 32'sd268311, -32'sd478590, -32'sd1568335, 32'sd90496, 32'sd992314, -32'sd727283, -32'sd651486, 32'sd1801116, 32'sd157797, 32'sd99929, -32'sd987612, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd620447, -32'sd697930, -32'sd102559, -32'sd630524, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd440729, -32'sd854932, -32'sd281264, -32'sd861847, 32'sd21721, 32'sd156931, 32'sd991377, -32'sd263363, 32'sd555440, -32'sd687552, -32'sd1187410, -32'sd1342976, 32'sd742513, 32'sd1491830, 32'sd982551, -32'sd696895, 32'sd376055, -32'sd1268384, 32'sd92934, -32'sd268650, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd190897, -32'sd680311, 32'sd169932, 32'sd1208674, -32'sd1011377, 32'sd895488, 32'sd617077, 32'sd567877, -32'sd599943, -32'sd619352, -32'sd889634, 32'sd201346, -32'sd1079621, 32'sd505354, -32'sd2540572, 32'sd305446, 32'sd1506726, -32'sd612006, -32'sd48932, -32'sd816486, 32'sd240362, -32'sd1448261, -32'sd846529, -32'sd762499, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd124258, -32'sd1061652, 32'sd617235, 32'sd329451, 32'sd557948, 32'sd852181, 32'sd911966, -32'sd44288, -32'sd1902618, -32'sd407158, 32'sd994544, -32'sd652069, -32'sd389447, -32'sd385145, 32'sd1356375, 32'sd321487, 32'sd1129823, -32'sd1927985, -32'sd678311, 32'sd678865, -32'sd304009, 32'sd671701, 32'sd483226, -32'sd144576, 32'sd734881, 32'sd0, 32'sd0, 32'sd790024, -32'sd749800, 32'sd415677, 32'sd1586953, -32'sd418739, -32'sd276533, -32'sd1497047, -32'sd1362764, -32'sd3034658, -32'sd3853722, -32'sd251811, 32'sd1473475, 32'sd777343, 32'sd920578, 32'sd697394, -32'sd294885, -32'sd9158, 32'sd382693, -32'sd150622, 32'sd424713, 32'sd2478912, 32'sd24423, 32'sd1862330, 32'sd1368766, 32'sd1829429, -32'sd956238, 32'sd206973, 32'sd0, -32'sd921307, -32'sd38445, 32'sd816593, 32'sd212014, -32'sd1675949, -32'sd933519, -32'sd140367, -32'sd2056375, -32'sd1213899, 32'sd662240, 32'sd1752117, 32'sd2180933, 32'sd1649153, 32'sd1794720, 32'sd1077469, 32'sd1106648, 32'sd573026, 32'sd121950, 32'sd597080, 32'sd219432, -32'sd355228, 32'sd269680, 32'sd295803, 32'sd307471, 32'sd186349, -32'sd134263, -32'sd888806, 32'sd0, -32'sd659483, -32'sd1354774, -32'sd832256, -32'sd374974, -32'sd1022839, -32'sd1978545, -32'sd1121929, 32'sd491608, -32'sd1927054, 32'sd909251, 32'sd1115730, -32'sd69819, 32'sd1173855, 32'sd365456, -32'sd963990, -32'sd357285, -32'sd181149, -32'sd1378543, -32'sd1113692, -32'sd1008899, -32'sd902155, 32'sd2653041, 32'sd3170444, 32'sd983829, -32'sd2838670, -32'sd1459101, 32'sd164960, 32'sd12890, 32'sd450320, -32'sd1669259, -32'sd419509, -32'sd815758, 32'sd1032845, 32'sd46431, -32'sd2241994, 32'sd486574, 32'sd622394, -32'sd506213, 32'sd1021271, 32'sd21792, -32'sd415575, -32'sd605886, 32'sd338094, 32'sd1262479, -32'sd224851, 32'sd444438, -32'sd599575, -32'sd618775, -32'sd1083832, -32'sd1265157, -32'sd186828, -32'sd56589, -32'sd1884796, -32'sd1241032, -32'sd405827, 32'sd888433, -32'sd214507, 32'sd1174029, -32'sd726574, -32'sd650944, 32'sd346167, -32'sd1187992, -32'sd256395, -32'sd554692, -32'sd840062, -32'sd1040189, -32'sd142980, 32'sd189135, 32'sd1425807, -32'sd1241157, -32'sd1305206, 32'sd88167, -32'sd1021572, 32'sd556561, -32'sd1332471, 32'sd1039652, 32'sd393303, 32'sd132226, -32'sd749422, 32'sd257090, -32'sd829036, -32'sd741596, 32'sd944389, 32'sd373678, 32'sd736791, -32'sd893476, -32'sd723210, -32'sd2054139, -32'sd759696, -32'sd2841458, -32'sd559817, -32'sd683821, -32'sd942032, -32'sd93673, 32'sd79608, 32'sd199671, 32'sd1573419, -32'sd1397088, -32'sd2128008, -32'sd2589817, 32'sd216421, 32'sd1706341, 32'sd1275874, -32'sd254324, 32'sd1574957, 32'sd554971, 32'sd690517, 32'sd2066036, 32'sd2404506, 32'sd1683531, 32'sd504473, -32'sd975739, 32'sd192568, -32'sd497149, -32'sd355280, -32'sd2669361, -32'sd1785389, -32'sd711143, -32'sd2094508, -32'sd2556704, -32'sd726463, 32'sd368364, 32'sd1745750, 32'sd2818857, 32'sd1600545, 32'sd49854, -32'sd2272271, -32'sd980290, 32'sd102718, 32'sd2186937, 32'sd378723, -32'sd1253683, 32'sd1088369, 32'sd1719064, -32'sd330847, 32'sd218649, -32'sd296227, 32'sd1057735, 32'sd575785, 32'sd607880, -32'sd594376, -32'sd1082515, 32'sd838495, -32'sd1631805, -32'sd596822, -32'sd1473237, -32'sd1414360, -32'sd1467092, -32'sd190408, 32'sd1147695, 32'sd1029012, -32'sd164117, 32'sd446609, 32'sd1673343, -32'sd489138, 32'sd1704945, 32'sd3215933, 32'sd2894774, 32'sd653403, -32'sd774843, 32'sd238308, 32'sd112838, 32'sd2204695, 32'sd2312353, -32'sd500613, -32'sd1350312, -32'sd243874, -32'sd233637, -32'sd271460, -32'sd1096633, 32'sd300717, -32'sd402985, 32'sd1595468, 32'sd55193, -32'sd363874, 32'sd34477, 32'sd729476, -32'sd1468292, -32'sd725111, 32'sd347698, 32'sd1808037, 32'sd2330885, 32'sd1059548, 32'sd914059, 32'sd216610, 32'sd588663, 32'sd1504568, 32'sd1294779, 32'sd735246, 32'sd639416, -32'sd37559, 32'sd656003, -32'sd2666587, -32'sd1156327, -32'sd1429756, -32'sd425850, -32'sd529198, 32'sd1094143, -32'sd817924, 32'sd1602982, 32'sd625429, -32'sd692364, -32'sd1028691, -32'sd1894057, -32'sd1103527, -32'sd1364074, -32'sd265413, 32'sd1480894, 32'sd2420021, 32'sd2971292, 32'sd461124, -32'sd927680, -32'sd379079, 32'sd476017, 32'sd1378067, -32'sd511481, 32'sd66884, 32'sd29117, 32'sd771604, 32'sd1636179, -32'sd553260, 32'sd810425, 32'sd61834, -32'sd50148, -32'sd873024, -32'sd271044, 32'sd1711003, -32'sd232231, -32'sd654493, -32'sd2236343, -32'sd2410197, -32'sd1658749, -32'sd2529246, 32'sd1879, 32'sd38195, 32'sd1040330, 32'sd2388228, -32'sd575737, 32'sd143258, 32'sd682983, 32'sd271034, 32'sd1143541, 32'sd487351, 32'sd253841, -32'sd225052, -32'sd1134927, -32'sd1801316, -32'sd516434, -32'sd1041095, 32'sd647078, 32'sd145335, -32'sd578079, -32'sd699550, 32'sd936754, -32'sd87678, 32'sd90853, -32'sd584880, -32'sd48424, -32'sd1076819, -32'sd935798, -32'sd1049471, 32'sd360735, -32'sd474450, 32'sd1032569, -32'sd729953, -32'sd348138, 32'sd1848152, 32'sd480544, 32'sd1355375, 32'sd1479977, -32'sd202850, 32'sd220275, -32'sd2223141, -32'sd1860800, -32'sd2053086, -32'sd1687995, -32'sd739813, -32'sd1087254, 32'sd293403, -32'sd488831, -32'sd443449, 32'sd293230, 32'sd631681, 32'sd1621325, 32'sd1515256, -32'sd1394294, -32'sd1066286, -32'sd672042, -32'sd3136762, -32'sd2400623, -32'sd2340838, 32'sd986419, -32'sd1557146, 32'sd498939, -32'sd723574, -32'sd187496, 32'sd2033313, 32'sd1008631, 32'sd203606, -32'sd1112205, -32'sd3077154, -32'sd225600, -32'sd1265695, -32'sd1342610, 32'sd525554, -32'sd257313, -32'sd98953, 32'sd0, -32'sd825420, -32'sd480593, 32'sd273200, 32'sd142227, -32'sd207104, -32'sd249547, -32'sd2811495, -32'sd3052074, -32'sd3006369, -32'sd4388641, -32'sd1916155, 32'sd1906104, 32'sd397946, -32'sd1920911, 32'sd229807, 32'sd862267, 32'sd2745696, 32'sd1703972, 32'sd985600, 32'sd344803, 32'sd591187, -32'sd2457301, -32'sd775300, -32'sd2170213, 32'sd942509, -32'sd1295158, -32'sd1117517, 32'sd408075, -32'sd974575, 32'sd753595, -32'sd1242452, 32'sd2251996, 32'sd1101176, 32'sd1055998, -32'sd272650, -32'sd142546, -32'sd506469, 32'sd184259, 32'sd1429100, 32'sd1584833, -32'sd365783, -32'sd2156464, -32'sd839413, 32'sd398031, 32'sd2474281, 32'sd1860348, -32'sd662239, 32'sd36824, -32'sd2069442, -32'sd733078, -32'sd1537356, 32'sd126299, -32'sd807228, 32'sd1348413, -32'sd1416567, 32'sd77237, -32'sd669607, -32'sd663155, 32'sd716188, 32'sd681230, 32'sd414217, 32'sd1591610, -32'sd271607, 32'sd91008, 32'sd334657, 32'sd36030, -32'sd297943, -32'sd1409132, -32'sd1155087, -32'sd1006323, -32'sd957356, 32'sd94474, 32'sd1559298, 32'sd2264487, -32'sd1060587, -32'sd595616, -32'sd1123339, -32'sd2989755, -32'sd1259053, 32'sd161012, -32'sd8522, 32'sd1005141, -32'sd319959, 32'sd0, -32'sd849514, -32'sd1348281, -32'sd996718, -32'sd312417, 32'sd2319291, 32'sd642662, -32'sd123783, -32'sd361739, 32'sd139940, 32'sd751478, 32'sd354213, -32'sd395929, 32'sd401675, -32'sd739923, 32'sd396416, -32'sd97464, 32'sd2267453, -32'sd64938, -32'sd939514, -32'sd3697145, -32'sd1425347, -32'sd2218224, -32'sd490084, 32'sd588061, -32'sd446757, -32'sd1353808, -32'sd83481, -32'sd11710, -32'sd930941, 32'sd1387957, 32'sd1112149, 32'sd704722, -32'sd1036438, -32'sd162320, -32'sd991450, -32'sd1504722, -32'sd674942, 32'sd1574137, 32'sd1711086, -32'sd1565522, 32'sd219216, 32'sd1408092, 32'sd1164231, 32'sd939366, 32'sd1122895, -32'sd525186, -32'sd2680870, -32'sd2770049, -32'sd1958729, -32'sd3500185, -32'sd1332105, -32'sd1830595, 32'sd77848, 32'sd78592, -32'sd160301, -32'sd183985, -32'sd420648, 32'sd935086, -32'sd509178, 32'sd278692, -32'sd1460906, -32'sd793629, 32'sd1404403, 32'sd107265, 32'sd481891, -32'sd378400, 32'sd174505, 32'sd2110620, 32'sd114690, 32'sd1236040, 32'sd1723611, -32'sd525267, -32'sd484132, -32'sd1437404, -32'sd2631435, -32'sd1902479, -32'sd3977626, -32'sd1608910, -32'sd56506, -32'sd583659, -32'sd67924, 32'sd1006626, 32'sd255417, 32'sd0, -32'sd349675, -32'sd539317, -32'sd247457, 32'sd724331, 32'sd395572, -32'sd1396002, 32'sd1182956, -32'sd534652, 32'sd293673, 32'sd490753, 32'sd1401384, 32'sd1155297, 32'sd432610, 32'sd1346363, -32'sd171954, -32'sd1005969, -32'sd1222299, -32'sd922035, -32'sd2167758, -32'sd527129, -32'sd2299671, -32'sd818710, -32'sd930517, -32'sd562827, 32'sd595261, -32'sd1877620, 32'sd0, 32'sd0, 32'sd0, 32'sd76607, 32'sd1726303, -32'sd796688, -32'sd2213937, -32'sd1847884, 32'sd1248035, -32'sd1362201, -32'sd1455037, 32'sd881930, 32'sd1063021, 32'sd625536, 32'sd2518427, 32'sd1839847, 32'sd1688246, -32'sd976241, -32'sd2052451, -32'sd3378349, -32'sd3137436, 32'sd952013, -32'sd1422142, -32'sd990476, 32'sd354803, -32'sd37706, 32'sd641006, -32'sd876682, 32'sd0, 32'sd0, 32'sd0, -32'sd914871, 32'sd782632, -32'sd1142171, -32'sd1398092, 32'sd57403, 32'sd566269, -32'sd1208793, 32'sd1032284, -32'sd36195, 32'sd403756, -32'sd931783, 32'sd1053435, 32'sd457745, 32'sd1876067, -32'sd1008938, -32'sd2805398, -32'sd1926438, 32'sd84141, -32'sd569932, -32'sd549943, -32'sd400908, -32'sd707673, -32'sd757465, 32'sd325392, 32'sd1348950, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd706863, 32'sd1406667, -32'sd169715, -32'sd1063271, 32'sd635224, 32'sd880801, 32'sd237869, -32'sd1533240, 32'sd74370, -32'sd110632, -32'sd1289644, -32'sd3466233, -32'sd1004804, 32'sd4525, -32'sd750585, -32'sd286396, -32'sd1038422, -32'sd852401, -32'sd179525, 32'sd233762, -32'sd1071690, -32'sd669005, -32'sd623035, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd71660, 32'sd140902, 32'sd452364, 32'sd1378119, 32'sd456149, 32'sd813525, -32'sd468998, -32'sd1359409, 32'sd432419, -32'sd1866979, 32'sd728912, -32'sd705762, -32'sd1481760, 32'sd80103, 32'sd740592, -32'sd51732, -32'sd701729, -32'sd697726, 32'sd668836, 32'sd410926, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd260765, 32'sd1673255, 32'sd1339869, 32'sd631536, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd698599, 32'sd1498705, 32'sd87375, 32'sd473265, 32'sd2045493, -32'sd57897, 32'sd574822, -32'sd279729, 32'sd835900, 32'sd279138, 32'sd693043, 32'sd1465603, 32'sd1758708, -32'sd1182283, -32'sd1738864, 32'sd1152964, 32'sd903715, -32'sd557320, 32'sd760610, 32'sd872750, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd331985, 32'sd632830, 32'sd792179, -32'sd884891, 32'sd1560703, 32'sd1674565, 32'sd818492, 32'sd412928, 32'sd310429, -32'sd1679872, -32'sd1740585, -32'sd84249, 32'sd186066, -32'sd1012689, 32'sd1610025, 32'sd349668, 32'sd705650, 32'sd43598, 32'sd1967317, 32'sd727254, -32'sd805958, -32'sd137803, 32'sd827556, 32'sd1062170, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1431939, 32'sd963997, 32'sd100923, -32'sd594376, -32'sd202788, -32'sd1034198, -32'sd739987, -32'sd1222166, -32'sd948925, -32'sd2393518, -32'sd2825503, 32'sd641092, -32'sd1695537, -32'sd1887649, -32'sd513239, -32'sd617311, -32'sd1930573, -32'sd1299000, 32'sd935244, 32'sd2050882, -32'sd1181929, -32'sd570361, 32'sd487056, 32'sd883332, -32'sd407908, 32'sd0, 32'sd0, 32'sd475852, -32'sd147741, 32'sd1135759, -32'sd1485999, -32'sd1834764, -32'sd706283, 32'sd155279, -32'sd666621, -32'sd1356260, -32'sd1214590, -32'sd884406, -32'sd48338, 32'sd492307, 32'sd1146279, 32'sd1343471, -32'sd322030, 32'sd1501065, 32'sd568103, -32'sd2616114, -32'sd259503, -32'sd281432, -32'sd760558, -32'sd644309, -32'sd976825, 32'sd88254, -32'sd792525, 32'sd286329, 32'sd0, 32'sd670694, 32'sd883407, 32'sd195875, -32'sd1184102, -32'sd1076413, -32'sd792439, -32'sd225716, -32'sd60624, -32'sd483025, 32'sd1421231, -32'sd1265433, -32'sd837112, 32'sd1597348, 32'sd130722, -32'sd1594475, 32'sd1072860, 32'sd126597, -32'sd1666535, -32'sd768218, -32'sd811685, -32'sd834288, -32'sd1796858, -32'sd1391400, -32'sd1109417, -32'sd261825, 32'sd1576207, -32'sd368427, 32'sd0, -32'sd434970, 32'sd403674, -32'sd191417, 32'sd924208, 32'sd1314461, -32'sd955945, -32'sd407015, 32'sd2841, 32'sd1954423, -32'sd1205435, -32'sd791592, 32'sd864040, 32'sd2677469, 32'sd747338, 32'sd1115444, 32'sd262163, 32'sd1341190, 32'sd1833456, -32'sd625269, -32'sd578637, 32'sd664217, -32'sd2358055, -32'sd1947911, -32'sd2966873, -32'sd1766745, -32'sd1396232, -32'sd35279, -32'sd40128, 32'sd353471, -32'sd577317, 32'sd195840, 32'sd167233, 32'sd142268, 32'sd836620, 32'sd298258, 32'sd1005450, 32'sd582375, -32'sd767931, 32'sd136447, -32'sd569139, 32'sd787896, 32'sd1348486, 32'sd2685257, 32'sd752792, 32'sd632672, 32'sd1669295, 32'sd235765, -32'sd1535474, -32'sd291569, -32'sd1314491, -32'sd1800094, -32'sd747605, 32'sd859018, -32'sd709634, -32'sd297701, 32'sd117718, -32'sd303810, 32'sd585304, 32'sd65304, 32'sd534045, -32'sd368088, 32'sd627198, 32'sd578598, 32'sd1220221, 32'sd1907250, 32'sd2260110, -32'sd144950, 32'sd1119696, 32'sd372983, 32'sd1296093, 32'sd2134586, -32'sd200051, -32'sd1474668, 32'sd2083272, 32'sd2808962, 32'sd1499714, 32'sd347270, -32'sd1024828, -32'sd2302036, -32'sd429345, -32'sd1038617, -32'sd42782, -32'sd478358, 32'sd1265789, -32'sd24087, 32'sd476880, 32'sd108166, -32'sd367503, 32'sd944888, -32'sd151618, 32'sd1895650, 32'sd668368, -32'sd1110514, 32'sd1911822, 32'sd1807428, -32'sd166547, -32'sd1331414, -32'sd408305, -32'sd1420786, -32'sd806516, 32'sd1186518, -32'sd451994, 32'sd2523455, 32'sd1306222, -32'sd1486459, -32'sd942082, -32'sd1534670, 32'sd853246, -32'sd1493673, -32'sd2092806, -32'sd355330, -32'sd625410, 32'sd759852, 32'sd358580, -32'sd2677215, -32'sd1132831, 32'sd593672, 32'sd1862327, 32'sd1367311, 32'sd380401, -32'sd539206, 32'sd140008, 32'sd1601872, -32'sd2193445, 32'sd857140, -32'sd3248705, -32'sd2501192, 32'sd1271022, -32'sd844228, 32'sd2020333, 32'sd2310393, 32'sd2402389, -32'sd1376227, -32'sd1194059, -32'sd1900887, -32'sd1975525, -32'sd707173, -32'sd390563, 32'sd465692, 32'sd659887, 32'sd415517, -32'sd1160314, 32'sd1013573, 32'sd895767, 32'sd766555, 32'sd1065504, 32'sd365092, 32'sd495867, -32'sd780276, -32'sd970757, 32'sd1304591, 32'sd436576, -32'sd2309560, -32'sd3363015, 32'sd604238, -32'sd214949, 32'sd774912, 32'sd2250746, 32'sd1186457, 32'sd2319671, 32'sd389397, 32'sd946581, -32'sd1406455, 32'sd301455, 32'sd1610299, 32'sd862584, 32'sd682426, -32'sd586025, 32'sd1077702, 32'sd1250564, -32'sd144235, -32'sd25418, -32'sd1799268, -32'sd175415, -32'sd784720, 32'sd627526, -32'sd48292, 32'sd5039, -32'sd748103, 32'sd1449023, -32'sd3291522, -32'sd3263819, -32'sd2112977, 32'sd64554, 32'sd1464693, 32'sd2590687, 32'sd2968741, 32'sd1818984, -32'sd219329, -32'sd445979, -32'sd163341, -32'sd1635960, 32'sd120001, 32'sd426622, -32'sd980875, 32'sd280601, 32'sd2584, 32'sd1432645, 32'sd192629, 32'sd11540, -32'sd43886, 32'sd558338, -32'sd652297, 32'sd929818, -32'sd519671, 32'sd805234, -32'sd745448, -32'sd498966, -32'sd2059536, -32'sd3759119, -32'sd446218, -32'sd1154237, 32'sd683834, 32'sd2388526, 32'sd1852808, 32'sd977236, 32'sd202952, -32'sd134075, -32'sd383839, -32'sd1360779, 32'sd984081, 32'sd12524, 32'sd1007092, -32'sd124403, 32'sd628715, 32'sd1281169, -32'sd1238697, -32'sd649477, -32'sd603371, 32'sd315217, -32'sd1345875, -32'sd1225452, -32'sd1771602, 32'sd958942, 32'sd462228, -32'sd303396, -32'sd1595922, -32'sd2924216, -32'sd1475134, 32'sd444173, 32'sd1469210, 32'sd1763386, 32'sd3154736, -32'sd230163, -32'sd807676, 32'sd448872, 32'sd2230991, -32'sd1555491, 32'sd578799, -32'sd526932, 32'sd605070, 32'sd211588, -32'sd2058673, -32'sd844049, -32'sd2010600, -32'sd965948, -32'sd2771093, -32'sd142904, 32'sd383369, -32'sd148481, 32'sd217658, 32'sd708185, -32'sd1853142, -32'sd4469702, -32'sd3842922, -32'sd1305645, -32'sd680167, 32'sd1039893, -32'sd466494, 32'sd1818608, 32'sd2030038, -32'sd1114569, -32'sd882819, 32'sd435102, -32'sd274162, -32'sd1244545, -32'sd91881, -32'sd322268, 32'sd1013955, 32'sd629856, 32'sd668294, 32'sd260184, -32'sd987497, -32'sd93275, -32'sd1787097, 32'sd412408, 32'sd993105, -32'sd1289849, -32'sd1567977, -32'sd823318, -32'sd1363145, -32'sd4761173, -32'sd1453909, 32'sd858053, 32'sd1912390, 32'sd198263, 32'sd968349, -32'sd931466, 32'sd570934, 32'sd655110, 32'sd352562, -32'sd537463, 32'sd2360094, 32'sd239264, -32'sd48474, -32'sd1676000, -32'sd1256059, 32'sd0, 32'sd28890, -32'sd913464, -32'sd1164801, -32'sd553265, -32'sd1196983, -32'sd1026618, -32'sd98981, -32'sd920719, -32'sd146033, -32'sd3259943, -32'sd3865304, -32'sd2964309, 32'sd687768, 32'sd1384507, 32'sd1210673, 32'sd2121090, 32'sd714170, 32'sd2031995, -32'sd1599744, -32'sd415671, -32'sd2578986, -32'sd1217344, -32'sd673498, -32'sd1626586, -32'sd1646309, -32'sd855547, 32'sd737163, 32'sd228405, 32'sd1543408, 32'sd844416, -32'sd685667, -32'sd2274329, -32'sd1697592, -32'sd967360, -32'sd602484, -32'sd1136975, -32'sd2277541, -32'sd3331947, -32'sd3437295, -32'sd628646, 32'sd1733426, 32'sd531125, 32'sd76104, 32'sd1356714, -32'sd652672, -32'sd61163, -32'sd398212, -32'sd1351230, -32'sd3631139, -32'sd539164, 32'sd784292, 32'sd1441710, 32'sd831898, 32'sd1288162, 32'sd901653, 32'sd27968, -32'sd613844, -32'sd976357, 32'sd358675, -32'sd1387451, -32'sd430931, -32'sd783300, 32'sd1766369, -32'sd884569, -32'sd1846985, -32'sd791254, -32'sd1603902, 32'sd2950282, 32'sd2541338, 32'sd2559326, 32'sd474917, 32'sd1151715, 32'sd1374504, -32'sd485233, -32'sd375561, -32'sd1862240, -32'sd2202758, -32'sd2348573, -32'sd718878, 32'sd1244339, -32'sd317274, 32'sd1311139, 32'sd337669, 32'sd0, 32'sd422300, 32'sd41863, 32'sd855398, -32'sd446454, -32'sd1233637, 32'sd42392, 32'sd872987, 32'sd1392641, -32'sd1049637, -32'sd1280140, 32'sd24017, 32'sd2990714, 32'sd1857343, 32'sd1324873, 32'sd873995, 32'sd1054674, -32'sd1606519, 32'sd305043, 32'sd259105, -32'sd1423545, 32'sd623514, -32'sd2248110, 32'sd768403, 32'sd2243370, -32'sd186701, 32'sd142484, -32'sd41860, -32'sd202834, 32'sd1168203, 32'sd883501, -32'sd456575, -32'sd1287648, -32'sd1000787, -32'sd1517604, -32'sd1583360, 32'sd67755, 32'sd149555, -32'sd864264, -32'sd1774929, 32'sd1760358, 32'sd1424286, -32'sd144341, 32'sd1036009, -32'sd935358, -32'sd277007, 32'sd1307768, 32'sd554751, -32'sd729762, 32'sd865917, 32'sd1248623, 32'sd1068490, 32'sd1916749, -32'sd1083654, -32'sd787392, -32'sd614609, -32'sd553984, -32'sd561178, 32'sd475060, -32'sd1186487, -32'sd1855893, -32'sd2150788, -32'sd9209, -32'sd1144953, 32'sd2286432, -32'sd398816, -32'sd2311736, -32'sd1770563, -32'sd557138, 32'sd358316, 32'sd1602680, 32'sd1127610, 32'sd1306413, 32'sd1825245, 32'sd457366, -32'sd2419615, -32'sd353390, -32'sd1986594, 32'sd52026, -32'sd624947, 32'sd506114, -32'sd28051, -32'sd933850, 32'sd417291, 32'sd0, -32'sd718381, 32'sd335694, 32'sd39274, -32'sd1500371, -32'sd855511, -32'sd381180, -32'sd492667, -32'sd806620, 32'sd277319, -32'sd1991361, 32'sd449520, -32'sd172491, 32'sd339047, 32'sd727864, -32'sd472800, -32'sd550839, -32'sd719192, -32'sd1432192, 32'sd1540732, 32'sd144009, -32'sd182956, -32'sd537867, -32'sd563006, -32'sd1439751, 32'sd203588, -32'sd23954, 32'sd0, 32'sd0, 32'sd0, -32'sd117031, -32'sd1226272, -32'sd2032352, -32'sd3233415, -32'sd459632, -32'sd805553, -32'sd1156573, -32'sd431734, -32'sd922595, -32'sd773612, -32'sd2644595, 32'sd1298818, 32'sd434993, -32'sd299948, 32'sd579713, 32'sd107973, 32'sd630241, 32'sd968362, 32'sd364274, -32'sd1120411, 32'sd289027, -32'sd252514, 32'sd264480, 32'sd297654, 32'sd6563, 32'sd0, 32'sd0, 32'sd0, 32'sd618982, -32'sd103036, -32'sd1297010, -32'sd2010153, -32'sd37597, -32'sd1037043, -32'sd2002670, -32'sd1662130, -32'sd326609, 32'sd4408, 32'sd191815, -32'sd162467, 32'sd1930366, 32'sd145942, 32'sd181594, 32'sd985650, 32'sd893507, 32'sd768369, 32'sd1190027, 32'sd340710, -32'sd638453, 32'sd816348, -32'sd101382, 32'sd807521, 32'sd14942, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd569401, 32'sd616381, -32'sd871774, -32'sd2013013, -32'sd1322883, 32'sd1676193, 32'sd2165562, 32'sd1333814, 32'sd22378, -32'sd988741, 32'sd1220302, 32'sd2153856, -32'sd852462, 32'sd447833, 32'sd690119, 32'sd2044922, 32'sd1789970, 32'sd1798031, -32'sd247502, 32'sd33877, 32'sd271554, 32'sd408583, -32'sd59214, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1281726, 32'sd42137, -32'sd379423, 32'sd1476226, 32'sd990151, -32'sd864730, 32'sd999685, 32'sd1440200, -32'sd59714, 32'sd230256, -32'sd7658, 32'sd647315, 32'sd488678, 32'sd194575, 32'sd416857, -32'sd328243, -32'sd592556, 32'sd786166, 32'sd1606140, 32'sd1782519, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1575611, -32'sd1448044, -32'sd1268692, -32'sd998659, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd758079, -32'sd1338125, -32'sd144415, -32'sd2154247, -32'sd520514, 32'sd1158235, 32'sd729865, -32'sd1417329, -32'sd1355029, -32'sd825284, 32'sd324286, 32'sd1217789, -32'sd51103, 32'sd130450, 32'sd285498, -32'sd192867, -32'sd2450962, -32'sd1970494, 32'sd188343, 32'sd698607, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd574587, -32'sd970312, 32'sd32218, 32'sd919946, -32'sd2299826, 32'sd960277, 32'sd988805, 32'sd2076709, 32'sd1771393, -32'sd981809, -32'sd481845, -32'sd743847, 32'sd478943, 32'sd670624, -32'sd1901890, -32'sd1338844, 32'sd540700, -32'sd701846, -32'sd1171400, 32'sd322694, -32'sd932470, -32'sd1493364, -32'sd1116221, -32'sd1464762, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd655283, -32'sd841604, 32'sd12728, -32'sd2467435, -32'sd4111956, -32'sd2517608, -32'sd831728, -32'sd190388, 32'sd797955, -32'sd676359, -32'sd295107, 32'sd557070, 32'sd478819, -32'sd554155, -32'sd79001, -32'sd798600, -32'sd357823, 32'sd509360, 32'sd773317, -32'sd15726, -32'sd1250996, 32'sd983391, -32'sd1541454, -32'sd1477071, -32'sd912148, 32'sd0, 32'sd0, 32'sd714083, 32'sd993927, -32'sd1856394, -32'sd221130, -32'sd1063087, -32'sd54787, -32'sd1211093, 32'sd1041894, 32'sd2253392, 32'sd2702373, 32'sd1387159, 32'sd78143, 32'sd544552, 32'sd2472121, 32'sd1662990, -32'sd1856177, -32'sd1172337, -32'sd991892, -32'sd343062, 32'sd2131171, 32'sd805342, 32'sd1130615, -32'sd296845, 32'sd151960, -32'sd392818, -32'sd835878, 32'sd971017, 32'sd0, -32'sd411541, 32'sd564722, 32'sd536881, 32'sd1638169, 32'sd754994, -32'sd1121390, 32'sd614627, 32'sd2020483, 32'sd1817460, 32'sd2546929, 32'sd1672385, 32'sd1496312, -32'sd482164, -32'sd663494, 32'sd204167, -32'sd155961, -32'sd2181594, -32'sd847404, -32'sd2409984, -32'sd402719, -32'sd788262, 32'sd143809, 32'sd1531459, 32'sd720669, -32'sd142787, -32'sd818939, -32'sd574743, 32'sd0, -32'sd1178089, 32'sd153423, 32'sd360706, -32'sd200792, -32'sd425691, 32'sd1738746, 32'sd1778147, 32'sd1109995, 32'sd1536808, 32'sd894285, 32'sd2943010, 32'sd1257601, 32'sd581458, -32'sd728838, -32'sd554884, -32'sd1331307, -32'sd205513, -32'sd2123932, 32'sd470494, -32'sd2031909, -32'sd1376198, -32'sd1409362, 32'sd623510, 32'sd1489667, -32'sd897764, -32'sd879866, 32'sd725867, -32'sd886163, 32'sd663305, 32'sd447255, -32'sd1257075, -32'sd10060, 32'sd1810904, -32'sd358696, 32'sd234187, -32'sd195555, 32'sd630471, 32'sd1407131, -32'sd87566, 32'sd687248, 32'sd2163292, 32'sd456716, -32'sd860654, -32'sd622763, 32'sd1251567, -32'sd169654, 32'sd175274, -32'sd151864, 32'sd2064943, 32'sd2354337, 32'sd502967, -32'sd1234102, 32'sd776420, 32'sd1504741, -32'sd482126, -32'sd629754, 32'sd104157, -32'sd1374274, -32'sd174324, -32'sd1210860, 32'sd394184, -32'sd124560, -32'sd383888, 32'sd1476654, 32'sd2874209, 32'sd1960542, 32'sd200057, -32'sd865801, -32'sd181220, 32'sd1731702, 32'sd883980, 32'sd162578, -32'sd711615, -32'sd940882, -32'sd29565, -32'sd956240, -32'sd163229, 32'sd248966, -32'sd710024, -32'sd1402427, 32'sd888852, 32'sd1163011, 32'sd1858031, -32'sd1947130, -32'sd404367, -32'sd859362, 32'sd539576, -32'sd857699, -32'sd99604, 32'sd711638, -32'sd593281, 32'sd2625722, 32'sd2587012, 32'sd1188138, -32'sd2368882, -32'sd5923177, -32'sd2960406, -32'sd309082, 32'sd38368, 32'sd743972, -32'sd628239, -32'sd272008, 32'sd2502239, -32'sd987598, -32'sd1565160, -32'sd1124174, 32'sd747438, 32'sd1681755, 32'sd533704, 32'sd1086338, 32'sd618718, -32'sd917775, -32'sd2103332, -32'sd2601273, 32'sd1470930, 32'sd105723, 32'sd1704922, 32'sd1947182, 32'sd1342605, 32'sd3562820, 32'sd3265964, 32'sd305279, -32'sd2757916, -32'sd3713804, -32'sd2823712, 32'sd1689938, -32'sd814376, -32'sd420315, 32'sd149864, 32'sd1859971, -32'sd255225, -32'sd137137, -32'sd832778, -32'sd1046420, 32'sd1535056, 32'sd2388452, -32'sd408478, -32'sd532846, 32'sd1018214, -32'sd1228880, -32'sd1475045, -32'sd248599, -32'sd768517, 32'sd768299, -32'sd227646, -32'sd561110, 32'sd1725586, 32'sd2308395, 32'sd2865687, 32'sd1337096, -32'sd220445, -32'sd1307762, -32'sd162396, -32'sd97175, -32'sd389202, -32'sd971299, -32'sd472823, -32'sd798396, 32'sd660796, -32'sd932561, -32'sd339459, -32'sd1943551, 32'sd171572, 32'sd1163269, -32'sd558803, 32'sd1640058, -32'sd1527263, -32'sd1227568, -32'sd826080, -32'sd2255555, 32'sd794060, -32'sd1183686, 32'sd613737, 32'sd3059700, 32'sd3069423, 32'sd1496320, 32'sd3411374, 32'sd101954, 32'sd1592694, 32'sd2023427, 32'sd1173754, -32'sd1535037, -32'sd1444159, -32'sd1280715, -32'sd1024952, -32'sd1501730, 32'sd66483, -32'sd823959, -32'sd94007, -32'sd2919297, -32'sd819156, 32'sd981617, -32'sd275979, -32'sd305584, -32'sd1344478, -32'sd916190, 32'sd211698, -32'sd1890959, 32'sd425626, -32'sd1203221, 32'sd821318, 32'sd1921720, 32'sd975850, 32'sd850454, 32'sd1767986, 32'sd2490736, 32'sd3664821, 32'sd288445, 32'sd1191767, 32'sd144285, 32'sd373622, -32'sd1789689, -32'sd812333, -32'sd62359, 32'sd2197787, -32'sd1112451, -32'sd822461, 32'sd981140, -32'sd1936720, -32'sd1783806, 32'sd317033, 32'sd975110, -32'sd1918961, 32'sd1052953, -32'sd880744, 32'sd147025, -32'sd1711384, -32'sd1084335, 32'sd2204276, 32'sd1582278, 32'sd568722, 32'sd243234, 32'sd1098718, 32'sd658387, 32'sd1087880, 32'sd29800, -32'sd1119312, -32'sd48006, -32'sd1081745, -32'sd1590473, 32'sd1785988, 32'sd1520866, -32'sd879259, -32'sd831221, 32'sd259117, -32'sd334463, -32'sd1073311, -32'sd657902, 32'sd1476455, 32'sd93652, -32'sd121667, 32'sd1282712, 32'sd186804, -32'sd1264222, -32'sd773620, -32'sd839281, 32'sd996284, 32'sd631187, -32'sd1015691, -32'sd1114142, 32'sd1948465, 32'sd2010206, 32'sd2686879, 32'sd937060, 32'sd1460868, 32'sd99134, -32'sd441325, 32'sd774720, -32'sd917496, 32'sd30787, 32'sd932654, 32'sd590215, -32'sd643035, 32'sd239162, -32'sd880734, 32'sd714991, 32'sd678734, -32'sd533619, 32'sd698212, 32'sd705563, 32'sd560567, -32'sd415225, -32'sd2685899, -32'sd26481, 32'sd409587, -32'sd2253416, -32'sd1397132, -32'sd1657986, -32'sd1723911, 32'sd1923049, 32'sd2643888, 32'sd1410176, 32'sd1224806, -32'sd1861394, -32'sd568874, 32'sd807177, -32'sd2162017, 32'sd1161543, 32'sd613259, 32'sd436184, -32'sd1132020, -32'sd1529902, 32'sd1674971, 32'sd504845, 32'sd163566, 32'sd1250335, 32'sd510372, 32'sd0, -32'sd55303, 32'sd27233, 32'sd835842, -32'sd721084, -32'sd557245, 32'sd8268, -32'sd3226510, -32'sd1454760, -32'sd534028, 32'sd2037323, 32'sd1332654, 32'sd144124, 32'sd984182, 32'sd1016051, -32'sd1036264, 32'sd783623, -32'sd3626743, -32'sd1530976, -32'sd153517, 32'sd1197218, -32'sd155305, 32'sd771042, -32'sd228032, 32'sd2039353, -32'sd174525, -32'sd1321780, -32'sd1326818, -32'sd1723036, 32'sd1417050, -32'sd67375, 32'sd905259, -32'sd1249139, -32'sd564394, 32'sd916603, -32'sd1463278, -32'sd1370565, 32'sd1256081, -32'sd286743, -32'sd295336, 32'sd107332, 32'sd537583, 32'sd1204350, -32'sd1432779, -32'sd2841251, -32'sd3524135, -32'sd2524388, -32'sd333670, 32'sd1387217, 32'sd388612, -32'sd1675223, -32'sd941657, 32'sd1980553, 32'sd613046, 32'sd329445, -32'sd1416412, -32'sd1470323, 32'sd757040, -32'sd335782, 32'sd2017264, -32'sd1393081, 32'sd238398, 32'sd1117438, -32'sd354972, 32'sd1768055, 32'sd2012638, -32'sd754043, -32'sd1616700, -32'sd319389, 32'sd2200002, 32'sd549135, 32'sd2305220, -32'sd2069979, -32'sd4111129, -32'sd2191790, -32'sd1527654, 32'sd1276469, 32'sd1493046, 32'sd1533857, -32'sd782327, 32'sd243574, -32'sd1146418, 32'sd346998, -32'sd1711139, 32'sd0, 32'sd1275547, -32'sd19852, 32'sd86918, 32'sd865314, -32'sd1329220, -32'sd595486, 32'sd45928, 32'sd1888403, 32'sd1333130, 32'sd719877, 32'sd905082, -32'sd678243, -32'sd250992, 32'sd1159179, 32'sd1254941, -32'sd827369, -32'sd1447150, -32'sd801752, -32'sd648376, 32'sd2645364, 32'sd215796, 32'sd687861, 32'sd1183622, -32'sd654818, -32'sd747357, 32'sd1203, -32'sd1343913, -32'sd1059181, -32'sd1558705, -32'sd783637, 32'sd1093875, -32'sd19137, -32'sd502789, 32'sd475247, 32'sd1773611, 32'sd1442967, 32'sd1574724, -32'sd840732, -32'sd1277021, -32'sd2571378, -32'sd991536, 32'sd257465, 32'sd4277015, 32'sd478702, 32'sd208757, -32'sd451124, 32'sd430222, 32'sd1660603, 32'sd2279869, 32'sd1039858, 32'sd465826, -32'sd936549, -32'sd534383, 32'sd576572, -32'sd469500, -32'sd1346458, 32'sd1021145, 32'sd453857, 32'sd328292, -32'sd592071, -32'sd2708939, -32'sd1921959, 32'sd1000117, 32'sd1244361, 32'sd768396, 32'sd2081323, 32'sd803304, -32'sd923754, -32'sd2065233, 32'sd327300, 32'sd631008, 32'sd764892, 32'sd274620, 32'sd1695062, 32'sd598189, 32'sd1494120, 32'sd867142, 32'sd656294, 32'sd1992021, -32'sd806207, 32'sd363190, -32'sd241718, -32'sd1086665, 32'sd0, -32'sd1381356, 32'sd1329114, -32'sd15001, 32'sd1753077, -32'sd367420, -32'sd646060, -32'sd14630, -32'sd67170, 32'sd393635, -32'sd411906, 32'sd131003, 32'sd86544, 32'sd1130519, -32'sd662185, -32'sd1265999, 32'sd1567612, 32'sd1394983, 32'sd1039313, 32'sd2781903, 32'sd209475, 32'sd679341, 32'sd982220, -32'sd463333, -32'sd1688423, -32'sd1374307, -32'sd1383824, 32'sd0, 32'sd0, 32'sd0, -32'sd212183, -32'sd1931888, -32'sd1701901, -32'sd1772108, -32'sd918928, 32'sd617214, -32'sd168648, 32'sd656785, -32'sd109635, 32'sd1320352, 32'sd624581, 32'sd1395292, -32'sd1807007, 32'sd200079, -32'sd96216, 32'sd295657, 32'sd1468923, 32'sd1656922, 32'sd929133, -32'sd210075, 32'sd1085546, 32'sd990486, -32'sd327051, -32'sd813657, -32'sd1156651, 32'sd0, 32'sd0, 32'sd0, 32'sd783029, -32'sd1816681, 32'sd967100, -32'sd217448, -32'sd2450784, -32'sd2238027, -32'sd835729, 32'sd1296603, 32'sd1161023, 32'sd1264906, 32'sd940389, 32'sd428220, -32'sd1010542, 32'sd1497801, -32'sd1385120, 32'sd628448, 32'sd501442, 32'sd568294, 32'sd118078, -32'sd1237663, -32'sd629940, 32'sd286401, -32'sd113922, -32'sd1886315, -32'sd688050, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd630609, -32'sd1534233, -32'sd2130408, -32'sd444781, 32'sd3665, 32'sd1703032, -32'sd1349740, -32'sd569804, 32'sd534080, 32'sd2163655, -32'sd422472, 32'sd354218, 32'sd785123, -32'sd64524, 32'sd1712739, -32'sd454659, -32'sd453992, 32'sd558529, 32'sd238452, 32'sd27395, 32'sd489690, 32'sd1160056, -32'sd984456, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd131406, -32'sd1449895, -32'sd1457162, -32'sd1703793, -32'sd479544, 32'sd1091970, 32'sd1364972, -32'sd877272, 32'sd758395, 32'sd276476, -32'sd724177, -32'sd1417311, -32'sd1870768, -32'sd716316, -32'sd582477, 32'sd226715, 32'sd504616, -32'sd2235461, -32'sd1380348, -32'sd531294, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd697992, 32'sd1581744, 32'sd1240270, 32'sd231190, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd97962, 32'sd429807, 32'sd2375367, 32'sd1664410, 32'sd918051, 32'sd1342903, -32'sd277424, 32'sd789527, 32'sd454923, 32'sd666699, -32'sd930225, 32'sd857398, -32'sd590928, 32'sd433234, 32'sd461026, 32'sd942206, 32'sd21882, 32'sd1893893, 32'sd436776, 32'sd759643, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1246977, 32'sd675171, 32'sd657212, -32'sd20096, 32'sd196763, 32'sd1009448, 32'sd1783388, -32'sd641586, -32'sd1241036, -32'sd524713, 32'sd1210904, -32'sd844881, 32'sd340307, 32'sd627579, -32'sd327484, -32'sd849258, 32'sd1201374, 32'sd994226, 32'sd178372, 32'sd1266658, 32'sd1542927, 32'sd2104104, 32'sd522817, 32'sd1275930, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1338354, 32'sd593935, 32'sd320554, -32'sd2063753, -32'sd60990, -32'sd359053, 32'sd996241, 32'sd880582, -32'sd148155, 32'sd710874, -32'sd1086928, -32'sd802438, -32'sd1527394, -32'sd783786, -32'sd821225, -32'sd1555595, 32'sd2051892, -32'sd336853, 32'sd278322, 32'sd1778400, -32'sd229191, -32'sd2750740, 32'sd118374, -32'sd752023, 32'sd382396, 32'sd0, 32'sd0, 32'sd473399, 32'sd119784, 32'sd6232, -32'sd1410359, -32'sd473082, 32'sd781549, 32'sd1936063, 32'sd913082, 32'sd1489468, 32'sd196175, 32'sd1529631, 32'sd2627981, 32'sd2971155, -32'sd67741, -32'sd396631, -32'sd2290023, -32'sd1517886, 32'sd367144, -32'sd43013, -32'sd679631, 32'sd2086785, 32'sd367203, -32'sd718009, -32'sd1105781, 32'sd263968, 32'sd82126, 32'sd381058, 32'sd0, 32'sd1372100, -32'sd414261, -32'sd459891, 32'sd754455, 32'sd1260773, 32'sd1120827, 32'sd3217177, 32'sd1398234, -32'sd453852, 32'sd2127266, 32'sd734567, 32'sd1891126, 32'sd1682209, -32'sd761472, 32'sd620354, 32'sd1943683, -32'sd1434695, 32'sd27934, 32'sd1108658, 32'sd585143, -32'sd869168, 32'sd290097, -32'sd1341807, -32'sd1550444, -32'sd420481, -32'sd194055, 32'sd300664, 32'sd0, 32'sd347620, 32'sd745646, 32'sd311461, 32'sd1684447, 32'sd111802, -32'sd393321, 32'sd750239, 32'sd126897, 32'sd847608, -32'sd916853, -32'sd562557, 32'sd41052, -32'sd806057, 32'sd939686, 32'sd1981811, 32'sd1068162, 32'sd2683518, 32'sd1525707, 32'sd456381, 32'sd59765, 32'sd695514, -32'sd230444, -32'sd1465772, -32'sd1270842, 32'sd977092, 32'sd838173, -32'sd93263, 32'sd868275, 32'sd578796, 32'sd1364726, 32'sd300680, 32'sd593903, -32'sd1043676, -32'sd496228, -32'sd399738, -32'sd743580, -32'sd1989227, -32'sd451077, -32'sd3059863, -32'sd2402429, -32'sd379905, 32'sd347256, 32'sd1184662, 32'sd844138, 32'sd1871126, 32'sd2004875, 32'sd1287890, 32'sd147821, 32'sd1261099, 32'sd123412, -32'sd1417766, -32'sd1240678, -32'sd343788, 32'sd168488, 32'sd1730448, 32'sd1020899, -32'sd790224, 32'sd110786, -32'sd985348, 32'sd111093, -32'sd1674201, -32'sd372520, -32'sd492139, 32'sd2401117, -32'sd2095606, -32'sd1146947, -32'sd175745, -32'sd2022122, -32'sd167381, -32'sd559211, -32'sd58002, -32'sd1634391, 32'sd552791, -32'sd1188380, 32'sd700316, 32'sd423866, 32'sd975485, 32'sd1489760, 32'sd629156, -32'sd2114796, -32'sd1315132, 32'sd265441, -32'sd862717, 32'sd859721, 32'sd164966, 32'sd641947, 32'sd1774192, 32'sd1120465, -32'sd2219477, -32'sd1181813, -32'sd1506287, -32'sd1006037, -32'sd2123574, -32'sd561623, 32'sd216201, -32'sd2171773, 32'sd426925, 32'sd535129, 32'sd2016932, -32'sd1028536, -32'sd2395017, -32'sd2687097, 32'sd85440, -32'sd409363, -32'sd53078, 32'sd1167632, 32'sd1353749, -32'sd163006, 32'sd1043629, -32'sd1437763, 32'sd215904, -32'sd220398, -32'sd183402, 32'sd932902, 32'sd1769085, 32'sd1178055, -32'sd1177390, 32'sd927404, 32'sd66543, 32'sd211952, -32'sd1499596, 32'sd477727, 32'sd621483, 32'sd337720, 32'sd4616, 32'sd2032180, -32'sd315533, -32'sd1445444, -32'sd1309694, -32'sd1551475, -32'sd380569, 32'sd454044, -32'sd895744, 32'sd65216, 32'sd1509713, 32'sd1566082, -32'sd1076409, 32'sd672619, 32'sd1078455, 32'sd59067, 32'sd1523546, -32'sd1071089, 32'sd992999, 32'sd444356, -32'sd410045, -32'sd1625820, -32'sd1174349, -32'sd1012882, -32'sd1121015, 32'sd1467857, -32'sd589514, -32'sd412531, -32'sd1094960, 32'sd696680, -32'sd1306262, -32'sd531549, 32'sd2013936, 32'sd319802, 32'sd179792, 32'sd1871473, 32'sd888644, 32'sd898254, 32'sd1925636, -32'sd1206931, -32'sd446871, 32'sd1660378, 32'sd1703431, 32'sd648916, 32'sd354426, 32'sd995216, -32'sd284229, 32'sd164038, 32'sd247568, -32'sd1843461, -32'sd881420, -32'sd1652100, 32'sd146943, 32'sd732573, -32'sd126405, -32'sd685049, 32'sd240837, 32'sd157101, 32'sd1282416, 32'sd3873440, 32'sd416572, 32'sd1537644, -32'sd96695, 32'sd981822, 32'sd322758, 32'sd280756, 32'sd982553, 32'sd1083689, 32'sd484525, -32'sd2078853, -32'sd1304666, -32'sd95203, 32'sd1546104, -32'sd673119, -32'sd503494, 32'sd277350, 32'sd736888, 32'sd403972, -32'sd217753, 32'sd338777, -32'sd2140521, -32'sd676278, 32'sd408561, 32'sd821286, -32'sd445626, 32'sd2797142, 32'sd2791118, 32'sd2108629, 32'sd2333993, -32'sd174729, -32'sd429353, -32'sd762600, -32'sd251149, 32'sd1635580, -32'sd451536, 32'sd1062084, -32'sd1059513, -32'sd624413, 32'sd483125, -32'sd629660, 32'sd1542547, 32'sd1576403, -32'sd744455, -32'sd172802, 32'sd2136670, 32'sd444068, 32'sd1051568, -32'sd1358233, 32'sd359343, 32'sd642365, 32'sd1189694, 32'sd2455405, 32'sd2459897, 32'sd1889808, 32'sd1606637, 32'sd2288165, -32'sd295879, -32'sd1369094, -32'sd285744, 32'sd173811, -32'sd201960, 32'sd581468, 32'sd308016, 32'sd315662, 32'sd1068910, 32'sd1062959, -32'sd250849, 32'sd301380, -32'sd341184, 32'sd46992, 32'sd298177, 32'sd1137161, -32'sd564060, 32'sd878398, -32'sd105589, -32'sd593293, -32'sd143161, 32'sd1136603, 32'sd1180487, 32'sd2963564, 32'sd1604540, -32'sd74522, -32'sd1373171, 32'sd959145, 32'sd588746, 32'sd922120, -32'sd469845, -32'sd41643, 32'sd163974, 32'sd672227, 32'sd887583, -32'sd1318612, 32'sd736253, 32'sd1081268, 32'sd257428, 32'sd417621, 32'sd482043, 32'sd1131658, -32'sd700069, -32'sd625047, -32'sd437604, 32'sd169869, 32'sd820390, -32'sd1382068, -32'sd156495, 32'sd229532, -32'sd1008558, -32'sd385570, -32'sd1646523, -32'sd2268997, -32'sd3070618, 32'sd214045, 32'sd42557, -32'sd493489, -32'sd1476174, 32'sd610678, 32'sd125370, 32'sd74616, 32'sd15659, -32'sd479310, -32'sd234112, -32'sd617622, -32'sd1296196, 32'sd0, -32'sd322152, 32'sd342226, -32'sd295907, -32'sd861246, -32'sd1665421, -32'sd2341336, 32'sd333292, -32'sd2992161, -32'sd1339354, -32'sd2150898, -32'sd2275214, -32'sd3233308, -32'sd211025, -32'sd180000, -32'sd2006308, -32'sd2106935, 32'sd74748, 32'sd1181433, 32'sd830614, 32'sd1162029, 32'sd1846945, -32'sd965757, 32'sd525412, 32'sd411626, 32'sd882578, -32'sd1033584, 32'sd168292, 32'sd33853, 32'sd546924, -32'sd101410, -32'sd1571301, -32'sd732626, -32'sd1715952, -32'sd1159153, -32'sd518553, -32'sd518317, -32'sd1392791, -32'sd3767653, -32'sd3388517, -32'sd3633599, -32'sd2151337, 32'sd1205542, -32'sd980696, -32'sd203754, 32'sd555178, -32'sd888340, -32'sd80250, -32'sd182219, -32'sd306149, -32'sd1161630, -32'sd2320967, -32'sd1294929, 32'sd703989, 32'sd2070113, 32'sd55632, 32'sd486029, 32'sd689107, 32'sd346989, -32'sd1287153, -32'sd2040778, -32'sd954038, -32'sd818453, -32'sd1844614, -32'sd490277, -32'sd1301941, -32'sd1009759, -32'sd3121456, -32'sd1639703, -32'sd664387, -32'sd74224, -32'sd602673, -32'sd1860429, -32'sd1556700, 32'sd1862798, 32'sd714795, -32'sd356978, -32'sd192923, -32'sd867813, -32'sd1435599, 32'sd46605, 32'sd997539, -32'sd218907, 32'sd1302445, 32'sd0, 32'sd268793, 32'sd463555, -32'sd543026, -32'sd680662, 32'sd274713, -32'sd321051, -32'sd966003, -32'sd349885, 32'sd498237, 32'sd338695, 32'sd583525, 32'sd640761, 32'sd1256490, 32'sd623259, -32'sd2789101, -32'sd2563432, 32'sd534469, -32'sd545027, -32'sd455683, -32'sd422131, 32'sd546643, -32'sd485502, -32'sd560372, 32'sd788235, -32'sd871468, 32'sd1730484, 32'sd760438, 32'sd838270, 32'sd277262, 32'sd1006669, 32'sd2279214, 32'sd2238503, 32'sd910743, 32'sd375216, 32'sd148238, -32'sd878143, 32'sd320652, 32'sd2191820, 32'sd1260699, 32'sd1495294, 32'sd345622, -32'sd936414, 32'sd302818, -32'sd1100921, -32'sd1193784, -32'sd380178, -32'sd1535787, 32'sd988273, -32'sd1022737, -32'sd713078, -32'sd1266997, -32'sd1738161, -32'sd196413, 32'sd1340235, 32'sd343289, 32'sd1226387, 32'sd90445, -32'sd54364, 32'sd1767821, 32'sd917521, -32'sd680333, 32'sd1805425, -32'sd253145, 32'sd1414994, 32'sd1135706, 32'sd1238559, 32'sd1476191, 32'sd1364378, 32'sd2139248, 32'sd2314101, -32'sd438301, -32'sd1222712, 32'sd883027, 32'sd1154862, -32'sd979112, -32'sd335047, -32'sd1651847, -32'sd3136353, -32'sd298804, -32'sd1582151, 32'sd1137172, 32'sd398679, 32'sd1112286, 32'sd0, 32'sd302385, 32'sd93987, 32'sd469591, 32'sd481575, 32'sd909487, 32'sd1736237, 32'sd1729437, 32'sd833580, 32'sd2750731, 32'sd2171882, 32'sd44417, -32'sd318579, 32'sd1505264, 32'sd138973, -32'sd1038206, 32'sd498074, 32'sd653501, 32'sd1642756, -32'sd402363, -32'sd3446, 32'sd150793, -32'sd613116, 32'sd171053, -32'sd57308, -32'sd1110288, -32'sd218507, 32'sd0, 32'sd0, 32'sd0, -32'sd536361, 32'sd1385760, 32'sd969731, 32'sd428176, -32'sd239883, 32'sd2337052, 32'sd2202286, -32'sd384765, 32'sd732332, -32'sd1712308, -32'sd463263, 32'sd801136, -32'sd1027117, -32'sd1155643, -32'sd1325554, 32'sd157656, -32'sd159322, -32'sd1285552, -32'sd831167, -32'sd359326, -32'sd362436, -32'sd175445, -32'sd422886, -32'sd172536, 32'sd409534, 32'sd0, 32'sd0, 32'sd0, 32'sd1108135, -32'sd1252603, -32'sd586859, 32'sd1713190, -32'sd172518, 32'sd448463, 32'sd545028, -32'sd1379112, -32'sd57372, -32'sd276231, -32'sd785004, 32'sd976357, 32'sd91873, -32'sd253687, -32'sd1027229, -32'sd64575, 32'sd793746, -32'sd1084490, -32'sd1323926, -32'sd1152354, -32'sd609237, 32'sd1042798, -32'sd250651, 32'sd1009284, 32'sd428968, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd690822, -32'sd594402, -32'sd324180, -32'sd122377, 32'sd25227, 32'sd340605, 32'sd958420, 32'sd826946, -32'sd1060680, -32'sd745873, -32'sd159585, -32'sd2183348, -32'sd459703, 32'sd942303, 32'sd1319033, 32'sd161581, 32'sd839607, -32'sd1274094, -32'sd200330, -32'sd509691, 32'sd930232, -32'sd127744, 32'sd427978, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1210590, 32'sd1564517, -32'sd29041, 32'sd1511801, -32'sd23019, -32'sd778311, 32'sd438120, 32'sd1525638, 32'sd530238, 32'sd362035, -32'sd464536, -32'sd1073735, -32'sd325587, -32'sd213057, 32'sd1280359, 32'sd590698, 32'sd465529, -32'sd347617, -32'sd362441, 32'sd406059, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd247845, 32'sd1118355, 32'sd1530120, 32'sd1258089, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd412159, -32'sd190007, -32'sd389368, 32'sd1065852, 32'sd121242, -32'sd1099582, 32'sd360961, 32'sd1318618, 32'sd1012606, 32'sd68829, -32'sd186593, 32'sd191391, 32'sd914077, -32'sd1079795, 32'sd295189, 32'sd2068493, 32'sd17620, 32'sd1613714, 32'sd1492188, 32'sd796018, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1313079, 32'sd341830, 32'sd953960, 32'sd1418873, 32'sd1576652, 32'sd689540, 32'sd188953, 32'sd707724, 32'sd771864, 32'sd1627201, 32'sd544069, 32'sd888521, 32'sd1585683, -32'sd685378, -32'sd1138860, 32'sd4416636, 32'sd2401822, 32'sd841665, -32'sd1095656, 32'sd1323001, 32'sd2277309, 32'sd2632527, -32'sd464203, 32'sd1660859, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd784145, 32'sd121193, -32'sd438909, 32'sd1651420, -32'sd305636, -32'sd1294841, 32'sd1890924, 32'sd1094296, 32'sd821769, -32'sd1756005, 32'sd16352, -32'sd2146585, -32'sd65895, 32'sd3018921, 32'sd771543, 32'sd251941, 32'sd1515643, 32'sd1183697, 32'sd454266, 32'sd1302840, 32'sd602036, 32'sd461168, 32'sd1085623, -32'sd782672, 32'sd1146048, 32'sd0, 32'sd0, 32'sd229667, 32'sd498674, -32'sd1346611, -32'sd1201925, -32'sd1365721, -32'sd707187, -32'sd3309439, -32'sd1226171, -32'sd357998, -32'sd72043, 32'sd561625, -32'sd757920, -32'sd934247, -32'sd1126424, -32'sd634183, 32'sd949038, 32'sd1664729, -32'sd559682, 32'sd1024219, 32'sd291570, 32'sd731978, -32'sd1396116, 32'sd1173695, 32'sd113063, -32'sd133200, -32'sd220577, -32'sd174553, 32'sd0, 32'sd78894, -32'sd545899, 32'sd1674380, -32'sd585292, -32'sd1378954, -32'sd674243, -32'sd1446175, -32'sd599129, -32'sd1383219, -32'sd402874, -32'sd2034160, 32'sd389780, -32'sd701906, -32'sd367913, -32'sd1104873, 32'sd1477441, 32'sd2462687, 32'sd1143153, 32'sd667923, 32'sd2018905, 32'sd510139, 32'sd478618, 32'sd1584093, 32'sd2091175, 32'sd168606, -32'sd192112, 32'sd360745, 32'sd0, 32'sd870390, 32'sd525714, 32'sd2260791, 32'sd177090, 32'sd819435, -32'sd9516, 32'sd1513581, -32'sd423591, -32'sd314515, -32'sd360467, 32'sd414247, 32'sd1741285, 32'sd620027, 32'sd963143, 32'sd862148, 32'sd1038707, -32'sd1058215, 32'sd51901, 32'sd1895003, -32'sd1132241, -32'sd1864894, -32'sd237699, 32'sd1890500, 32'sd1069012, 32'sd191005, 32'sd440451, 32'sd1849546, 32'sd1301111, 32'sd578043, -32'sd587702, -32'sd1242401, 32'sd199537, -32'sd627248, 32'sd1685547, -32'sd49058, 32'sd382615, -32'sd1660899, -32'sd282943, -32'sd308225, 32'sd829149, 32'sd822561, 32'sd107162, -32'sd1322067, -32'sd1838109, -32'sd1796738, 32'sd254240, -32'sd2931353, -32'sd1675365, -32'sd4707870, -32'sd3785400, -32'sd1473871, -32'sd466282, -32'sd249507, -32'sd1885237, -32'sd1084040, 32'sd228836, 32'sd200755, -32'sd2768579, -32'sd3220291, -32'sd1813949, -32'sd1466275, 32'sd738969, 32'sd154902, 32'sd1584234, -32'sd991860, 32'sd539523, 32'sd2064584, -32'sd67157, -32'sd2610, -32'sd421972, -32'sd3307783, -32'sd2053564, -32'sd1684003, -32'sd4368242, -32'sd4277299, -32'sd4032551, -32'sd5120317, -32'sd5203570, -32'sd2624777, -32'sd2438426, -32'sd2474657, -32'sd1227049, 32'sd1081845, 32'sd572276, -32'sd1231843, 32'sd240051, -32'sd789810, -32'sd1545495, -32'sd135822, -32'sd1390263, 32'sd1073117, 32'sd458732, 32'sd1064724, -32'sd227521, -32'sd790036, 32'sd1494623, -32'sd1874901, -32'sd1825440, -32'sd1593467, -32'sd4203932, -32'sd2494586, -32'sd3744679, -32'sd3496441, -32'sd2621751, -32'sd2234758, -32'sd1680978, -32'sd1466532, 32'sd626703, -32'sd1316450, 32'sd1238864, -32'sd802177, -32'sd397208, 32'sd797846, -32'sd976523, 32'sd431793, 32'sd760154, 32'sd1498848, 32'sd1922305, 32'sd1134939, -32'sd81050, -32'sd478665, -32'sd668156, 32'sd187900, 32'sd52853, -32'sd1870758, -32'sd2365326, -32'sd2828555, -32'sd2880839, -32'sd211627, -32'sd600285, -32'sd1505429, -32'sd1356588, -32'sd1524178, -32'sd2124989, 32'sd993664, 32'sd1991177, 32'sd826772, -32'sd861124, -32'sd1509765, 32'sd432984, 32'sd166508, -32'sd408685, -32'sd1908902, -32'sd1074974, -32'sd1219264, 32'sd952006, -32'sd283005, 32'sd1437953, -32'sd1722659, 32'sd236797, 32'sd1436358, 32'sd283845, -32'sd655285, 32'sd822726, -32'sd1476601, 32'sd224955, -32'sd1537693, -32'sd613571, 32'sd1308841, 32'sd88121, -32'sd547470, -32'sd52869, 32'sd3043232, 32'sd2012041, 32'sd1099208, -32'sd201032, 32'sd395233, 32'sd1061015, 32'sd309333, -32'sd419398, -32'sd118214, -32'sd1299884, -32'sd1353027, -32'sd1100246, 32'sd1022730, -32'sd748658, 32'sd657868, 32'sd104683, 32'sd1617978, -32'sd408538, 32'sd2129969, 32'sd2704011, -32'sd185177, 32'sd35891, -32'sd606589, -32'sd1439009, -32'sd108049, -32'sd895980, -32'sd667102, 32'sd2455795, 32'sd128224, 32'sd131027, -32'sd499592, -32'sd712443, -32'sd496429, 32'sd491375, 32'sd674323, -32'sd1555435, -32'sd621511, -32'sd3330691, -32'sd1148888, -32'sd1585133, 32'sd614055, 32'sd1306151, 32'sd1030940, -32'sd784417, -32'sd740041, -32'sd223842, 32'sd2456088, 32'sd3101668, 32'sd1999210, 32'sd1523141, 32'sd893018, 32'sd913382, 32'sd1062972, -32'sd605692, -32'sd1252126, -32'sd593900, -32'sd170134, -32'sd114239, -32'sd1192446, -32'sd13092, -32'sd862297, 32'sd244032, -32'sd426626, 32'sd284624, -32'sd383222, -32'sd622331, -32'sd1426021, -32'sd349064, 32'sd769124, -32'sd1269535, -32'sd112285, 32'sd1986807, 32'sd326220, -32'sd627729, 32'sd1872229, 32'sd1994780, 32'sd2115315, 32'sd3625818, 32'sd1370760, 32'sd1913472, 32'sd1439670, -32'sd924939, -32'sd838202, -32'sd238921, -32'sd1329171, -32'sd1999093, 32'sd853048, -32'sd47127, -32'sd84725, 32'sd4627, -32'sd835322, -32'sd821653, -32'sd62627, 32'sd370057, -32'sd920698, 32'sd1625283, -32'sd1316087, -32'sd595898, -32'sd1759258, -32'sd435896, 32'sd840771, 32'sd1663940, 32'sd1443601, 32'sd1397437, 32'sd1714398, 32'sd3395447, 32'sd1922557, 32'sd1956075, 32'sd2416376, -32'sd420531, 32'sd1636784, -32'sd41771, -32'sd77537, 32'sd1570054, -32'sd180653, -32'sd1687727, -32'sd889131, 32'sd297713, 32'sd529785, -32'sd1011795, -32'sd1112109, -32'sd1583170, -32'sd2178257, -32'sd311246, -32'sd1670048, -32'sd2234537, -32'sd1496730, 32'sd1132283, 32'sd352897, -32'sd36740, -32'sd389409, -32'sd434485, 32'sd741487, 32'sd187063, 32'sd3896196, 32'sd1073895, 32'sd1432594, 32'sd1720158, 32'sd2532813, 32'sd2275096, 32'sd2869187, 32'sd1880455, -32'sd8219, 32'sd1076793, 32'sd863143, 32'sd0, 32'sd634734, -32'sd161280, 32'sd1023703, -32'sd384209, -32'sd650220, 32'sd914928, -32'sd747824, 32'sd320784, -32'sd171149, 32'sd347151, -32'sd641745, 32'sd125361, -32'sd1457281, -32'sd2015397, -32'sd1395084, 32'sd1402438, 32'sd2623298, 32'sd1832349, -32'sd157639, 32'sd1907461, 32'sd2831972, 32'sd1588645, -32'sd427884, 32'sd7428, -32'sd859598, 32'sd33709, 32'sd895254, -32'sd21098, 32'sd175216, 32'sd1662923, -32'sd375392, -32'sd713634, 32'sd499888, -32'sd495795, 32'sd150070, 32'sd1003857, 32'sd470203, -32'sd577190, -32'sd397507, -32'sd1044341, 32'sd148573, 32'sd777405, -32'sd1125371, -32'sd105988, 32'sd1826135, 32'sd1413228, 32'sd2414158, 32'sd2002703, 32'sd2147052, 32'sd1522398, 32'sd769957, -32'sd595294, 32'sd1169950, 32'sd895304, 32'sd140397, 32'sd265829, -32'sd1595710, 32'sd1982693, -32'sd1241170, -32'sd733075, -32'sd730738, -32'sd2100660, 32'sd53480, 32'sd1155754, 32'sd584437, 32'sd136864, 32'sd1056010, -32'sd1017632, -32'sd1011839, 32'sd1013555, -32'sd1577186, 32'sd496337, 32'sd1428215, 32'sd552972, 32'sd328530, 32'sd967412, -32'sd104448, 32'sd443887, 32'sd2223745, -32'sd660512, 32'sd1690811, 32'sd8279, 32'sd1321821, 32'sd0, -32'sd109833, 32'sd557392, -32'sd776743, 32'sd408555, 32'sd164527, -32'sd188962, -32'sd493525, -32'sd620213, 32'sd1092594, 32'sd461317, 32'sd513937, -32'sd670407, 32'sd769898, -32'sd362944, -32'sd428243, -32'sd812164, 32'sd668251, -32'sd343297, 32'sd2006067, 32'sd1858939, 32'sd1834966, 32'sd2072154, 32'sd101985, -32'sd646030, 32'sd549850, -32'sd700061, 32'sd451316, 32'sd484767, -32'sd1032181, -32'sd870046, -32'sd1645496, -32'sd160302, 32'sd1084996, 32'sd527791, 32'sd1002274, -32'sd47696, 32'sd633697, 32'sd286376, -32'sd538309, 32'sd1447831, -32'sd394898, 32'sd24941, -32'sd995659, -32'sd1167769, -32'sd1776159, -32'sd838278, 32'sd1951764, 32'sd2456431, 32'sd35579, 32'sd1098454, 32'sd1116543, -32'sd1569004, -32'sd2661, 32'sd679191, 32'sd573422, 32'sd522026, 32'sd987258, 32'sd436860, 32'sd150764, -32'sd707809, 32'sd558257, 32'sd1282398, 32'sd2009200, -32'sd147210, 32'sd1432300, 32'sd899348, 32'sd741291, -32'sd748040, -32'sd1006030, -32'sd1768458, -32'sd1738465, -32'sd3065072, -32'sd2554119, -32'sd2094336, 32'sd148896, -32'sd530300, 32'sd135006, 32'sd277691, -32'sd742688, -32'sd916041, -32'sd429302, -32'sd634041, 32'sd180607, 32'sd0, 32'sd679472, 32'sd296466, -32'sd422758, 32'sd593065, 32'sd891168, 32'sd571757, 32'sd116864, 32'sd78145, 32'sd755785, 32'sd1165361, -32'sd332674, -32'sd121449, 32'sd946569, -32'sd2506600, -32'sd2829973, -32'sd1899279, -32'sd2212589, -32'sd3460944, -32'sd1812851, -32'sd1437297, -32'sd1652277, -32'sd13630, -32'sd2990019, 32'sd361914, 32'sd599769, -32'sd1973338, 32'sd0, 32'sd0, 32'sd0, -32'sd132785, 32'sd774351, 32'sd274197, -32'sd242692, -32'sd90794, 32'sd682667, -32'sd306679, -32'sd1602313, -32'sd2229131, -32'sd1655420, -32'sd1150332, -32'sd302818, -32'sd1238098, -32'sd736209, -32'sd707937, -32'sd1847231, -32'sd1623255, -32'sd2967820, -32'sd1557870, -32'sd242487, 32'sd415724, -32'sd3138493, -32'sd356836, 32'sd1113559, 32'sd807132, 32'sd0, 32'sd0, 32'sd0, 32'sd230131, 32'sd1000180, -32'sd822583, 32'sd891881, 32'sd45491, -32'sd831621, -32'sd1302205, 32'sd1703113, -32'sd1036707, 32'sd372689, -32'sd166270, -32'sd802327, -32'sd254780, 32'sd1455432, 32'sd2004537, -32'sd3189648, -32'sd1819300, -32'sd1160799, -32'sd1445935, -32'sd401527, -32'sd1771168, -32'sd2301863, -32'sd962728, 32'sd464136, -32'sd499094, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1087876, 32'sd1314298, 32'sd598442, -32'sd4403, 32'sd49008, -32'sd875331, 32'sd890615, -32'sd1112805, -32'sd1191311, 32'sd1655058, 32'sd843978, 32'sd2061178, -32'sd1651312, 32'sd284317, 32'sd706001, -32'sd848437, -32'sd292145, 32'sd1539721, -32'sd214379, 32'sd386969, -32'sd968092, 32'sd689664, 32'sd1024239, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1278289, 32'sd899151, 32'sd784584, -32'sd247835, -32'sd142717, 32'sd829689, 32'sd417692, 32'sd1380578, 32'sd1040816, 32'sd1337599, 32'sd573245, -32'sd302706, 32'sd1335273, 32'sd651084, 32'sd576181, -32'sd624683, 32'sd386598, -32'sd854047, -32'sd860946, 32'sd696557, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd151185, 32'sd354285, -32'sd158149, 32'sd298746, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd658113, 32'sd216015, 32'sd739978, 32'sd905405, 32'sd616998, 32'sd743448, 32'sd1103926, 32'sd791522, 32'sd1858802, 32'sd1589087, 32'sd225217, 32'sd1434566, 32'sd154471, 32'sd1474913, 32'sd233948, 32'sd1568182, 32'sd1254374, 32'sd274374, 32'sd1557158, 32'sd173247, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd301359, -32'sd440842, 32'sd241907, 32'sd334085, 32'sd295692, -32'sd799862, -32'sd199335, -32'sd549948, 32'sd715, 32'sd3125894, -32'sd255917, -32'sd194469, 32'sd1600869, 32'sd534764, -32'sd339804, 32'sd2881095, 32'sd1176873, 32'sd3119693, 32'sd2032915, 32'sd1278005, 32'sd1023483, 32'sd1184624, 32'sd638114, -32'sd104809, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1023679, 32'sd580083, -32'sd105633, -32'sd1732348, -32'sd737380, -32'sd2170791, 32'sd1962308, 32'sd1222082, 32'sd247002, 32'sd1453028, 32'sd2342742, 32'sd3239611, 32'sd1700141, 32'sd804973, -32'sd487037, 32'sd318925, -32'sd145609, -32'sd170356, 32'sd974166, 32'sd41452, -32'sd2363107, -32'sd1074388, -32'sd1614239, -32'sd835858, 32'sd252121, 32'sd0, 32'sd0, 32'sd770137, -32'sd1128110, 32'sd1721280, -32'sd62339, -32'sd773288, 32'sd407959, -32'sd1414363, 32'sd960852, -32'sd123432, -32'sd151690, -32'sd574321, -32'sd537087, 32'sd674760, 32'sd198593, 32'sd1012441, 32'sd926431, 32'sd994251, 32'sd783907, -32'sd320336, 32'sd1278558, 32'sd857336, 32'sd430867, -32'sd559162, -32'sd930824, 32'sd750831, -32'sd1767376, 32'sd1750440, 32'sd0, 32'sd985914, 32'sd405663, -32'sd1836637, -32'sd1232687, -32'sd1324634, -32'sd2939499, 32'sd68766, 32'sd52033, 32'sd1745391, 32'sd1182760, -32'sd1104896, -32'sd1876114, 32'sd1224048, 32'sd402274, 32'sd711764, 32'sd104984, 32'sd1770576, 32'sd484225, 32'sd895134, 32'sd1048796, 32'sd1231731, 32'sd1825299, 32'sd1715361, 32'sd1408304, -32'sd415965, -32'sd300716, -32'sd196633, 32'sd0, 32'sd1315712, -32'sd20060, -32'sd77406, 32'sd1257313, 32'sd817059, -32'sd586010, -32'sd1919389, 32'sd182416, 32'sd323926, 32'sd588286, -32'sd249914, 32'sd1602503, 32'sd725990, 32'sd135354, -32'sd381877, 32'sd433697, 32'sd1254918, 32'sd2804210, 32'sd511029, -32'sd435010, -32'sd1227114, 32'sd1297458, -32'sd1602162, 32'sd1821336, 32'sd281277, 32'sd992034, -32'sd1463153, 32'sd1105002, 32'sd131090, -32'sd180558, 32'sd15641, 32'sd1806283, -32'sd750405, -32'sd2472542, -32'sd1143842, 32'sd53720, -32'sd827066, 32'sd806622, 32'sd2395614, 32'sd1359938, 32'sd413444, 32'sd1169621, -32'sd69339, 32'sd705716, 32'sd2601640, 32'sd3030502, 32'sd1084351, 32'sd2072877, 32'sd2191590, -32'sd179322, -32'sd344808, -32'sd1189534, 32'sd817868, 32'sd196230, -32'sd110515, 32'sd804088, 32'sd1927874, -32'sd92743, 32'sd620166, 32'sd374918, -32'sd1014027, -32'sd2768015, 32'sd594372, 32'sd576127, -32'sd238484, -32'sd557325, 32'sd1955591, 32'sd3442431, 32'sd1008097, 32'sd989640, 32'sd293234, 32'sd967087, -32'sd439239, 32'sd296535, 32'sd1401907, 32'sd1449593, 32'sd1535056, -32'sd316601, -32'sd1473923, -32'sd227639, 32'sd535234, 32'sd1302699, -32'sd1091203, 32'sd790142, 32'sd2407073, -32'sd982738, 32'sd404604, 32'sd1197570, -32'sd594548, 32'sd233143, -32'sd235892, 32'sd362892, -32'sd2348249, -32'sd2567354, 32'sd307428, 32'sd1166088, 32'sd2504815, -32'sd674889, -32'sd2480174, -32'sd4904971, -32'sd4414175, -32'sd732274, 32'sd331495, 32'sd1299708, -32'sd623278, 32'sd1180551, -32'sd1421283, 32'sd514132, -32'sd506857, -32'sd880709, 32'sd156780, 32'sd1149850, 32'sd1142563, 32'sd1716947, -32'sd791632, 32'sd1458886, -32'sd564814, -32'sd1549880, -32'sd1818156, -32'sd31274, -32'sd775193, 32'sd1505442, 32'sd2309090, 32'sd1841591, 32'sd2136460, -32'sd3542784, -32'sd4252239, -32'sd3820433, -32'sd2484626, -32'sd348101, 32'sd189809, -32'sd1091480, -32'sd1158394, -32'sd1192957, -32'sd2698757, -32'sd759504, -32'sd526363, 32'sd273241, 32'sd960289, 32'sd1635399, 32'sd1633881, -32'sd365756, 32'sd1706015, -32'sd1118785, 32'sd1239176, -32'sd234411, -32'sd256630, 32'sd146365, 32'sd2177564, 32'sd865419, 32'sd2898074, 32'sd2519944, 32'sd77554, -32'sd4789234, -32'sd2812415, -32'sd1412563, 32'sd643881, 32'sd1719559, -32'sd740044, -32'sd2220511, -32'sd2221100, -32'sd3205131, -32'sd2529532, -32'sd1560780, -32'sd65162, 32'sd725487, 32'sd5247, 32'sd500464, -32'sd313835, 32'sd47574, -32'sd1170541, 32'sd292248, -32'sd735371, 32'sd382659, 32'sd1165548, 32'sd1542638, 32'sd942334, 32'sd1962972, 32'sd1465739, -32'sd732487, -32'sd2354302, -32'sd4510863, -32'sd1404393, -32'sd113956, -32'sd696729, 32'sd2295608, -32'sd2872770, -32'sd1429980, -32'sd540670, -32'sd3478108, -32'sd2818257, -32'sd619674, -32'sd1271475, 32'sd699852, 32'sd61468, -32'sd8902, -32'sd457777, 32'sd1513201, -32'sd353082, 32'sd1252441, 32'sd1107260, 32'sd1995040, 32'sd1780978, 32'sd1688954, 32'sd1491861, 32'sd1800767, -32'sd853319, -32'sd474025, -32'sd2879239, -32'sd2141607, -32'sd3175488, -32'sd2420340, -32'sd716361, -32'sd447421, 32'sd704758, -32'sd777898, -32'sd571957, -32'sd2591923, -32'sd2507315, 32'sd1313928, -32'sd960119, -32'sd996057, -32'sd335389, -32'sd212110, -32'sd639226, 32'sd224608, -32'sd1224557, 32'sd1283064, 32'sd644908, -32'sd717646, -32'sd63741, 32'sd992927, 32'sd551151, -32'sd846483, -32'sd961945, -32'sd584197, -32'sd2244361, -32'sd3112233, -32'sd2332646, -32'sd881053, -32'sd1985485, -32'sd800999, 32'sd405028, 32'sd106030, 32'sd486812, -32'sd945323, -32'sd2223968, 32'sd194748, -32'sd2467256, 32'sd413557, 32'sd1350456, -32'sd454203, 32'sd7541, 32'sd1796970, 32'sd254897, -32'sd290379, 32'sd428871, -32'sd2197691, -32'sd562364, -32'sd2994924, -32'sd1407348, -32'sd217420, -32'sd1655443, -32'sd1425972, -32'sd514813, -32'sd1630590, -32'sd1871033, -32'sd1083024, 32'sd49027, 32'sd1370963, 32'sd62568, -32'sd1079664, 32'sd1407937, -32'sd621038, -32'sd334577, 32'sd442273, -32'sd1699572, -32'sd353775, 32'sd777937, 32'sd73631, 32'sd572632, 32'sd987601, 32'sd618123, -32'sd2341496, -32'sd1714153, -32'sd2611562, -32'sd1697675, -32'sd2055903, -32'sd759046, 32'sd898807, 32'sd293454, -32'sd80298, -32'sd2871130, -32'sd1651669, -32'sd910313, -32'sd1126884, 32'sd820068, 32'sd1359690, 32'sd476638, 32'sd564444, 32'sd1499921, 32'sd2240524, -32'sd490039, -32'sd330153, -32'sd649748, 32'sd304042, -32'sd717820, 32'sd0, 32'sd237438, -32'sd817719, 32'sd147481, -32'sd1967116, -32'sd1671027, -32'sd590245, 32'sd1191986, -32'sd2521341, -32'sd1704681, 32'sd1108834, -32'sd1925734, -32'sd1575479, -32'sd707033, -32'sd2366394, -32'sd3227400, -32'sd1843556, 32'sd145618, 32'sd2046777, 32'sd1860880, 32'sd1093540, 32'sd1296402, 32'sd1270705, -32'sd1013148, 32'sd1112012, -32'sd430286, -32'sd211779, 32'sd1186207, -32'sd74499, 32'sd1469732, 32'sd943172, 32'sd499657, -32'sd1293005, -32'sd2891186, -32'sd1692314, -32'sd724737, -32'sd977541, 32'sd47216, -32'sd211524, -32'sd1194429, 32'sd581712, -32'sd2592048, -32'sd2702738, -32'sd2946959, -32'sd1122610, -32'sd133317, 32'sd1304404, 32'sd394447, 32'sd1120902, 32'sd904153, -32'sd694251, 32'sd99701, -32'sd1144650, -32'sd1345038, 32'sd270173, -32'sd713589, 32'sd157861, 32'sd385677, 32'sd1563653, 32'sd836328, -32'sd309454, -32'sd881072, -32'sd1253958, -32'sd945951, -32'sd2433001, -32'sd1019614, -32'sd3311204, -32'sd526844, -32'sd622253, -32'sd70685, -32'sd1280417, -32'sd2163217, -32'sd633802, 32'sd1762839, 32'sd982448, -32'sd1570604, 32'sd1468104, -32'sd895660, 32'sd852149, -32'sd576220, -32'sd53057, -32'sd5034, -32'sd658556, -32'sd921002, 32'sd0, -32'sd705687, -32'sd1495509, 32'sd1679043, 32'sd411570, -32'sd1802307, -32'sd924262, -32'sd1154500, -32'sd120793, -32'sd220710, -32'sd1015867, 32'sd162794, 32'sd481893, 32'sd356819, 32'sd779274, -32'sd46776, -32'sd807676, -32'sd664998, -32'sd1575163, -32'sd691110, 32'sd507860, 32'sd98797, 32'sd1120627, 32'sd892808, -32'sd123200, -32'sd1423190, -32'sd821427, 32'sd660854, 32'sd760852, 32'sd479826, 32'sd308287, 32'sd14733, 32'sd34105, -32'sd2293378, -32'sd1518572, -32'sd2097844, 32'sd143986, 32'sd862641, 32'sd948257, 32'sd1343322, 32'sd2333575, 32'sd2356031, 32'sd1483759, 32'sd2059427, 32'sd232494, -32'sd567976, 32'sd482129, -32'sd1752037, -32'sd266365, 32'sd807053, 32'sd2169075, 32'sd354685, -32'sd1511103, -32'sd304123, 32'sd204669, -32'sd283025, 32'sd473933, 32'sd672907, -32'sd316382, -32'sd1387364, -32'sd744419, -32'sd1496197, -32'sd2541868, -32'sd2010325, 32'sd39624, 32'sd949259, -32'sd1012570, 32'sd2364386, 32'sd2718807, 32'sd2617200, -32'sd58506, 32'sd2601155, 32'sd3095622, -32'sd1081475, 32'sd157076, 32'sd72169, 32'sd450181, -32'sd1447528, 32'sd1031612, 32'sd1123854, -32'sd1438046, -32'sd2227819, 32'sd755821, 32'sd1092767, 32'sd0, 32'sd926762, -32'sd474497, 32'sd194460, -32'sd1115775, 32'sd682816, -32'sd636870, 32'sd260300, 32'sd585242, 32'sd1829220, 32'sd1955938, 32'sd2370541, 32'sd744829, 32'sd1304002, 32'sd1167868, 32'sd280510, -32'sd532268, 32'sd1901603, 32'sd1325562, 32'sd1104566, -32'sd2115962, -32'sd253636, -32'sd67978, 32'sd1550484, -32'sd1759027, -32'sd1719141, -32'sd182889, 32'sd0, 32'sd0, 32'sd0, 32'sd42975, -32'sd391823, 32'sd635262, 32'sd1298032, 32'sd619288, 32'sd1097218, 32'sd2721143, 32'sd3518700, 32'sd2269373, 32'sd192481, 32'sd1724293, -32'sd161111, 32'sd605150, 32'sd1632033, 32'sd1417691, 32'sd2124276, 32'sd1710730, 32'sd2509060, -32'sd1018631, -32'sd553088, -32'sd50250, -32'sd1762786, 32'sd21147, 32'sd824989, 32'sd381240, 32'sd0, 32'sd0, 32'sd0, -32'sd269397, 32'sd626375, -32'sd214799, -32'sd282532, 32'sd523196, 32'sd1876529, 32'sd1083755, 32'sd2754264, 32'sd109358, 32'sd706327, 32'sd1505875, 32'sd2145831, -32'sd1759162, -32'sd109140, -32'sd392436, 32'sd218324, 32'sd302391, 32'sd239972, 32'sd1890966, -32'sd848623, 32'sd134675, -32'sd119267, 32'sd45421, -32'sd112464, 32'sd1225751, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd339430, 32'sd717728, -32'sd2486484, -32'sd388576, 32'sd577966, -32'sd436513, 32'sd2009430, 32'sd719274, 32'sd879085, 32'sd2473037, 32'sd955386, -32'sd65710, 32'sd1527808, 32'sd2069569, 32'sd589911, 32'sd1184557, 32'sd661945, -32'sd1342173, -32'sd957440, -32'sd820855, -32'sd416026, -32'sd204132, 32'sd393978, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1584280, 32'sd226725, -32'sd300752, 32'sd1445549, 32'sd1076395, 32'sd219296, 32'sd253741, 32'sd783957, 32'sd1091426, 32'sd1737012, 32'sd184003, 32'sd681044, -32'sd395582, 32'sd2173197, 32'sd31090, 32'sd63907, -32'sd17015, -32'sd251920, -32'sd195707, 32'sd325071, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd697995, -32'sd754669, 32'sd1245828, 32'sd1434839, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd600847, 32'sd881991, 32'sd1420787, 32'sd28539, -32'sd756489, 32'sd1255535, -32'sd174264, -32'sd1431226, -32'sd1871593, -32'sd269558, 32'sd328647, 32'sd107947, 32'sd1297844, -32'sd1244650, -32'sd1115551, -32'sd168978, -32'sd431027, -32'sd1010087, -32'sd214734, -32'sd317972, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd247388, -32'sd944274, -32'sd1994173, -32'sd1539860, 32'sd46667, 32'sd1047586, -32'sd720511, -32'sd1609090, -32'sd497675, -32'sd334446, -32'sd2855119, -32'sd645001, -32'sd2249854, -32'sd1570476, 32'sd541537, -32'sd1435313, -32'sd290305, 32'sd1421014, -32'sd755147, 32'sd329668, -32'sd2209607, -32'sd874294, 32'sd432532, -32'sd176660, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd175787, 32'sd1206524, 32'sd352909, 32'sd727521, -32'sd868548, -32'sd715472, -32'sd1771099, 32'sd1046109, -32'sd533933, -32'sd2107210, -32'sd1126474, -32'sd2484571, -32'sd914996, 32'sd1027038, 32'sd808657, -32'sd1652517, -32'sd2856477, -32'sd1046331, -32'sd350602, -32'sd867933, 32'sd655884, -32'sd1017715, 32'sd1258499, 32'sd399634, 32'sd562813, 32'sd0, 32'sd0, -32'sd507290, 32'sd862384, 32'sd81823, -32'sd523824, -32'sd1091999, -32'sd246180, -32'sd1080072, -32'sd3392897, -32'sd1301328, -32'sd1777648, -32'sd1094171, 32'sd271996, -32'sd1460644, -32'sd1146529, -32'sd669629, -32'sd582185, -32'sd267975, 32'sd182163, -32'sd907562, 32'sd1410378, -32'sd507774, 32'sd905522, -32'sd1849921, -32'sd1567404, 32'sd818983, 32'sd1332754, 32'sd197299, 32'sd0, -32'sd604938, -32'sd1651775, 32'sd473702, 32'sd38626, -32'sd2194694, -32'sd1987261, -32'sd2098121, -32'sd1465779, -32'sd1810817, -32'sd1986, 32'sd86636, 32'sd56409, 32'sd3718438, 32'sd1977290, 32'sd1077697, -32'sd1573349, -32'sd1071782, -32'sd37859, 32'sd1155993, -32'sd521709, -32'sd2478359, -32'sd226017, -32'sd3072711, -32'sd1437605, -32'sd1052811, 32'sd660609, -32'sd356992, 32'sd0, -32'sd366353, -32'sd423416, -32'sd1619884, -32'sd333011, -32'sd2924450, -32'sd1776096, -32'sd658775, -32'sd775839, -32'sd427366, -32'sd207511, 32'sd315001, 32'sd563685, 32'sd555490, 32'sd103763, 32'sd383980, 32'sd1477417, 32'sd1436961, 32'sd1809874, -32'sd4033, 32'sd963632, 32'sd993762, 32'sd721100, -32'sd1178871, -32'sd496265, -32'sd247449, -32'sd2044996, 32'sd942451, 32'sd552269, -32'sd247608, 32'sd233938, -32'sd318193, 32'sd965470, -32'sd2436486, -32'sd2509019, -32'sd1052720, -32'sd668952, 32'sd58557, 32'sd955904, 32'sd446130, 32'sd112200, -32'sd791021, 32'sd69832, 32'sd46699, 32'sd1553618, 32'sd1236898, 32'sd2391720, 32'sd2267720, 32'sd580692, -32'sd170613, -32'sd156670, 32'sd487196, 32'sd1629702, 32'sd450428, -32'sd2445193, -32'sd375128, 32'sd315663, 32'sd276600, 32'sd1149970, -32'sd1349461, -32'sd780123, -32'sd29595, 32'sd171402, -32'sd1417684, -32'sd241174, -32'sd639032, 32'sd954826, -32'sd350745, -32'sd219252, -32'sd1072676, 32'sd1276708, 32'sd3950988, 32'sd4429859, 32'sd2759101, 32'sd686959, 32'sd2081556, 32'sd48662, 32'sd645106, -32'sd803911, 32'sd1028668, 32'sd734140, 32'sd1609757, -32'sd1198547, -32'sd843065, -32'sd1138814, -32'sd1341708, -32'sd804798, -32'sd994461, 32'sd834918, -32'sd1325561, 32'sd2104453, 32'sd463467, -32'sd895956, 32'sd300914, 32'sd1327934, -32'sd477245, -32'sd152360, 32'sd1114096, 32'sd423893, 32'sd1228317, 32'sd1969011, 32'sd715825, 32'sd1149880, 32'sd1191389, 32'sd3791161, 32'sd1169317, -32'sd658191, 32'sd9140, 32'sd983153, -32'sd37382, -32'sd999688, -32'sd703367, 32'sd515392, 32'sd48682, -32'sd941396, 32'sd1174229, 32'sd355566, 32'sd936095, 32'sd198430, -32'sd1064812, -32'sd702333, 32'sd100250, 32'sd1069846, 32'sd1683238, 32'sd460707, -32'sd674207, 32'sd55654, 32'sd305556, -32'sd889554, -32'sd781239, -32'sd316279, 32'sd321309, 32'sd2161122, 32'sd2083926, 32'sd1175915, 32'sd411703, 32'sd1195929, -32'sd423550, -32'sd1130508, -32'sd396698, 32'sd419954, 32'sd1116258, 32'sd443014, -32'sd327177, -32'sd1143711, 32'sd910853, 32'sd312692, -32'sd211208, -32'sd1264384, -32'sd1859683, 32'sd1136507, -32'sd425262, -32'sd1469103, -32'sd552677, -32'sd2219486, -32'sd2502811, -32'sd627693, -32'sd731777, -32'sd690579, 32'sd409016, 32'sd2396119, 32'sd1612549, 32'sd835163, -32'sd1612362, 32'sd1241014, 32'sd1210364, 32'sd1379972, -32'sd1289791, 32'sd959685, 32'sd614915, -32'sd1959838, 32'sd730890, 32'sd1322469, 32'sd1260823, 32'sd1773272, -32'sd387574, -32'sd1232087, -32'sd2354375, 32'sd293, 32'sd630000, -32'sd2297007, -32'sd1520858, -32'sd880835, 32'sd240560, -32'sd392008, -32'sd825769, 32'sd1509686, 32'sd3981956, 32'sd2524599, 32'sd1049332, 32'sd246285, 32'sd773110, -32'sd390440, -32'sd255847, -32'sd342429, 32'sd435975, -32'sd110040, -32'sd1252084, 32'sd646497, 32'sd36257, -32'sd99897, 32'sd252581, 32'sd1805083, 32'sd1622484, -32'sd1280466, -32'sd2426416, -32'sd853011, -32'sd2024519, 32'sd1041863, -32'sd871567, 32'sd959321, -32'sd701368, -32'sd1436699, -32'sd1181495, 32'sd1314891, 32'sd3144205, 32'sd1604344, 32'sd999967, 32'sd317812, -32'sd424711, -32'sd3782930, -32'sd350272, 32'sd74295, -32'sd887968, -32'sd792967, -32'sd158906, -32'sd1025118, -32'sd1339712, 32'sd2354260, -32'sd341253, 32'sd2515553, 32'sd1307759, 32'sd2170626, 32'sd1694272, 32'sd507101, 32'sd1890566, 32'sd7071, -32'sd73519, 32'sd1280075, -32'sd1367008, -32'sd2549160, -32'sd175798, 32'sd2717209, 32'sd2120598, 32'sd245464, 32'sd1034100, 32'sd326030, -32'sd344498, -32'sd1212610, -32'sd579611, 32'sd2970920, -32'sd476986, -32'sd302438, -32'sd622737, 32'sd335162, -32'sd419041, 32'sd1344412, 32'sd2466394, 32'sd1125477, 32'sd3162566, 32'sd2405809, 32'sd1408262, 32'sd1803009, -32'sd1407950, -32'sd199845, -32'sd1410209, 32'sd468946, -32'sd1838909, -32'sd498367, 32'sd772619, 32'sd423683, 32'sd1126008, 32'sd1215881, 32'sd391096, 32'sd154932, -32'sd1350512, 32'sd618235, 32'sd478384, 32'sd2278824, -32'sd643171, -32'sd732568, -32'sd1041194, -32'sd544996, -32'sd804333, 32'sd1199365, 32'sd792257, 32'sd740367, 32'sd1252284, 32'sd1470252, 32'sd523344, -32'sd495834, -32'sd704491, 32'sd272097, 32'sd1182262, 32'sd191536, -32'sd87195, 32'sd95646, 32'sd309257, 32'sd1868906, -32'sd1416932, -32'sd1249167, -32'sd813810, 32'sd4396, -32'sd1848916, -32'sd390077, -32'sd1277557, 32'sd618789, -32'sd478435, 32'sd0, -32'sd1037316, 32'sd143712, -32'sd462149, 32'sd742101, -32'sd1103727, -32'sd517381, 32'sd1272341, 32'sd1515155, 32'sd3722855, 32'sd1754357, 32'sd1314525, -32'sd662069, -32'sd749972, -32'sd1179709, 32'sd290539, 32'sd524527, 32'sd506835, -32'sd794515, -32'sd458446, 32'sd1209983, 32'sd610769, -32'sd1094650, -32'sd1761379, 32'sd777707, 32'sd1047170, -32'sd721185, 32'sd665409, 32'sd1129525, 32'sd851434, 32'sd221755, -32'sd2175919, -32'sd1446592, -32'sd1763599, -32'sd749312, 32'sd811726, 32'sd339417, 32'sd1091037, 32'sd2116419, 32'sd1465479, 32'sd416711, 32'sd236447, 32'sd2042951, -32'sd145058, -32'sd1806498, 32'sd226418, -32'sd466299, 32'sd563946, 32'sd1152253, 32'sd1951235, -32'sd1139337, -32'sd544540, 32'sd388779, -32'sd770157, -32'sd864727, -32'sd524232, 32'sd418064, -32'sd544413, 32'sd250224, 32'sd656760, -32'sd2335133, -32'sd1847739, -32'sd138300, 32'sd1076179, 32'sd983781, -32'sd1291983, -32'sd506798, 32'sd836334, 32'sd2828818, 32'sd2194090, 32'sd1147390, -32'sd879891, 32'sd844805, -32'sd829930, 32'sd1512177, 32'sd2217101, -32'sd1059268, 32'sd1748450, -32'sd1647459, -32'sd1962275, 32'sd742866, -32'sd1032493, -32'sd508836, -32'sd1128555, 32'sd0, 32'sd1427645, -32'sd2661048, -32'sd163833, 32'sd527288, 32'sd806051, 32'sd37072, 32'sd228604, -32'sd721852, -32'sd2364030, -32'sd767136, -32'sd309946, 32'sd1720855, 32'sd689603, 32'sd49462, -32'sd2042641, -32'sd257972, 32'sd369542, 32'sd1762193, 32'sd1449516, 32'sd177683, 32'sd2731222, -32'sd1128280, -32'sd2115937, -32'sd585282, 32'sd1123384, 32'sd1006503, -32'sd637568, 32'sd238717, -32'sd1268457, -32'sd450988, 32'sd125703, 32'sd952823, 32'sd1015158, 32'sd1959731, 32'sd1594067, -32'sd433751, -32'sd2568065, -32'sd352255, -32'sd215076, 32'sd1041869, -32'sd1075894, 32'sd84495, -32'sd1712200, 32'sd793526, -32'sd1786879, 32'sd347518, 32'sd498646, 32'sd471342, 32'sd761772, 32'sd1249361, -32'sd1400970, -32'sd911694, 32'sd609310, 32'sd1764165, -32'sd719592, 32'sd70375, -32'sd1323843, 32'sd20564, 32'sd654420, -32'sd649719, 32'sd1457979, 32'sd2406131, -32'sd176583, 32'sd228901, 32'sd957808, -32'sd71024, 32'sd420129, 32'sd295660, -32'sd847396, -32'sd1744603, -32'sd1370523, -32'sd634778, 32'sd231946, 32'sd903085, -32'sd515460, -32'sd432758, 32'sd2176874, 32'sd930181, -32'sd1477652, -32'sd682604, -32'sd763686, 32'sd2058505, 32'sd72104, 32'sd0, -32'sd818334, -32'sd256652, 32'sd326313, -32'sd2106478, -32'sd1558096, 32'sd576846, 32'sd54395, 32'sd891063, -32'sd397478, -32'sd1117255, 32'sd988921, 32'sd202265, -32'sd186014, -32'sd381800, 32'sd735814, -32'sd730173, -32'sd1297164, -32'sd1352059, -32'sd764421, 32'sd1640114, -32'sd48799, 32'sd1351658, 32'sd842695, -32'sd172310, 32'sd371289, -32'sd469544, 32'sd0, 32'sd0, 32'sd0, 32'sd108038, 32'sd1527648, 32'sd1673492, 32'sd297826, -32'sd539032, -32'sd320472, 32'sd978263, 32'sd859576, -32'sd1009635, -32'sd1715234, -32'sd597619, -32'sd1741486, -32'sd986454, -32'sd769097, 32'sd385856, -32'sd938142, -32'sd335117, 32'sd1450018, 32'sd951185, -32'sd115629, -32'sd246175, 32'sd445766, 32'sd1732943, -32'sd575335, -32'sd190863, 32'sd0, 32'sd0, 32'sd0, 32'sd1022813, -32'sd820949, 32'sd87245, 32'sd1436624, -32'sd51431, 32'sd366003, 32'sd979322, 32'sd181526, -32'sd756306, -32'sd568650, -32'sd1996741, -32'sd3440535, -32'sd771249, -32'sd1507847, -32'sd2371243, -32'sd2959325, -32'sd1104949, -32'sd112017, 32'sd433311, -32'sd556654, 32'sd721280, -32'sd601282, 32'sd90144, 32'sd1321864, -32'sd773987, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5538, -32'sd130788, 32'sd1315185, 32'sd1427814, 32'sd994888, 32'sd1081279, -32'sd3310922, -32'sd1871905, -32'sd316419, -32'sd24572, 32'sd639433, 32'sd956471, 32'sd809029, -32'sd177997, -32'sd1051141, -32'sd1046840, 32'sd288874, -32'sd1163830, -32'sd398682, -32'sd930422, -32'sd995934, -32'sd444362, 32'sd106551, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd887778, -32'sd936233, -32'sd100999, -32'sd1332, -32'sd105015, -32'sd159775, 32'sd1245462, 32'sd1461367, -32'sd1021826, -32'sd1866862, -32'sd1261121, -32'sd236194, -32'sd183309, 32'sd548043, 32'sd8713, -32'sd399412, -32'sd346531, -32'sd918877, -32'sd762318, -32'sd739294, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd797822, 32'sd1256295, 32'sd194900, 32'sd1651896, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd73006, -32'sd342860, -32'sd326724, -32'sd773462, 32'sd349894, 32'sd40747, 32'sd837095, 32'sd76496, 32'sd321804, -32'sd366393, -32'sd1316816, 32'sd119846, -32'sd527780, 32'sd1046919, -32'sd36529, 32'sd1411627, 32'sd851524, 32'sd280503, 32'sd803718, -32'sd130535, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd751115, -32'sd89608, -32'sd222121, -32'sd983447, -32'sd400675, -32'sd955460, -32'sd250344, -32'sd1949604, -32'sd569618, 32'sd1545113, 32'sd1647797, 32'sd554206, 32'sd1334204, 32'sd853595, 32'sd1969327, 32'sd1548989, 32'sd332119, 32'sd1629367, 32'sd1421562, 32'sd2093035, 32'sd1691241, 32'sd323764, 32'sd957433, -32'sd253831, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd90164, -32'sd158303, 32'sd521077, 32'sd966799, 32'sd795239, -32'sd1503871, -32'sd3286845, 32'sd1727349, -32'sd202811, 32'sd698044, -32'sd593096, 32'sd1877892, 32'sd1015364, -32'sd1743687, -32'sd170074, -32'sd1972257, -32'sd659426, -32'sd1228890, 32'sd117717, 32'sd1554738, -32'sd110376, 32'sd1049622, 32'sd537909, 32'sd459718, -32'sd2531379, 32'sd0, 32'sd0, 32'sd504363, 32'sd162665, 32'sd297029, 32'sd944294, 32'sd715359, 32'sd318603, -32'sd236053, -32'sd2409504, 32'sd500261, -32'sd835479, -32'sd141590, -32'sd420922, -32'sd1799322, -32'sd3377855, -32'sd3364581, -32'sd198851, 32'sd271688, 32'sd170658, -32'sd438262, -32'sd1299130, 32'sd363245, -32'sd102572, -32'sd893512, -32'sd929878, -32'sd1782830, -32'sd738943, 32'sd842839, 32'sd0, -32'sd269476, -32'sd1339114, 32'sd423387, 32'sd1686819, 32'sd1159678, -32'sd703171, -32'sd982202, -32'sd518525, -32'sd976547, -32'sd309048, 32'sd451286, -32'sd1921011, -32'sd1539311, -32'sd437134, -32'sd925228, -32'sd1307176, 32'sd1068468, -32'sd555227, 32'sd2188987, -32'sd521184, 32'sd1285409, -32'sd83279, 32'sd502808, 32'sd214676, -32'sd2635711, -32'sd1055790, -32'sd27148, 32'sd0, -32'sd297636, -32'sd1082191, 32'sd171101, -32'sd2280968, 32'sd21722, 32'sd1501228, 32'sd470296, -32'sd1537098, -32'sd1312335, -32'sd1110161, -32'sd654148, -32'sd377684, -32'sd1181725, -32'sd2708671, 32'sd115232, -32'sd837915, -32'sd1230450, -32'sd264654, 32'sd619473, 32'sd3197189, 32'sd2362051, 32'sd931082, -32'sd472539, -32'sd969657, -32'sd272188, -32'sd761247, 32'sd1772724, 32'sd467309, 32'sd281921, 32'sd172859, -32'sd1332168, 32'sd196360, -32'sd1159963, 32'sd1284974, -32'sd468396, 32'sd500240, 32'sd556617, 32'sd543999, -32'sd102392, 32'sd562073, -32'sd1760427, -32'sd2723186, 32'sd1846905, 32'sd1240062, 32'sd385214, 32'sd1120105, 32'sd172325, 32'sd2220230, 32'sd1188675, 32'sd1471657, 32'sd1130948, -32'sd2158771, -32'sd472507, 32'sd1710495, 32'sd34494, 32'sd740689, 32'sd618792, -32'sd901076, -32'sd359166, -32'sd636953, -32'sd607270, -32'sd970634, 32'sd1102913, 32'sd778106, 32'sd1636090, 32'sd2020299, 32'sd3157301, 32'sd1549964, -32'sd307146, 32'sd309527, -32'sd1561152, 32'sd726559, 32'sd12210, 32'sd91200, -32'sd610924, 32'sd640491, 32'sd1493260, 32'sd1007948, -32'sd2569363, -32'sd1173480, 32'sd1821774, 32'sd448865, -32'sd550672, 32'sd622980, 32'sd635894, -32'sd2154548, -32'sd340942, -32'sd303486, -32'sd2279145, -32'sd2121410, -32'sd1641076, -32'sd1906025, -32'sd2269890, 32'sd2342187, 32'sd3746926, 32'sd650458, 32'sd385253, -32'sd2498868, -32'sd985843, -32'sd1651528, -32'sd675652, -32'sd1425913, -32'sd1745164, 32'sd458590, 32'sd325105, -32'sd1762923, -32'sd1438684, -32'sd1112617, 32'sd2931855, -32'sd917471, -32'sd1893655, 32'sd1068848, 32'sd1535997, -32'sd142940, -32'sd1832122, -32'sd239149, -32'sd1851361, -32'sd2275327, -32'sd2535002, -32'sd1925822, -32'sd2395379, 32'sd289744, 32'sd3760255, -32'sd302136, -32'sd1059592, -32'sd2795145, -32'sd2124425, 32'sd1104089, -32'sd363588, -32'sd2349040, -32'sd2375418, -32'sd1648963, -32'sd2146373, -32'sd1746170, -32'sd3297684, -32'sd511933, 32'sd963697, 32'sd617150, -32'sd1974973, 32'sd1424507, -32'sd193941, -32'sd1045697, 32'sd713044, 32'sd773148, -32'sd2308598, -32'sd2436, -32'sd2061831, -32'sd917834, -32'sd2097210, -32'sd469809, 32'sd3262573, 32'sd2625345, 32'sd865620, -32'sd1728509, -32'sd1551043, 32'sd1250952, -32'sd334771, -32'sd849550, 32'sd56326, 32'sd944855, -32'sd604507, -32'sd592673, -32'sd1246046, -32'sd1158487, -32'sd471852, 32'sd722324, -32'sd567532, 32'sd527715, -32'sd523704, 32'sd1167529, 32'sd698405, -32'sd553427, -32'sd1640189, -32'sd805722, -32'sd1790943, -32'sd2386429, -32'sd2074561, -32'sd899133, 32'sd1954569, 32'sd2023434, -32'sd1603329, -32'sd2366773, -32'sd1462826, -32'sd619163, 32'sd222896, -32'sd88952, -32'sd988826, 32'sd1673529, 32'sd702457, 32'sd617020, -32'sd1406979, -32'sd1174305, -32'sd490152, 32'sd280980, 32'sd120928, -32'sd343695, 32'sd837850, -32'sd594076, -32'sd841633, 32'sd305017, 32'sd647201, -32'sd14243, -32'sd1238693, -32'sd2297062, -32'sd1492684, 32'sd1648833, 32'sd179406, -32'sd970708, -32'sd2424407, -32'sd2812101, -32'sd328474, 32'sd427499, 32'sd133516, 32'sd840362, 32'sd2165119, 32'sd707493, 32'sd1004191, 32'sd1881152, -32'sd576283, -32'sd3071962, -32'sd1189891, 32'sd157467, -32'sd39751, 32'sd773321, 32'sd806776, 32'sd802797, -32'sd326806, 32'sd310203, 32'sd79188, -32'sd2073724, 32'sd19944, -32'sd2325686, 32'sd480094, 32'sd2587228, 32'sd1629018, -32'sd423276, -32'sd123569, -32'sd1225241, 32'sd1592600, 32'sd524613, -32'sd2277121, 32'sd1782530, 32'sd928556, 32'sd3272956, 32'sd3362010, 32'sd1717090, -32'sd1224400, -32'sd2021820, 32'sd943947, 32'sd621473, 32'sd720313, -32'sd721382, 32'sd270035, -32'sd389464, -32'sd691248, -32'sd2425902, -32'sd2443361, -32'sd1674866, -32'sd699667, -32'sd581382, 32'sd577950, 32'sd2654958, 32'sd1312640, -32'sd651958, -32'sd502408, 32'sd1130611, 32'sd1454753, 32'sd883848, 32'sd1243708, 32'sd1368780, 32'sd1645177, 32'sd771359, 32'sd1187666, -32'sd1589587, -32'sd757575, -32'sd2619084, 32'sd200790, 32'sd478786, -32'sd586856, -32'sd16043, 32'sd472642, -32'sd2264093, -32'sd1511205, -32'sd1545163, -32'sd243911, -32'sd1645240, -32'sd1801100, 32'sd329252, 32'sd1310275, -32'sd780974, 32'sd346470, -32'sd488740, -32'sd527472, -32'sd615492, 32'sd532345, 32'sd760220, 32'sd186451, 32'sd199887, -32'sd2020326, -32'sd1058180, -32'sd1495066, -32'sd109650, -32'sd2647538, -32'sd793047, 32'sd993128, 32'sd1223129, 32'sd211466, 32'sd0, 32'sd471030, -32'sd1287460, 32'sd101568, 32'sd1122834, 32'sd986308, -32'sd2821858, -32'sd1502446, 32'sd1078699, -32'sd272261, 32'sd2015769, -32'sd433444, -32'sd1815518, -32'sd1373174, 32'sd1290447, 32'sd24233, 32'sd1606112, -32'sd1541755, -32'sd452475, -32'sd1875109, -32'sd781567, -32'sd1934365, -32'sd1573998, -32'sd1736930, -32'sd2730831, 32'sd472647, -32'sd920269, -32'sd416709, -32'sd626982, 32'sd633896, 32'sd601124, -32'sd370156, 32'sd265477, -32'sd2241886, -32'sd2084746, -32'sd692271, 32'sd1150955, 32'sd688307, 32'sd346861, 32'sd1055492, 32'sd401307, 32'sd497420, 32'sd1593721, 32'sd2159963, -32'sd733057, -32'sd621806, -32'sd57754, 32'sd12872, -32'sd2758077, -32'sd2216927, -32'sd974679, -32'sd827900, -32'sd1464306, -32'sd1795706, -32'sd2274770, 32'sd643990, 32'sd193631, -32'sd724711, 32'sd509554, -32'sd984462, 32'sd360860, 32'sd141079, -32'sd2076300, -32'sd2021087, 32'sd1067520, 32'sd1010657, 32'sd2572091, 32'sd1415503, 32'sd947853, -32'sd1752953, 32'sd874558, -32'sd353551, -32'sd926851, -32'sd3214723, -32'sd551160, 32'sd1391338, -32'sd337846, -32'sd1695719, -32'sd399087, 32'sd1236501, 32'sd1265257, -32'sd334309, -32'sd982653, 32'sd1521544, 32'sd0, -32'sd1163032, 32'sd928628, -32'sd1925746, -32'sd1472113, -32'sd2594488, -32'sd593609, -32'sd2316943, -32'sd1032229, 32'sd802582, 32'sd2410078, 32'sd2328639, 32'sd911488, -32'sd2562305, -32'sd1012224, -32'sd2379807, -32'sd2071371, -32'sd2041601, -32'sd493039, -32'sd759824, -32'sd1780785, -32'sd1378780, -32'sd475985, 32'sd1174696, 32'sd1169856, -32'sd74047, -32'sd492427, 32'sd861390, -32'sd180979, 32'sd551025, 32'sd261748, -32'sd587263, -32'sd1882426, -32'sd3058687, -32'sd3418538, -32'sd2526629, -32'sd1181476, -32'sd858919, -32'sd1008482, 32'sd472963, 32'sd1712912, 32'sd1148985, -32'sd1030883, -32'sd1740551, -32'sd1671853, -32'sd916604, -32'sd1717401, -32'sd2388276, -32'sd3532044, -32'sd248606, 32'sd2123119, 32'sd2417622, 32'sd2120048, -32'sd67951, 32'sd28702, 32'sd527873, -32'sd986911, -32'sd84240, 32'sd573527, -32'sd584505, -32'sd1863637, -32'sd732044, -32'sd2145302, 32'sd285121, -32'sd1284757, 32'sd390338, -32'sd673358, -32'sd1121606, 32'sd1794105, 32'sd3072630, 32'sd1551755, 32'sd1482748, 32'sd90, -32'sd1962684, -32'sd1124650, -32'sd1037274, -32'sd1802886, -32'sd254673, 32'sd1119683, -32'sd490287, -32'sd749194, 32'sd1361600, 32'sd1762930, -32'sd344439, 32'sd0, 32'sd863338, -32'sd410897, 32'sd564667, -32'sd3220712, -32'sd2001957, -32'sd1086104, -32'sd583806, 32'sd1529415, 32'sd1863909, -32'sd150872, -32'sd1235383, 32'sd1559735, 32'sd2136322, 32'sd420781, -32'sd1814969, 32'sd530563, -32'sd553780, -32'sd1160869, -32'sd1385641, -32'sd923984, 32'sd1123280, 32'sd1373243, 32'sd1015820, -32'sd1100662, 32'sd1070221, -32'sd187124, 32'sd0, 32'sd0, 32'sd0, -32'sd51298, 32'sd553670, -32'sd1896092, -32'sd1890434, -32'sd801425, -32'sd1128268, -32'sd2065892, -32'sd2274125, -32'sd610241, -32'sd32990, 32'sd1861527, 32'sd455354, -32'sd455752, 32'sd611966, 32'sd1994558, -32'sd75842, -32'sd2531701, -32'sd1803089, -32'sd1657419, -32'sd364946, -32'sd983949, -32'sd1643517, -32'sd742790, -32'sd649772, 32'sd1148540, 32'sd0, 32'sd0, 32'sd0, -32'sd182425, -32'sd82610, -32'sd145860, 32'sd983134, -32'sd658036, 32'sd371948, -32'sd2451761, -32'sd1557248, -32'sd508250, -32'sd685052, 32'sd1667995, -32'sd510995, 32'sd1483111, 32'sd4095411, -32'sd17692, -32'sd936100, 32'sd160374, -32'sd910389, -32'sd1442087, -32'sd1858636, -32'sd1433585, 32'sd525260, 32'sd1297860, -32'sd101626, 32'sd272929, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd464419, -32'sd1270064, -32'sd1713960, 32'sd447663, 32'sd448785, 32'sd1900885, 32'sd468058, 32'sd515913, -32'sd1307035, -32'sd682706, 32'sd1955688, -32'sd944812, -32'sd668457, -32'sd396905, -32'sd653860, 32'sd156537, -32'sd427972, 32'sd637122, -32'sd802869, -32'sd947940, 32'sd193375, 32'sd312538, 32'sd1047927, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd288484, -32'sd505767, 32'sd546993, -32'sd231018, 32'sd351775, 32'sd513717, -32'sd642531, -32'sd489447, -32'sd915444, 32'sd1008036, -32'sd275073, 32'sd203428, -32'sd533352, 32'sd812006, 32'sd556138, 32'sd657511, -32'sd243157, -32'sd175913, -32'sd584003, -32'sd257273, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1929677, -32'sd738918, -32'sd769634, -32'sd61933, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1813, 32'sd406387, 32'sd826447, -32'sd1370269, -32'sd551992, -32'sd709482, 32'sd321795, 32'sd1193723, -32'sd1099316, -32'sd929670, 32'sd619928, 32'sd1817364, -32'sd217737, -32'sd74985, 32'sd1261737, 32'sd601950, -32'sd803116, 32'sd979676, 32'sd262514, 32'sd22938, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd99351, -32'sd136364, -32'sd384786, -32'sd33894, -32'sd621840, -32'sd1451602, -32'sd584040, -32'sd1261707, 32'sd701206, -32'sd1323204, -32'sd103024, -32'sd2667463, -32'sd1260270, 32'sd2235924, 32'sd1313673, -32'sd599328, -32'sd594163, 32'sd1258028, -32'sd1059813, -32'sd131818, 32'sd243249, 32'sd578820, 32'sd670360, -32'sd205694, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd881143, -32'sd38079, 32'sd500016, 32'sd236645, -32'sd250081, -32'sd2287679, -32'sd974250, 32'sd898958, 32'sd326831, 32'sd576589, -32'sd612068, 32'sd185213, 32'sd62493, 32'sd1052921, -32'sd2638156, -32'sd3192526, -32'sd1926053, -32'sd1708101, -32'sd1371855, 32'sd632830, 32'sd777106, 32'sd220218, -32'sd1430013, -32'sd718034, -32'sd234585, 32'sd0, 32'sd0, -32'sd45975, 32'sd892342, 32'sd1164711, -32'sd616272, -32'sd668335, -32'sd2628475, 32'sd99351, 32'sd38623, 32'sd1641022, 32'sd722273, 32'sd637606, -32'sd2559829, -32'sd3102268, 32'sd773107, 32'sd654137, 32'sd916344, 32'sd1501389, -32'sd1127592, -32'sd1108436, -32'sd2157328, -32'sd1787580, -32'sd2280807, -32'sd263402, -32'sd1988020, -32'sd481755, -32'sd540345, -32'sd127605, 32'sd0, -32'sd183446, -32'sd826660, -32'sd651934, -32'sd1327697, -32'sd814958, 32'sd348023, 32'sd1877306, -32'sd1139970, 32'sd356121, 32'sd928468, 32'sd1397720, 32'sd1752405, 32'sd1611978, 32'sd3672077, -32'sd1099240, -32'sd865352, -32'sd253417, -32'sd3208036, -32'sd1939816, 32'sd602235, 32'sd2212286, -32'sd305591, -32'sd2612587, -32'sd1082666, -32'sd726008, 32'sd985800, -32'sd1124192, 32'sd0, -32'sd295902, -32'sd509431, 32'sd1283531, -32'sd1107146, 32'sd2090179, 32'sd2314255, 32'sd1610233, 32'sd214820, -32'sd236784, 32'sd1937936, 32'sd1438854, 32'sd4040806, 32'sd1144459, -32'sd1090888, -32'sd521946, -32'sd4129890, -32'sd2511130, -32'sd2525266, -32'sd864091, -32'sd506591, 32'sd634520, -32'sd1451284, -32'sd157640, -32'sd566520, 32'sd1259640, 32'sd1224677, 32'sd211765, -32'sd132434, 32'sd690269, -32'sd744001, 32'sd1587378, -32'sd1607833, 32'sd689290, 32'sd2206334, 32'sd986993, 32'sd1133826, 32'sd437103, 32'sd795480, 32'sd878169, 32'sd997485, -32'sd478361, -32'sd150740, -32'sd1858114, -32'sd404218, -32'sd814463, -32'sd908228, 32'sd1245597, 32'sd1261913, 32'sd2527057, 32'sd1229741, -32'sd1290374, -32'sd1382802, 32'sd667198, -32'sd1489754, 32'sd1098160, -32'sd489162, -32'sd932452, 32'sd119217, -32'sd1070562, 32'sd205450, 32'sd1520234, 32'sd2034982, 32'sd2948319, 32'sd1638994, 32'sd617193, 32'sd2282361, 32'sd629544, 32'sd1813122, 32'sd169239, -32'sd570961, -32'sd156125, 32'sd1066815, 32'sd1108837, 32'sd829289, 32'sd2899700, 32'sd2757146, 32'sd1582356, 32'sd2618501, 32'sd2317901, 32'sd1525346, 32'sd1403592, 32'sd672258, 32'sd1647856, 32'sd195176, -32'sd901314, 32'sd529928, -32'sd1069023, 32'sd716735, -32'sd258781, 32'sd1384951, 32'sd1268462, -32'sd456144, -32'sd349460, 32'sd1836067, 32'sd3378064, 32'sd1195007, 32'sd1795641, 32'sd1479041, 32'sd2088925, 32'sd1757675, 32'sd1096826, 32'sd2965572, 32'sd2878945, 32'sd4475687, 32'sd2350681, 32'sd3127102, 32'sd527652, 32'sd1871730, 32'sd1990939, 32'sd893202, 32'sd1234092, -32'sd416530, -32'sd646682, 32'sd393644, -32'sd2386291, -32'sd405712, -32'sd894231, 32'sd45047, -32'sd301009, 32'sd115466, -32'sd1787463, 32'sd616026, 32'sd1623847, 32'sd878680, 32'sd892762, 32'sd1447250, 32'sd2962844, -32'sd137934, 32'sd98552, 32'sd4286829, 32'sd4220122, 32'sd2767781, 32'sd2534627, 32'sd1686259, -32'sd6555, 32'sd3133819, 32'sd1700606, -32'sd472468, 32'sd924802, 32'sd217055, -32'sd656194, 32'sd255601, -32'sd1388229, -32'sd995037, 32'sd959605, 32'sd1033172, 32'sd1431475, -32'sd1479769, -32'sd1873701, -32'sd1133763, 32'sd1034359, -32'sd3536082, -32'sd2047099, -32'sd1247723, -32'sd41601, -32'sd674324, -32'sd554050, 32'sd990149, 32'sd1000650, 32'sd1195693, 32'sd856765, 32'sd634000, -32'sd1011897, 32'sd538587, 32'sd239492, 32'sd1439722, 32'sd1293477, 32'sd438777, 32'sd618648, 32'sd479515, -32'sd119974, -32'sd779512, -32'sd1128227, -32'sd1188008, 32'sd2030568, 32'sd2069065, 32'sd1352532, -32'sd2252295, -32'sd345657, -32'sd1560374, -32'sd1542185, -32'sd2031243, -32'sd1745644, -32'sd3162851, 32'sd63402, -32'sd1978575, -32'sd760057, -32'sd1635609, 32'sd1136266, -32'sd112696, -32'sd1547763, -32'sd854660, 32'sd2113612, -32'sd354604, -32'sd1018542, -32'sd380807, 32'sd1317770, 32'sd1694657, 32'sd313417, -32'sd1067765, -32'sd2100605, -32'sd1209960, 32'sd752435, 32'sd2699689, 32'sd346518, 32'sd1119551, -32'sd1046397, -32'sd1871203, -32'sd2836588, -32'sd2671611, -32'sd2940077, -32'sd736068, -32'sd337053, -32'sd2419183, -32'sd4003530, -32'sd1530090, -32'sd727448, -32'sd1383822, -32'sd1613698, -32'sd465467, 32'sd2087530, -32'sd441875, -32'sd254584, 32'sd1914994, 32'sd632162, -32'sd1355902, 32'sd280476, -32'sd1974333, -32'sd2908730, -32'sd1776767, -32'sd1263868, 32'sd556461, 32'sd380635, 32'sd1737269, 32'sd73967, -32'sd1374205, -32'sd2999964, -32'sd2549972, -32'sd2429310, -32'sd2510867, -32'sd703440, -32'sd3069014, -32'sd3979650, -32'sd1919472, -32'sd433744, -32'sd1179991, 32'sd116560, -32'sd2266040, -32'sd1971605, -32'sd1417245, 32'sd621273, -32'sd124575, -32'sd1836836, -32'sd2121048, 32'sd278239, 32'sd948380, -32'sd1664898, 32'sd164155, 32'sd485046, -32'sd184871, 32'sd1495411, 32'sd1462100, -32'sd176984, -32'sd2309743, -32'sd1340604, -32'sd3724253, -32'sd1907673, -32'sd3607950, -32'sd1581036, -32'sd2691442, -32'sd2968342, -32'sd2815512, 32'sd951061, -32'sd2249355, 32'sd1072401, -32'sd1535152, 32'sd21716, -32'sd707135, 32'sd10250, 32'sd631114, 32'sd491069, -32'sd1693776, 32'sd897367, 32'sd492173, -32'sd298766, 32'sd674540, -32'sd198062, 32'sd522893, 32'sd3300305, 32'sd659438, -32'sd1262588, -32'sd3837007, -32'sd2649885, -32'sd1063525, -32'sd862159, -32'sd1605361, 32'sd982941, -32'sd424171, -32'sd102218, -32'sd1698309, 32'sd672115, -32'sd171718, 32'sd1612934, -32'sd1016187, 32'sd2615937, -32'sd1540248, 32'sd157578, 32'sd0, 32'sd950852, 32'sd927613, 32'sd49444, 32'sd1235932, 32'sd1570886, 32'sd943228, 32'sd1922783, 32'sd2951612, 32'sd3040303, 32'sd1101094, -32'sd963792, -32'sd1623951, -32'sd1600732, -32'sd1131449, 32'sd398245, 32'sd1433293, 32'sd659941, 32'sd257697, -32'sd1416115, 32'sd119843, -32'sd1680141, -32'sd1380808, -32'sd894370, 32'sd12971, -32'sd1326620, 32'sd133968, 32'sd700247, -32'sd395200, -32'sd478665, 32'sd229120, -32'sd1368038, -32'sd875017, 32'sd654214, 32'sd1765673, 32'sd2495440, 32'sd1199848, -32'sd267891, 32'sd1038148, -32'sd395211, -32'sd1074459, 32'sd1804762, 32'sd1365589, 32'sd426280, 32'sd958905, 32'sd330885, -32'sd283423, -32'sd1175257, -32'sd662942, 32'sd762018, -32'sd1378338, 32'sd1121944, -32'sd528177, -32'sd976239, 32'sd479172, 32'sd735393, 32'sd776883, -32'sd1146681, -32'sd1480306, -32'sd1151233, 32'sd1611208, -32'sd513214, 32'sd1225465, 32'sd1324754, -32'sd371241, 32'sd371135, -32'sd2155848, -32'sd1329763, 32'sd1167037, 32'sd1199945, 32'sd454933, 32'sd378779, 32'sd284750, 32'sd19798, 32'sd34570, -32'sd354901, -32'sd1523098, -32'sd425708, -32'sd594767, -32'sd1093378, 32'sd1252738, -32'sd919125, 32'sd481410, 32'sd1829271, 32'sd0, 32'sd50352, 32'sd1664893, 32'sd20978, -32'sd963531, 32'sd699469, -32'sd828029, 32'sd1143168, -32'sd1125967, -32'sd2060411, 32'sd626395, 32'sd404642, 32'sd2129680, 32'sd1339709, 32'sd2131153, 32'sd2475814, 32'sd587337, -32'sd1922200, -32'sd2002176, -32'sd2058842, -32'sd755927, -32'sd846019, -32'sd851674, -32'sd1619671, 32'sd121234, -32'sd2409135, -32'sd1664766, 32'sd389890, 32'sd545821, -32'sd1146525, 32'sd142652, 32'sd2351741, -32'sd886138, -32'sd1509854, -32'sd598990, 32'sd337068, 32'sd732379, 32'sd317878, -32'sd261097, 32'sd1630244, 32'sd48350, 32'sd566283, 32'sd89780, 32'sd1564006, 32'sd58502, -32'sd1039385, -32'sd1942561, -32'sd1129935, -32'sd1279860, 32'sd97677, -32'sd543825, -32'sd1182703, 32'sd666882, 32'sd492116, -32'sd296315, 32'sd96575, -32'sd495435, 32'sd67043, 32'sd98682, -32'sd1260570, -32'sd535703, -32'sd533415, 32'sd1446802, 32'sd665933, 32'sd1586364, -32'sd184461, 32'sd1277705, 32'sd1096209, 32'sd2047770, -32'sd220366, 32'sd614238, 32'sd259904, -32'sd1378181, 32'sd513265, 32'sd762005, -32'sd882215, 32'sd306197, 32'sd239102, -32'sd414061, -32'sd546367, -32'sd110497, 32'sd980474, -32'sd652874, 32'sd306240, 32'sd0, 32'sd387265, 32'sd509327, -32'sd760195, -32'sd1425410, -32'sd1354379, -32'sd751958, 32'sd526956, -32'sd770976, -32'sd1090823, -32'sd230331, 32'sd1951496, 32'sd2943082, -32'sd411549, 32'sd164876, 32'sd389164, 32'sd1216459, -32'sd188257, 32'sd115994, 32'sd1258059, 32'sd390707, -32'sd1216673, 32'sd446676, 32'sd1003793, 32'sd1103040, 32'sd682560, 32'sd160579, 32'sd0, 32'sd0, 32'sd0, -32'sd1236489, -32'sd703465, -32'sd728752, 32'sd269065, -32'sd966125, -32'sd1172244, -32'sd1697342, -32'sd1904083, -32'sd647355, 32'sd261749, -32'sd146535, -32'sd1089184, -32'sd526948, 32'sd782946, -32'sd203143, -32'sd442209, 32'sd159556, 32'sd108784, 32'sd1318244, -32'sd318571, -32'sd1506473, 32'sd2803, -32'sd522713, -32'sd98694, 32'sd645287, 32'sd0, 32'sd0, 32'sd0, 32'sd584111, 32'sd724260, 32'sd1245962, 32'sd660921, 32'sd1663657, 32'sd1517649, -32'sd1087265, 32'sd305355, -32'sd1461449, 32'sd1522952, -32'sd598128, 32'sd17453, 32'sd1748169, 32'sd312919, 32'sd506977, -32'sd363565, 32'sd298328, -32'sd490382, 32'sd65242, 32'sd1236279, 32'sd570762, -32'sd39310, 32'sd2110938, -32'sd1742274, -32'sd109019, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd773699, -32'sd1235671, 32'sd69999, -32'sd250110, -32'sd264422, 32'sd245506, -32'sd873885, 32'sd976334, -32'sd1370530, -32'sd578611, 32'sd777239, -32'sd396937, 32'sd805276, 32'sd1195527, 32'sd1006714, 32'sd1354702, 32'sd1994243, 32'sd1443095, -32'sd710290, 32'sd1099560, -32'sd1098651, -32'sd567659, 32'sd6658, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd847061, -32'sd503990, 32'sd888482, -32'sd616279, -32'sd306230, -32'sd1607222, 32'sd623720, -32'sd757466, 32'sd1465244, 32'sd88314, 32'sd611035, -32'sd1230385, 32'sd1127205, 32'sd509390, -32'sd819174, -32'sd3492, 32'sd115613, 32'sd402723, -32'sd475759, -32'sd341737, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd494123, 32'sd102830, -32'sd445053, 32'sd673182, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd172881, 32'sd487389, -32'sd867250, -32'sd738529, 32'sd316385, 32'sd146471, -32'sd105718, 32'sd239017, 32'sd1341114, -32'sd821449, 32'sd731645, -32'sd162592, -32'sd1746871, 32'sd1222669, 32'sd738552, 32'sd65185, 32'sd645110, 32'sd691949, -32'sd629988, 32'sd222891, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd108068, 32'sd757719, -32'sd708952, 32'sd1498428, 32'sd1399288, 32'sd727513, 32'sd1387176, -32'sd266546, -32'sd70231, 32'sd369844, 32'sd201434, -32'sd882834, -32'sd2377184, 32'sd303624, -32'sd1381592, -32'sd1226411, -32'sd282073, 32'sd357808, -32'sd1000661, -32'sd860035, 32'sd97422, 32'sd1189499, 32'sd396340, -32'sd226392, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1236172, -32'sd645745, 32'sd362699, 32'sd55982, -32'sd138906, 32'sd884704, 32'sd1143519, 32'sd599713, 32'sd2168136, 32'sd438729, 32'sd563327, -32'sd1939709, 32'sd438017, 32'sd637371, 32'sd839511, -32'sd197674, -32'sd118803, 32'sd521314, -32'sd165856, 32'sd1510032, 32'sd1105185, -32'sd12568, -32'sd1187142, 32'sd1178366, 32'sd1277017, 32'sd0, 32'sd0, -32'sd38085, 32'sd1044794, -32'sd104406, 32'sd48238, -32'sd399903, -32'sd1761591, -32'sd936725, -32'sd675256, -32'sd3433974, -32'sd1588874, 32'sd677664, 32'sd392886, 32'sd1302167, -32'sd191738, -32'sd689070, -32'sd969706, -32'sd802556, -32'sd1988640, -32'sd1164774, -32'sd2169650, -32'sd1686292, 32'sd352686, 32'sd1823135, -32'sd217180, -32'sd479791, 32'sd1356930, -32'sd292940, 32'sd0, -32'sd392563, 32'sd835229, -32'sd688364, -32'sd437038, -32'sd224587, 32'sd423869, 32'sd227093, -32'sd210163, -32'sd1264367, -32'sd133009, -32'sd2727136, -32'sd1271399, 32'sd735609, 32'sd1722056, 32'sd352446, 32'sd1008150, -32'sd2898316, -32'sd3883188, -32'sd3084120, -32'sd725441, 32'sd464044, -32'sd1429630, 32'sd621054, -32'sd851512, -32'sd519278, -32'sd396345, -32'sd884716, 32'sd0, 32'sd204365, -32'sd657273, -32'sd1207988, -32'sd243564, 32'sd943807, -32'sd878043, 32'sd153723, -32'sd1781458, 32'sd3132657, 32'sd2094127, -32'sd560172, 32'sd496647, 32'sd1533034, 32'sd1394871, 32'sd371873, -32'sd348159, 32'sd41083, 32'sd501269, 32'sd883021, 32'sd2190751, 32'sd2549576, 32'sd2935930, 32'sd103907, 32'sd740116, -32'sd639376, 32'sd265758, 32'sd210960, 32'sd581091, 32'sd388927, -32'sd96402, 32'sd1713293, -32'sd339340, 32'sd124327, -32'sd283366, 32'sd1420583, 32'sd1394548, 32'sd501664, 32'sd2500474, 32'sd1509583, 32'sd555234, 32'sd538359, 32'sd803641, -32'sd1734063, 32'sd1327536, 32'sd1536390, 32'sd1175297, 32'sd1602286, 32'sd905487, 32'sd1490091, 32'sd45575, -32'sd1853397, -32'sd25538, -32'sd89387, -32'sd857670, 32'sd519398, -32'sd640392, 32'sd952543, -32'sd469861, 32'sd1984603, 32'sd274580, 32'sd1033813, -32'sd1364655, 32'sd1984240, 32'sd188639, 32'sd2278527, 32'sd3774218, 32'sd3570609, 32'sd3625665, 32'sd4209717, 32'sd2833793, 32'sd3022587, 32'sd2936782, 32'sd1370104, 32'sd2066037, 32'sd525156, 32'sd1290599, -32'sd343550, 32'sd2244339, 32'sd1821415, 32'sd386264, 32'sd333247, -32'sd376175, 32'sd997436, 32'sd1047091, 32'sd100749, 32'sd119422, -32'sd2113754, -32'sd18296, -32'sd1134306, 32'sd706728, 32'sd2339363, 32'sd2058095, 32'sd2233755, 32'sd2267248, 32'sd2373285, 32'sd2994957, 32'sd2478726, 32'sd3645245, 32'sd2115355, 32'sd1753472, 32'sd1408166, 32'sd757767, -32'sd2217620, -32'sd527394, 32'sd736049, 32'sd1225528, 32'sd2096887, 32'sd1184123, 32'sd90899, 32'sd191328, 32'sd634644, 32'sd357673, -32'sd90096, -32'sd1630004, 32'sd378864, -32'sd726571, -32'sd423597, 32'sd1014583, 32'sd2285318, 32'sd2745040, 32'sd1444792, 32'sd1286367, -32'sd823142, -32'sd196297, -32'sd19023, -32'sd1213425, -32'sd627343, 32'sd17556, -32'sd2049409, -32'sd2377717, -32'sd653263, -32'sd889179, -32'sd1129213, 32'sd2267082, 32'sd1455195, 32'sd1416613, 32'sd421278, 32'sd484310, -32'sd133678, -32'sd405542, -32'sd1340397, -32'sd655228, 32'sd324378, 32'sd712821, -32'sd276505, 32'sd148329, 32'sd141000, 32'sd3663285, -32'sd274178, -32'sd2103864, -32'sd2071589, -32'sd2464410, -32'sd4046103, -32'sd4526607, -32'sd1973898, -32'sd1607290, -32'sd3140274, -32'sd689469, -32'sd2520370, -32'sd1535943, 32'sd1118074, 32'sd2269608, 32'sd522282, 32'sd257962, -32'sd1361098, 32'sd1100393, -32'sd1526237, 32'sd1044886, -32'sd1323543, 32'sd452250, 32'sd452705, 32'sd335500, 32'sd131695, -32'sd1596516, -32'sd1813839, -32'sd75775, -32'sd3553067, -32'sd5178600, -32'sd4018461, -32'sd3194308, -32'sd3643663, -32'sd3049509, -32'sd168459, -32'sd402016, 32'sd118930, -32'sd374568, 32'sd196337, -32'sd492110, -32'sd891159, -32'sd2100380, -32'sd651223, -32'sd1171711, 32'sd1607713, 32'sd738870, 32'sd944934, -32'sd73063, -32'sd957696, -32'sd953533, -32'sd629648, -32'sd1133979, -32'sd1690929, -32'sd3088135, -32'sd4436067, -32'sd4315938, -32'sd5598590, -32'sd3743668, -32'sd1076660, -32'sd1972026, -32'sd2490846, 32'sd43355, -32'sd1863759, -32'sd540831, -32'sd1062175, 32'sd1076505, -32'sd2040737, -32'sd3817640, -32'sd1418167, 32'sd926018, -32'sd213755, 32'sd2218988, 32'sd655677, -32'sd31375, 32'sd1155362, 32'sd151963, -32'sd819677, 32'sd297105, -32'sd171777, -32'sd2093654, -32'sd3763844, -32'sd3942259, -32'sd4220487, -32'sd3007618, -32'sd4474636, -32'sd421944, -32'sd1344275, 32'sd471751, -32'sd97347, 32'sd517008, 32'sd746144, 32'sd281042, 32'sd2940454, 32'sd1869194, -32'sd60498, -32'sd1156088, 32'sd1351961, 32'sd1665059, -32'sd145274, -32'sd308709, 32'sd50252, -32'sd184835, 32'sd387502, -32'sd648953, -32'sd249924, -32'sd1289951, -32'sd2522062, -32'sd2871004, -32'sd4373123, -32'sd3119062, -32'sd2843238, -32'sd1154018, -32'sd1205575, 32'sd749395, 32'sd1370892, 32'sd683696, 32'sd2187881, -32'sd49465, 32'sd2750634, 32'sd1234868, 32'sd1939080, -32'sd627806, 32'sd250960, -32'sd649774, -32'sd421241, 32'sd903777, 32'sd205195, 32'sd912858, -32'sd1948927, 32'sd208669, -32'sd800653, 32'sd1084478, -32'sd834019, -32'sd697553, 32'sd333549, -32'sd1640709, -32'sd1673848, -32'sd215587, 32'sd392891, 32'sd1290840, 32'sd934760, -32'sd873216, 32'sd1685751, 32'sd1300321, 32'sd263888, 32'sd3093613, 32'sd1369094, 32'sd2567753, 32'sd1746739, 32'sd1582523, 32'sd1630494, 32'sd160840, 32'sd1016394, 32'sd307477, 32'sd1630940, 32'sd57038, -32'sd18224, 32'sd897332, -32'sd1195336, 32'sd0, 32'sd655140, -32'sd673481, 32'sd321896, 32'sd958124, -32'sd1087613, -32'sd1618306, -32'sd117029, 32'sd546464, 32'sd1058770, 32'sd431475, 32'sd240627, -32'sd135668, 32'sd499594, 32'sd2930377, 32'sd2507349, 32'sd1504195, 32'sd375055, -32'sd291124, 32'sd1372112, 32'sd344360, -32'sd473343, -32'sd2046630, -32'sd2757594, 32'sd239563, -32'sd1134376, -32'sd1241734, 32'sd1040640, 32'sd121477, 32'sd1352820, -32'sd595610, -32'sd1547528, -32'sd574461, -32'sd720646, 32'sd459256, -32'sd531969, -32'sd254143, 32'sd137502, 32'sd1115106, -32'sd284240, 32'sd946580, 32'sd1404926, 32'sd1766155, 32'sd2803440, 32'sd831145, 32'sd168367, -32'sd727954, 32'sd1451362, 32'sd1298017, -32'sd2396725, -32'sd2979275, 32'sd207962, -32'sd1645047, -32'sd559335, -32'sd1802539, 32'sd1064520, -32'sd384152, -32'sd328455, 32'sd409873, 32'sd357056, 32'sd910345, 32'sd115671, 32'sd513163, 32'sd695356, 32'sd363620, -32'sd346987, -32'sd1339263, 32'sd351078, -32'sd188227, 32'sd2846108, 32'sd1335487, 32'sd205469, -32'sd235098, -32'sd1446847, -32'sd2834894, -32'sd167501, -32'sd582939, -32'sd2284053, -32'sd621465, -32'sd358886, 32'sd505469, -32'sd1204961, -32'sd1080265, 32'sd642880, 32'sd0, -32'sd1082667, 32'sd1296330, 32'sd1700965, 32'sd825135, 32'sd1096329, 32'sd1228993, 32'sd1351290, 32'sd1582741, 32'sd563908, 32'sd114061, -32'sd768150, 32'sd1773812, 32'sd495114, 32'sd1442991, 32'sd1708840, -32'sd284156, -32'sd2375326, -32'sd1490219, -32'sd1730845, -32'sd1283485, -32'sd122197, -32'sd148551, -32'sd99940, -32'sd606840, -32'sd236798, -32'sd908013, -32'sd591227, 32'sd569554, 32'sd132625, 32'sd878567, -32'sd632416, 32'sd1319100, 32'sd147203, 32'sd1549257, 32'sd661060, -32'sd696654, -32'sd796887, 32'sd1415789, 32'sd1000056, 32'sd2821914, 32'sd539278, -32'sd296804, -32'sd185730, -32'sd987097, -32'sd1611802, -32'sd537125, 32'sd1097307, -32'sd692533, 32'sd231239, 32'sd417254, 32'sd815507, 32'sd825016, -32'sd541710, -32'sd443834, 32'sd263978, -32'sd72246, -32'sd596835, 32'sd56850, -32'sd1208515, 32'sd1771815, -32'sd118917, -32'sd98421, -32'sd1348156, 32'sd973835, 32'sd101638, 32'sd2644636, 32'sd2466482, 32'sd629551, -32'sd1389, -32'sd847598, 32'sd178031, -32'sd456794, 32'sd730816, 32'sd467081, -32'sd862446, -32'sd1026819, -32'sd678692, 32'sd1447468, -32'sd337903, 32'sd551513, -32'sd1675763, -32'sd81726, -32'sd10677, 32'sd0, 32'sd541365, -32'sd1602731, -32'sd2648512, 32'sd893305, 32'sd138562, 32'sd1438007, 32'sd987074, -32'sd213157, 32'sd283040, 32'sd37044, 32'sd784857, 32'sd275437, -32'sd1019390, 32'sd1511482, 32'sd1238579, 32'sd1751761, 32'sd905225, 32'sd1230415, -32'sd1064129, -32'sd1694717, 32'sd41652, 32'sd816378, 32'sd1314718, 32'sd1116064, -32'sd1070809, 32'sd1080425, 32'sd0, 32'sd0, 32'sd0, 32'sd1572592, -32'sd856035, -32'sd672333, 32'sd352998, 32'sd920629, -32'sd44850, -32'sd190870, 32'sd1266210, 32'sd804951, -32'sd730026, -32'sd1291093, 32'sd689455, 32'sd948561, 32'sd795266, -32'sd234770, -32'sd60414, -32'sd1122548, -32'sd3060423, 32'sd487992, -32'sd104436, 32'sd914661, -32'sd728447, 32'sd767495, -32'sd75752, 32'sd167789, 32'sd0, 32'sd0, 32'sd0, 32'sd799382, 32'sd1756144, 32'sd1469088, 32'sd700988, 32'sd1083150, 32'sd1435474, 32'sd575200, 32'sd1865121, 32'sd2296086, -32'sd756776, 32'sd1134801, -32'sd398649, -32'sd535564, 32'sd2177298, 32'sd255724, 32'sd540172, -32'sd2465376, 32'sd781776, -32'sd78968, -32'sd117971, 32'sd278414, 32'sd738969, 32'sd489150, 32'sd1220409, -32'sd552938, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd84638, -32'sd599486, -32'sd1750880, 32'sd214448, 32'sd1563203, -32'sd220012, 32'sd1535481, -32'sd1821553, -32'sd2328690, -32'sd1355274, 32'sd1179498, 32'sd118433, 32'sd851619, -32'sd2885918, -32'sd732812, -32'sd873365, -32'sd738435, -32'sd1593664, -32'sd1671921, -32'sd308961, -32'sd710798, -32'sd1067807, -32'sd579850, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd5431, -32'sd627853, 32'sd841566, -32'sd799569, 32'sd340692, -32'sd465741, 32'sd1448684, 32'sd685431, -32'sd1106513, 32'sd611749, 32'sd2527878, 32'sd1507826, 32'sd1462994, 32'sd1572135, 32'sd1094783, -32'sd1537343, -32'sd212418, 32'sd508455, -32'sd881226, 32'sd191562, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1986169, 32'sd1317338, 32'sd2392023, 32'sd2372322, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd307545, 32'sd747314, 32'sd929677, -32'sd781083, -32'sd903347, 32'sd1860912, 32'sd119172, 32'sd1836978, 32'sd1293763, 32'sd227190, -32'sd868324, 32'sd945502, 32'sd1375610, 32'sd1075906, -32'sd431360, 32'sd1028753, -32'sd101230, 32'sd740357, -32'sd345867, 32'sd806432, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2174200, -32'sd1018287, 32'sd661208, -32'sd361094, 32'sd1966359, 32'sd899848, 32'sd912732, 32'sd254133, 32'sd2772038, 32'sd369717, 32'sd980131, -32'sd1524960, 32'sd977575, -32'sd494818, 32'sd1597175, 32'sd2696458, -32'sd389882, 32'sd1512565, -32'sd619732, 32'sd1641060, -32'sd689715, 32'sd390962, 32'sd1187662, 32'sd2817107, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2600666, 32'sd918691, 32'sd273163, -32'sd682612, 32'sd62569, -32'sd1432571, -32'sd345366, -32'sd848715, 32'sd767505, 32'sd1586501, 32'sd587464, 32'sd1376783, 32'sd1074977, 32'sd2406080, 32'sd2367133, 32'sd1306627, -32'sd1552026, -32'sd1390330, -32'sd1651782, 32'sd1123787, 32'sd2222811, -32'sd73441, -32'sd352536, -32'sd559916, -32'sd1397270, 32'sd0, 32'sd0, 32'sd923178, 32'sd605330, -32'sd105104, -32'sd1698007, -32'sd1406738, -32'sd783896, -32'sd120238, -32'sd363168, -32'sd909792, 32'sd1141091, -32'sd340616, 32'sd424413, 32'sd1943242, 32'sd672790, -32'sd1209316, -32'sd1669068, -32'sd250196, -32'sd643003, -32'sd631703, -32'sd2108658, -32'sd1237289, 32'sd1320932, 32'sd645384, -32'sd1748583, -32'sd515130, 32'sd1600978, -32'sd684432, 32'sd0, 32'sd1248767, 32'sd575071, 32'sd450110, 32'sd645653, 32'sd8670, 32'sd416880, -32'sd2091403, 32'sd1256822, 32'sd1832849, 32'sd286236, 32'sd3108447, 32'sd1416236, 32'sd1874867, -32'sd1275369, -32'sd1745045, -32'sd2642179, -32'sd2546924, -32'sd1631322, -32'sd1317519, -32'sd814926, 32'sd156213, -32'sd326930, -32'sd198420, 32'sd703950, 32'sd2468337, 32'sd1974722, 32'sd1149280, 32'sd0, 32'sd1141111, -32'sd106829, -32'sd264291, -32'sd894162, -32'sd657524, -32'sd2662424, -32'sd613479, -32'sd340099, -32'sd671281, 32'sd1934516, 32'sd2317053, 32'sd2490114, 32'sd163488, 32'sd888439, -32'sd1147720, -32'sd1962632, -32'sd122307, -32'sd2444542, -32'sd940193, 32'sd87936, 32'sd1902952, 32'sd1314638, -32'sd1329345, 32'sd856933, 32'sd2555059, 32'sd808320, -32'sd310004, 32'sd1987623, 32'sd875639, 32'sd478207, -32'sd601403, 32'sd228793, -32'sd565062, -32'sd1524931, -32'sd2077393, -32'sd1418421, -32'sd969551, 32'sd220948, 32'sd1430654, 32'sd2052077, 32'sd957689, -32'sd87115, 32'sd468048, 32'sd1751386, 32'sd1232734, 32'sd1916227, 32'sd1673775, 32'sd2030515, 32'sd1927895, 32'sd1393311, 32'sd1305852, 32'sd28293, 32'sd508560, 32'sd1673579, -32'sd1143786, 32'sd336984, 32'sd378814, 32'sd824954, -32'sd102243, 32'sd1743777, -32'sd983552, -32'sd54120, -32'sd1098513, -32'sd1238946, 32'sd513116, 32'sd333607, 32'sd1067357, 32'sd1775467, 32'sd2742414, 32'sd1603901, 32'sd1619763, 32'sd501761, 32'sd2903026, 32'sd2112286, 32'sd4131656, 32'sd4317034, 32'sd3278767, 32'sd2158160, 32'sd3059962, 32'sd2564642, 32'sd1865179, 32'sd1463138, -32'sd662635, 32'sd1684789, 32'sd378382, 32'sd1607969, 32'sd1959788, 32'sd2083114, 32'sd562649, -32'sd796230, -32'sd2055838, -32'sd2109730, -32'sd720544, -32'sd1275475, 32'sd1132270, 32'sd1057890, 32'sd2939993, 32'sd1734962, -32'sd780527, 32'sd3205924, -32'sd601702, 32'sd1848753, 32'sd1986878, 32'sd1662676, 32'sd966345, 32'sd1689910, 32'sd232413, 32'sd1810294, -32'sd959331, 32'sd604634, 32'sd1370289, 32'sd1018227, -32'sd485139, 32'sd1750112, 32'sd662865, 32'sd536700, 32'sd215933, -32'sd161962, -32'sd862562, -32'sd886933, -32'sd992901, 32'sd2107665, 32'sd178812, 32'sd1888001, 32'sd1579817, -32'sd967683, 32'sd1255647, 32'sd1657895, -32'sd1255431, 32'sd254717, -32'sd1162859, 32'sd802211, 32'sd1070848, -32'sd540291, -32'sd434367, -32'sd909777, -32'sd1379831, -32'sd128571, 32'sd1207325, 32'sd1312812, 32'sd530956, -32'sd424058, 32'sd1012787, -32'sd93878, -32'sd1951132, 32'sd526238, -32'sd933661, -32'sd971901, 32'sd599653, 32'sd466658, 32'sd523566, 32'sd2107203, -32'sd31821, -32'sd53735, 32'sd101973, -32'sd1387294, -32'sd2016281, -32'sd2315606, -32'sd2909052, -32'sd2649841, 32'sd727460, -32'sd1632607, -32'sd613364, -32'sd1660467, -32'sd1209535, 32'sd150156, 32'sd1233501, 32'sd1476724, 32'sd1051437, -32'sd670428, 32'sd187047, -32'sd469867, -32'sd818216, -32'sd1681139, -32'sd1235300, -32'sd987646, 32'sd117487, -32'sd1445676, -32'sd25468, 32'sd1225823, -32'sd1009219, -32'sd1655453, -32'sd767026, -32'sd1707240, -32'sd811224, -32'sd2284536, -32'sd2784711, -32'sd862632, 32'sd261720, 32'sd1218487, -32'sd707431, -32'sd128527, -32'sd1421526, -32'sd2206261, 32'sd1060256, 32'sd1011002, 32'sd930096, 32'sd718014, 32'sd1123912, -32'sd2363708, 32'sd1376426, -32'sd183560, 32'sd99575, -32'sd2431223, -32'sd854883, -32'sd1010732, -32'sd2206027, 32'sd771118, 32'sd752483, 32'sd345802, -32'sd414087, 32'sd215916, -32'sd80798, -32'sd435468, -32'sd2000972, -32'sd2211192, -32'sd2330011, -32'sd997718, -32'sd1857991, -32'sd3035899, -32'sd1142497, 32'sd661569, 32'sd658283, 32'sd2320049, 32'sd1016013, -32'sd1350068, -32'sd945757, -32'sd1547349, 32'sd908982, -32'sd3023918, -32'sd494742, -32'sd2720283, -32'sd2556256, -32'sd1722071, -32'sd1612195, 32'sd1729422, 32'sd3103555, 32'sd1580045, 32'sd608740, 32'sd1709436, 32'sd727493, -32'sd1453238, 32'sd290228, -32'sd2928033, -32'sd1487157, -32'sd1940055, -32'sd997863, -32'sd2060645, 32'sd539174, 32'sd268779, 32'sd1449603, -32'sd23640, 32'sd98888, -32'sd665132, -32'sd1485537, 32'sd100621, -32'sd1419116, -32'sd3409135, -32'sd2205133, -32'sd1754027, -32'sd2921707, -32'sd1027132, 32'sd680071, 32'sd1881162, 32'sd2999810, 32'sd1500877, -32'sd1397598, -32'sd604127, -32'sd167578, -32'sd266277, -32'sd2333500, -32'sd1298267, -32'sd489622, -32'sd1756699, -32'sd2495045, -32'sd1466758, 32'sd1456867, 32'sd1630504, 32'sd1264608, 32'sd616477, 32'sd385119, 32'sd127236, -32'sd1825647, 32'sd1248231, -32'sd1187159, -32'sd1159197, -32'sd1992332, -32'sd2631313, -32'sd2717375, 32'sd888168, 32'sd3190130, 32'sd2642782, 32'sd3119425, 32'sd657991, -32'sd1892214, -32'sd1933500, -32'sd437894, -32'sd2519873, -32'sd2399406, -32'sd2027290, 32'sd61577, 32'sd2214006, 32'sd472034, 32'sd1027350, 32'sd2014922, 32'sd1239809, 32'sd1559668, 32'sd0, 32'sd382272, -32'sd200714, -32'sd1120385, -32'sd312935, 32'sd175249, 32'sd383100, 32'sd1098402, -32'sd1247347, -32'sd922249, 32'sd2268543, 32'sd5401044, 32'sd5676586, 32'sd2036125, -32'sd1630532, -32'sd2629687, -32'sd2177326, -32'sd538503, -32'sd997368, -32'sd1496134, 32'sd573470, 32'sd1088760, 32'sd3148272, 32'sd1581590, 32'sd79041, 32'sd2474802, 32'sd1212257, 32'sd418214, 32'sd99019, -32'sd233207, -32'sd244878, 32'sd397608, -32'sd666492, -32'sd2144850, 32'sd389208, 32'sd1370544, 32'sd735819, 32'sd1912878, 32'sd2552020, 32'sd3835420, 32'sd4260297, -32'sd502670, -32'sd4395721, -32'sd5669058, -32'sd2128693, 32'sd636515, -32'sd1651294, -32'sd225547, 32'sd877808, -32'sd408775, 32'sd1312689, 32'sd200472, 32'sd1919756, 32'sd2023782, 32'sd3260577, 32'sd966125, 32'sd142196, 32'sd737700, -32'sd753784, 32'sd218999, -32'sd1662244, -32'sd1566929, -32'sd574875, -32'sd4253, 32'sd1058336, 32'sd627501, 32'sd3453896, 32'sd4505753, 32'sd2913913, -32'sd2002031, -32'sd3759026, -32'sd3868328, -32'sd1135672, -32'sd1057808, -32'sd1268615, -32'sd33967, 32'sd1461929, -32'sd188967, -32'sd1523721, -32'sd23213, 32'sd972564, 32'sd2450495, 32'sd2527117, -32'sd120650, 32'sd0, -32'sd64166, 32'sd211415, -32'sd266208, -32'sd2113448, 32'sd1005809, 32'sd43327, 32'sd119956, 32'sd1548409, 32'sd631531, 32'sd3288576, 32'sd4360879, 32'sd33741, -32'sd3333706, -32'sd4834653, -32'sd2474076, -32'sd389225, -32'sd791511, 32'sd237531, -32'sd174815, 32'sd186428, -32'sd1449998, -32'sd185843, -32'sd379789, 32'sd156344, 32'sd976353, 32'sd721365, 32'sd2475763, 32'sd678790, 32'sd1036468, 32'sd1548888, 32'sd1429550, 32'sd1607315, 32'sd596234, -32'sd350054, 32'sd1326531, 32'sd591574, 32'sd3696808, 32'sd2161640, 32'sd867730, 32'sd1320673, -32'sd1473741, -32'sd2351119, -32'sd3164709, -32'sd1312454, -32'sd76567, -32'sd2247080, -32'sd1044073, 32'sd1076351, 32'sd972532, 32'sd61487, 32'sd98682, 32'sd479289, 32'sd1885920, -32'sd598833, 32'sd1430506, -32'sd627946, -32'sd828406, 32'sd152150, -32'sd950990, -32'sd991315, 32'sd1443458, -32'sd171211, 32'sd33096, 32'sd2469721, 32'sd2885963, 32'sd506333, -32'sd971502, -32'sd2171212, -32'sd453576, -32'sd2029167, -32'sd1116166, -32'sd3124964, -32'sd1306878, 32'sd185417, -32'sd1143350, 32'sd1266732, 32'sd314818, 32'sd320828, -32'sd593713, -32'sd206365, 32'sd1650345, -32'sd172071, 32'sd1109539, 32'sd0, -32'sd836878, 32'sd429037, -32'sd257657, -32'sd776049, 32'sd1165406, 32'sd2466304, -32'sd863243, 32'sd178817, 32'sd1430570, 32'sd2105282, 32'sd730503, 32'sd251428, -32'sd1441149, 32'sd186755, 32'sd631239, 32'sd189609, -32'sd375689, -32'sd1915373, 32'sd2140013, -32'sd604905, -32'sd1966607, -32'sd1554310, -32'sd2474275, 32'sd1162714, 32'sd727458, 32'sd109792, 32'sd0, 32'sd0, 32'sd0, 32'sd53310, -32'sd1657508, -32'sd2340239, -32'sd1937410, -32'sd211173, -32'sd216873, 32'sd699465, -32'sd541587, 32'sd319744, 32'sd1244471, 32'sd3387142, 32'sd2037905, 32'sd829980, -32'sd1251524, 32'sd483296, -32'sd1463149, 32'sd592221, 32'sd929302, -32'sd1954298, -32'sd167002, 32'sd165716, -32'sd136928, 32'sd920753, 32'sd384539, 32'sd568165, 32'sd0, 32'sd0, 32'sd0, -32'sd95553, 32'sd868353, 32'sd1804494, -32'sd1072392, -32'sd1723283, 32'sd751481, 32'sd520124, 32'sd864132, -32'sd1483657, 32'sd316545, 32'sd141834, 32'sd927620, -32'sd1194456, -32'sd1126453, -32'sd1480502, 32'sd1011892, -32'sd774417, -32'sd3163234, -32'sd2238167, -32'sd1859197, -32'sd1178989, 32'sd651645, -32'sd621066, 32'sd154782, 32'sd364825, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2197561, -32'sd77905, 32'sd1631302, 32'sd273930, 32'sd405232, 32'sd903693, -32'sd493987, 32'sd1060230, 32'sd739581, -32'sd1769327, -32'sd643121, -32'sd1660078, -32'sd1412649, 32'sd444644, 32'sd1268131, -32'sd916100, 32'sd1441009, 32'sd564832, 32'sd135218, 32'sd1282266, -32'sd921219, 32'sd1241531, 32'sd1573671, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2132439, 32'sd1283940, 32'sd1378930, 32'sd1089966, 32'sd86246, -32'sd1418491, 32'sd553178, 32'sd956313, -32'sd747442, 32'sd1820028, 32'sd2230582, 32'sd1447046, 32'sd1560553, 32'sd726487, 32'sd280232, 32'sd2309043, 32'sd1527940, 32'sd923463, -32'sd1061787, 32'sd1055625, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd92702, 32'sd250098, 32'sd272310, 32'sd1719339, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd512513, -32'sd676056, 32'sd485169, 32'sd893006, -32'sd236803, -32'sd290248, 32'sd2345205, 32'sd2240299, 32'sd1042631, 32'sd413677, -32'sd1088412, 32'sd196829, -32'sd626943, -32'sd203606, -32'sd609428, -32'sd183845, 32'sd1755114, 32'sd666051, 32'sd1460888, 32'sd745849, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1478842, 32'sd1204325, 32'sd446828, 32'sd82277, 32'sd1895910, 32'sd1562515, 32'sd1707137, 32'sd1395656, 32'sd81300, 32'sd899134, -32'sd605614, -32'sd1763282, -32'sd664555, -32'sd825033, 32'sd55878, 32'sd1154192, 32'sd1638075, 32'sd1795103, 32'sd755968, 32'sd2124717, 32'sd1596918, -32'sd201856, 32'sd674134, 32'sd554238, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd170244, 32'sd737034, 32'sd1214850, 32'sd747394, 32'sd1194384, -32'sd1150759, -32'sd170924, 32'sd514251, -32'sd1977066, -32'sd1640839, -32'sd248413, -32'sd2495894, -32'sd507714, -32'sd1904208, -32'sd257104, -32'sd138651, 32'sd1893757, 32'sd1466563, 32'sd1301934, 32'sd1428012, -32'sd95626, -32'sd1022419, 32'sd51382, -32'sd2568820, 32'sd1266557, 32'sd0, 32'sd0, -32'sd50066, 32'sd160915, 32'sd412930, 32'sd86189, -32'sd640265, -32'sd1222428, -32'sd1677655, 32'sd286944, -32'sd2220317, -32'sd2085439, 32'sd1959968, -32'sd892617, 32'sd927154, -32'sd963424, 32'sd808965, -32'sd46518, -32'sd1537358, -32'sd1226078, -32'sd2133379, -32'sd1775793, 32'sd494153, -32'sd442934, -32'sd10245, -32'sd674205, 32'sd311102, 32'sd1264188, -32'sd749243, 32'sd0, 32'sd864965, -32'sd1199674, -32'sd1723963, 32'sd77822, 32'sd301014, -32'sd2079618, 32'sd420834, -32'sd2248680, -32'sd2656341, -32'sd2617917, -32'sd1930412, -32'sd2658177, -32'sd1844321, -32'sd2987166, -32'sd1978143, -32'sd1778057, -32'sd2037231, -32'sd494737, -32'sd1542115, 32'sd1541249, -32'sd676839, 32'sd546156, 32'sd881132, 32'sd934496, -32'sd406035, -32'sd957915, -32'sd647180, 32'sd0, 32'sd686512, 32'sd928937, 32'sd1005142, 32'sd1064835, 32'sd421652, 32'sd2080383, 32'sd773667, -32'sd58538, -32'sd2013773, -32'sd3762838, -32'sd3378908, -32'sd3911573, -32'sd1889273, -32'sd869731, -32'sd3124375, -32'sd1958550, 32'sd677094, 32'sd59541, 32'sd1237259, 32'sd111757, 32'sd928823, 32'sd1092307, -32'sd1040433, -32'sd538491, 32'sd1551272, 32'sd1487916, -32'sd89168, 32'sd592098, 32'sd294577, -32'sd2124139, 32'sd467269, 32'sd1064428, -32'sd454044, -32'sd1100772, 32'sd1017107, 32'sd1513261, -32'sd2337902, -32'sd2998207, -32'sd1820908, -32'sd2084421, -32'sd1917721, -32'sd739330, 32'sd2244498, 32'sd1312145, -32'sd288917, 32'sd1165151, 32'sd1352794, 32'sd945839, 32'sd1981396, 32'sd2427946, 32'sd1524723, 32'sd289360, 32'sd166413, 32'sd1798412, 32'sd664183, 32'sd806399, -32'sd1298963, -32'sd1311387, -32'sd2187130, -32'sd816258, -32'sd1108424, -32'sd2305964, -32'sd2596885, -32'sd1426663, -32'sd2178575, -32'sd1718149, -32'sd1717484, -32'sd2273257, 32'sd247927, -32'sd300030, -32'sd284473, 32'sd1235717, 32'sd1389911, 32'sd33133, 32'sd600913, 32'sd2738824, 32'sd1696700, 32'sd145126, 32'sd861475, 32'sd1561639, 32'sd261072, 32'sd872401, 32'sd739070, -32'sd230946, 32'sd242154, 32'sd266321, 32'sd1302339, -32'sd2208838, -32'sd1940886, -32'sd4096103, -32'sd2194247, -32'sd1000944, -32'sd70997, -32'sd1788452, -32'sd1946444, 32'sd1449801, 32'sd3291398, 32'sd31565, 32'sd1162, -32'sd364592, 32'sd1333608, -32'sd1544054, 32'sd69571, 32'sd720479, 32'sd737499, 32'sd1851525, -32'sd54335, 32'sd89268, 32'sd1666831, -32'sd809887, -32'sd272530, 32'sd305391, -32'sd202689, 32'sd997646, 32'sd541374, 32'sd713223, -32'sd2278008, -32'sd2903034, -32'sd1022337, -32'sd925922, -32'sd651579, -32'sd1067992, -32'sd651814, 32'sd2152160, 32'sd418864, 32'sd1866990, 32'sd1742440, 32'sd246035, -32'sd676019, -32'sd2226242, -32'sd1597984, -32'sd1504608, 32'sd142976, 32'sd2078168, 32'sd1866658, 32'sd708390, 32'sd975956, -32'sd4130, -32'sd1056893, -32'sd36070, -32'sd1644683, 32'sd1116408, -32'sd209134, -32'sd30734, -32'sd569827, -32'sd934631, 32'sd525005, -32'sd265435, -32'sd3046371, -32'sd423940, 32'sd1890484, 32'sd250031, 32'sd1884632, -32'sd501552, -32'sd60677, 32'sd1199950, -32'sd2357611, -32'sd2079888, -32'sd2113339, -32'sd2158248, -32'sd1625242, -32'sd1074353, 32'sd546757, 32'sd1697168, 32'sd858872, 32'sd1304473, -32'sd39449, 32'sd585424, 32'sd247037, 32'sd733112, 32'sd112042, -32'sd492935, -32'sd1615431, -32'sd478013, 32'sd66958, 32'sd1349843, -32'sd251737, -32'sd1983259, -32'sd521995, 32'sd1636970, 32'sd1709419, 32'sd2309163, 32'sd311457, -32'sd305055, -32'sd1838509, -32'sd1528812, -32'sd2756448, -32'sd3205902, -32'sd2312706, -32'sd834746, -32'sd836327, 32'sd795932, -32'sd1474639, 32'sd1129579, 32'sd627851, -32'sd90438, -32'sd140401, -32'sd368797, 32'sd2150615, -32'sd1198025, -32'sd2008801, 32'sd238133, 32'sd200769, 32'sd22603, 32'sd6397, -32'sd1166210, 32'sd732473, 32'sd2388899, 32'sd2641814, 32'sd4313875, -32'sd831627, -32'sd360282, 32'sd151151, -32'sd3329256, -32'sd1813288, -32'sd2122843, -32'sd255474, -32'sd1015581, -32'sd385335, -32'sd1840924, -32'sd847951, 32'sd1210910, -32'sd1266226, 32'sd2503176, 32'sd925361, 32'sd379023, 32'sd747009, -32'sd1268189, 32'sd144677, 32'sd872083, -32'sd120313, -32'sd868889, -32'sd660530, 32'sd413458, -32'sd512846, 32'sd433096, 32'sd354031, 32'sd639201, -32'sd2111451, -32'sd68170, -32'sd2968161, -32'sd1887854, -32'sd267036, 32'sd247308, -32'sd602045, -32'sd2675257, -32'sd190935, 32'sd1053082, -32'sd1134522, 32'sd376473, 32'sd1053151, 32'sd1827319, 32'sd1535572, -32'sd1888571, 32'sd764763, -32'sd514631, 32'sd2649320, 32'sd622824, -32'sd405771, -32'sd1561902, 32'sd88070, 32'sd712621, -32'sd682991, 32'sd1190617, 32'sd591043, -32'sd329459, -32'sd3115117, -32'sd1636708, -32'sd858407, 32'sd38198, -32'sd578790, 32'sd461494, -32'sd2128787, -32'sd2457363, 32'sd261006, -32'sd859246, -32'sd1058811, -32'sd1055366, 32'sd798850, 32'sd1093411, 32'sd386174, 32'sd29685, -32'sd149295, 32'sd1594709, 32'sd549141, -32'sd1272064, -32'sd790480, -32'sd1598814, -32'sd2414509, 32'sd549625, 32'sd571885, 32'sd711154, -32'sd1321598, 32'sd32579, -32'sd1148569, -32'sd551303, -32'sd1862749, -32'sd1015026, 32'sd348646, -32'sd1391448, -32'sd1300945, -32'sd440329, -32'sd754926, -32'sd1165635, -32'sd1951478, -32'sd605431, -32'sd835833, 32'sd0, 32'sd473624, -32'sd710095, 32'sd266456, 32'sd1432476, 32'sd1951233, 32'sd1395852, 32'sd1206687, -32'sd956974, -32'sd1552064, -32'sd1294601, -32'sd545355, -32'sd3374093, -32'sd1992585, 32'sd949789, 32'sd1070752, -32'sd588808, 32'sd1242814, -32'sd381231, 32'sd246590, -32'sd449865, -32'sd1225562, 32'sd1211942, -32'sd1224104, -32'sd540257, -32'sd689059, -32'sd2323146, 32'sd458896, 32'sd32494, 32'sd1284364, -32'sd364606, 32'sd1993450, 32'sd1589770, -32'sd45097, 32'sd1082152, 32'sd2508891, -32'sd589940, 32'sd140819, -32'sd48658, -32'sd1628171, -32'sd2776773, 32'sd696499, 32'sd2055979, 32'sd2696110, 32'sd1477707, 32'sd1589775, 32'sd311071, -32'sd842281, -32'sd526780, 32'sd493078, -32'sd1300382, -32'sd860681, -32'sd1456194, -32'sd70278, -32'sd1450951, 32'sd675882, 32'sd864078, 32'sd293351, -32'sd899682, -32'sd1251130, -32'sd1014499, 32'sd2379787, 32'sd1628857, 32'sd1355862, 32'sd513213, 32'sd785265, 32'sd2158866, 32'sd1809097, 32'sd1516993, 32'sd1706491, 32'sd2960042, 32'sd2657752, 32'sd1788243, -32'sd655410, -32'sd1245027, -32'sd691195, -32'sd761408, -32'sd363403, 32'sd751644, 32'sd168579, 32'sd355682, 32'sd101739, -32'sd1488182, 32'sd430229, 32'sd0, 32'sd96847, 32'sd1574751, -32'sd1402018, 32'sd152788, 32'sd868702, 32'sd890216, -32'sd733103, 32'sd1140014, 32'sd579467, 32'sd2748401, 32'sd2304725, 32'sd561254, 32'sd2253703, 32'sd3088566, 32'sd974008, 32'sd1573083, 32'sd502055, -32'sd2381243, -32'sd26995, -32'sd877140, -32'sd1791657, -32'sd134887, 32'sd58200, 32'sd1436129, 32'sd28564, -32'sd745285, 32'sd881336, 32'sd493734, -32'sd269846, -32'sd504856, 32'sd1564287, -32'sd522732, -32'sd148024, 32'sd77488, -32'sd148307, -32'sd473708, 32'sd689561, 32'sd2556396, 32'sd2131079, 32'sd1947073, 32'sd2046877, -32'sd823899, 32'sd233844, 32'sd536943, 32'sd84028, -32'sd1853855, -32'sd768527, -32'sd1687928, -32'sd942087, 32'sd201203, 32'sd624387, 32'sd1238544, -32'sd538500, -32'sd1117047, 32'sd586421, 32'sd84567, 32'sd387090, 32'sd1246817, 32'sd657440, -32'sd658343, -32'sd1826278, 32'sd41598, 32'sd573391, -32'sd1496507, 32'sd1046155, 32'sd296317, 32'sd1413582, 32'sd1812899, 32'sd64689, -32'sd1323385, -32'sd524561, -32'sd1906730, -32'sd1100566, -32'sd2245519, -32'sd1134808, -32'sd949403, -32'sd2017027, -32'sd37896, -32'sd281405, 32'sd2410299, 32'sd529489, 32'sd599436, 32'sd805990, 32'sd0, 32'sd1253564, -32'sd196604, -32'sd1062681, -32'sd1576863, 32'sd798248, -32'sd574870, -32'sd314196, 32'sd197491, -32'sd824149, 32'sd336431, -32'sd1736746, -32'sd1146970, -32'sd1689836, -32'sd348741, -32'sd1217578, -32'sd2251725, -32'sd1107892, -32'sd461497, -32'sd1009928, -32'sd847323, -32'sd1068909, -32'sd152031, 32'sd1811132, -32'sd220341, 32'sd828005, 32'sd1008960, 32'sd0, 32'sd0, 32'sd0, 32'sd877251, -32'sd1347681, 32'sd393020, -32'sd1091087, -32'sd394445, -32'sd1302350, 32'sd231009, -32'sd1141145, -32'sd2390949, -32'sd2579955, -32'sd1207528, -32'sd3043385, -32'sd3402978, -32'sd1793879, -32'sd1697983, -32'sd2051048, -32'sd1675343, 32'sd175600, 32'sd636376, -32'sd1123936, -32'sd830823, 32'sd1313465, -32'sd547004, 32'sd124506, -32'sd317455, 32'sd0, 32'sd0, 32'sd0, 32'sd519887, -32'sd905470, 32'sd473925, 32'sd764040, 32'sd785263, 32'sd510939, -32'sd941381, -32'sd1936048, -32'sd1536789, -32'sd1841105, -32'sd605054, 32'sd103642, -32'sd587274, 32'sd1824050, 32'sd1841957, 32'sd1104433, 32'sd148931, 32'sd542827, 32'sd913182, 32'sd964095, 32'sd968994, 32'sd2034730, 32'sd792771, -32'sd1149543, 32'sd837350, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1069738, -32'sd1320439, -32'sd464630, -32'sd1193080, 32'sd365491, -32'sd1402854, 32'sd25732, 32'sd1563993, 32'sd2253870, 32'sd1260815, -32'sd121735, 32'sd212546, 32'sd1048266, -32'sd735713, 32'sd253162, 32'sd1278587, 32'sd388463, -32'sd884428, 32'sd894959, -32'sd492180, -32'sd58631, 32'sd1564746, 32'sd578057, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2205531, 32'sd1612161, 32'sd620628, 32'sd2032401, -32'sd767282, -32'sd112203, 32'sd214055, 32'sd1048967, 32'sd388607, -32'sd469942, 32'sd1497816, 32'sd572672, -32'sd399231, -32'sd500948, 32'sd1063847, -32'sd122121, -32'sd216671, 32'sd259179, -32'sd134517, 32'sd2018676, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd612057, -32'sd278060, 32'sd572348, 32'sd482442, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd444935, 32'sd889091, -32'sd299793, 32'sd1924802, 32'sd1635271, -32'sd316319, 32'sd698897, -32'sd87911, 32'sd32904, 32'sd1226008, 32'sd475702, 32'sd911733, 32'sd506058, 32'sd661173, 32'sd217544, 32'sd1128699, 32'sd606434, 32'sd1698920, -32'sd560846, 32'sd341766, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd436654, 32'sd763755, 32'sd628774, 32'sd1266370, -32'sd378850, -32'sd121140, -32'sd1257020, -32'sd850514, 32'sd497320, -32'sd456578, -32'sd244513, 32'sd464302, 32'sd450906, 32'sd2623274, 32'sd368623, 32'sd415877, 32'sd444869, 32'sd894761, 32'sd918008, 32'sd563444, 32'sd1156852, -32'sd108750, -32'sd136789, 32'sd395394, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd962174, -32'sd583498, 32'sd517152, -32'sd822385, -32'sd479616, 32'sd1267801, -32'sd50685, -32'sd710097, 32'sd863234, -32'sd862429, -32'sd819298, -32'sd452919, 32'sd159271, 32'sd3433934, 32'sd2244474, -32'sd1914706, 32'sd456465, -32'sd1545588, -32'sd77401, -32'sd68753, -32'sd738191, -32'sd40384, 32'sd1259063, -32'sd1076203, 32'sd303737, 32'sd0, 32'sd0, 32'sd1016427, 32'sd5351, 32'sd1357158, 32'sd329034, 32'sd223787, 32'sd1298470, 32'sd612096, 32'sd130236, 32'sd2254901, 32'sd2174896, 32'sd576023, 32'sd1304597, 32'sd425305, -32'sd649516, 32'sd1364110, 32'sd1291351, 32'sd825995, 32'sd1767757, 32'sd1343593, -32'sd249504, -32'sd737882, -32'sd2291088, -32'sd1569028, -32'sd985098, -32'sd589254, -32'sd205663, 32'sd1039440, 32'sd0, 32'sd354159, -32'sd305560, -32'sd70713, 32'sd146406, 32'sd639448, -32'sd267221, -32'sd184384, 32'sd943397, 32'sd836905, 32'sd1010696, -32'sd338589, 32'sd167454, 32'sd1277220, 32'sd1052171, 32'sd8299, 32'sd785615, -32'sd146990, -32'sd98555, -32'sd781800, 32'sd323202, 32'sd787315, -32'sd1564948, -32'sd260164, 32'sd1010648, 32'sd611316, -32'sd1307522, 32'sd152130, 32'sd0, 32'sd1191199, -32'sd768552, 32'sd153466, 32'sd607530, 32'sd115050, -32'sd477261, -32'sd330603, 32'sd1281603, 32'sd357475, -32'sd1069337, -32'sd867231, -32'sd555663, -32'sd585832, 32'sd1007711, 32'sd541761, 32'sd2619817, 32'sd2504720, -32'sd1222243, 32'sd667829, -32'sd1024316, -32'sd1214594, 32'sd956525, 32'sd1429707, 32'sd316783, -32'sd361116, 32'sd582613, -32'sd593142, 32'sd594092, 32'sd48110, 32'sd821428, 32'sd677018, 32'sd87320, 32'sd747228, 32'sd1274977, 32'sd263971, 32'sd481709, 32'sd1221018, 32'sd61378, -32'sd749019, 32'sd624246, -32'sd1318717, 32'sd235482, 32'sd988414, 32'sd2083324, 32'sd2501850, 32'sd194660, 32'sd941874, 32'sd51171, 32'sd1164902, -32'sd775102, 32'sd903121, 32'sd967826, 32'sd874527, 32'sd1365488, -32'sd186767, 32'sd637378, -32'sd38988, 32'sd1449232, 32'sd2245907, -32'sd320936, 32'sd1554527, -32'sd855598, 32'sd60233, 32'sd1956573, 32'sd1846598, 32'sd1710702, -32'sd597750, -32'sd1874478, -32'sd378668, -32'sd306636, 32'sd1884142, -32'sd1290362, 32'sd429026, 32'sd275222, -32'sd739256, -32'sd1301823, -32'sd74698, 32'sd1348434, 32'sd2300311, 32'sd2212174, 32'sd177485, 32'sd1515188, -32'sd50807, 32'sd1470004, 32'sd367387, -32'sd98847, -32'sd1228109, 32'sd453951, 32'sd577455, 32'sd873845, -32'sd7237, 32'sd3312287, 32'sd1186600, 32'sd2030371, -32'sd574348, 32'sd498918, -32'sd237539, -32'sd1594426, -32'sd1978423, -32'sd3035744, -32'sd158188, -32'sd2370622, -32'sd1336472, -32'sd726295, -32'sd717233, 32'sd975091, 32'sd240833, 32'sd1195164, 32'sd880488, -32'sd203072, -32'sd1145025, 32'sd1595910, 32'sd1007599, -32'sd1172644, 32'sd1212475, 32'sd1020623, -32'sd47929, -32'sd489612, 32'sd384661, 32'sd1833347, 32'sd2620703, -32'sd301020, 32'sd142159, -32'sd340520, -32'sd1690185, -32'sd695574, -32'sd1707396, -32'sd1752204, -32'sd1852338, -32'sd277919, -32'sd859946, 32'sd605989, -32'sd736573, -32'sd1402099, -32'sd1349491, -32'sd1191121, -32'sd595757, 32'sd623385, 32'sd684600, 32'sd99971, 32'sd505721, -32'sd256937, -32'sd296132, 32'sd1362233, 32'sd495273, -32'sd53830, 32'sd235721, 32'sd803957, 32'sd1057010, 32'sd2700619, 32'sd1623434, 32'sd2284339, 32'sd2467718, 32'sd1863525, 32'sd2199735, -32'sd331158, -32'sd559546, 32'sd946705, 32'sd534501, -32'sd825556, -32'sd1897914, -32'sd2713088, -32'sd3202091, -32'sd755230, -32'sd1801190, -32'sd390090, -32'sd348372, 32'sd241984, 32'sd953127, -32'sd620862, -32'sd1546880, -32'sd943602, 32'sd839258, 32'sd68024, -32'sd571461, 32'sd1445383, 32'sd273332, 32'sd3250770, 32'sd3754292, 32'sd3323506, 32'sd4310584, 32'sd4146207, 32'sd2416938, 32'sd1134048, 32'sd2084673, 32'sd2689561, 32'sd981342, -32'sd398628, -32'sd1284712, -32'sd959406, -32'sd1295126, -32'sd3943101, -32'sd2121460, -32'sd1059704, -32'sd228823, 32'sd99822, -32'sd1046563, -32'sd2357655, -32'sd130457, -32'sd638168, -32'sd994946, -32'sd1247364, 32'sd193056, 32'sd992546, 32'sd533554, 32'sd1310549, 32'sd3200602, 32'sd3954594, 32'sd5023375, 32'sd5485772, 32'sd2850625, 32'sd1731793, 32'sd1479934, 32'sd2855067, -32'sd479740, 32'sd430184, -32'sd50899, 32'sd1102700, 32'sd133925, -32'sd1564731, -32'sd85989, -32'sd739504, 32'sd630374, 32'sd2108959, 32'sd528491, 32'sd297378, -32'sd1500915, -32'sd2413227, -32'sd2548567, -32'sd3704090, -32'sd462034, -32'sd144658, -32'sd1912952, 32'sd1080002, 32'sd476310, 32'sd2362703, 32'sd2095853, 32'sd2481669, 32'sd1598189, 32'sd1130217, 32'sd1043868, -32'sd150435, -32'sd1564774, -32'sd1302273, -32'sd221000, 32'sd1050190, 32'sd606306, 32'sd1402164, 32'sd27584, -32'sd587920, 32'sd162069, 32'sd1615296, 32'sd287888, 32'sd661977, -32'sd387923, -32'sd2279867, -32'sd3701001, -32'sd4166863, -32'sd4025920, -32'sd1898183, -32'sd3492314, -32'sd2916885, -32'sd273192, 32'sd721719, 32'sd985401, 32'sd401006, 32'sd955598, 32'sd762661, 32'sd395872, 32'sd623110, 32'sd47397, -32'sd314262, -32'sd150002, 32'sd329409, 32'sd2066043, 32'sd1891017, 32'sd525620, -32'sd479213, 32'sd955773, 32'sd106801, -32'sd586518, -32'sd663478, 32'sd2069506, -32'sd473284, -32'sd2039484, -32'sd2544981, -32'sd3447489, -32'sd4215545, -32'sd5842694, -32'sd5885842, -32'sd5074966, -32'sd2837394, -32'sd1825038, -32'sd1070498, -32'sd489229, -32'sd768877, 32'sd1622069, 32'sd612959, 32'sd885082, 32'sd804151, -32'sd174083, 32'sd65667, 32'sd831195, 32'sd1162117, -32'sd459701, 32'sd248528, 32'sd618747, 32'sd0, 32'sd1110439, -32'sd1073152, 32'sd768286, -32'sd1073857, -32'sd1047736, 32'sd558032, -32'sd7619, -32'sd1504319, -32'sd4184257, -32'sd5969924, -32'sd5737278, -32'sd7364009, -32'sd5047031, -32'sd2901056, -32'sd2470074, -32'sd1365952, -32'sd806308, -32'sd1406512, 32'sd944210, -32'sd439763, -32'sd268995, -32'sd1009900, 32'sd1714413, 32'sd353775, 32'sd649298, 32'sd538908, -32'sd205305, 32'sd97619, -32'sd601097, 32'sd1157658, 32'sd2477302, 32'sd1588956, 32'sd807608, 32'sd1435266, 32'sd740232, -32'sd997933, -32'sd1654971, -32'sd2937811, -32'sd3217120, -32'sd4894309, -32'sd4672751, -32'sd3019329, -32'sd3056948, 32'sd1086342, 32'sd397378, -32'sd589453, 32'sd1429035, 32'sd85254, 32'sd1627598, -32'sd1321513, -32'sd109827, 32'sd768330, -32'sd759576, -32'sd574556, 32'sd446656, 32'sd842848, 32'sd398059, 32'sd783319, 32'sd495418, 32'sd1677817, 32'sd2355707, 32'sd2035386, 32'sd1450516, 32'sd1296679, 32'sd512093, 32'sd2457320, 32'sd363943, -32'sd1819577, -32'sd3326346, -32'sd1587688, -32'sd1843400, -32'sd900750, -32'sd1015347, -32'sd1653556, 32'sd1393428, -32'sd1438655, 32'sd454937, 32'sd96681, 32'sd481596, 32'sd1470581, -32'sd621367, -32'sd1982051, -32'sd2600786, 32'sd0, -32'sd442704, -32'sd113856, 32'sd1427729, 32'sd1098506, 32'sd1023830, 32'sd300338, -32'sd61816, 32'sd409952, 32'sd1245535, 32'sd3068290, 32'sd1990480, 32'sd527901, -32'sd1554835, -32'sd765552, 32'sd35933, -32'sd590190, -32'sd18865, -32'sd826541, 32'sd908889, -32'sd1618516, 32'sd309662, 32'sd903189, 32'sd151800, 32'sd662083, -32'sd1175231, -32'sd540433, 32'sd783170, 32'sd1236728, 32'sd576164, 32'sd469139, -32'sd1376970, 32'sd821759, 32'sd2747000, 32'sd1255730, 32'sd976529, 32'sd449543, 32'sd485605, 32'sd872394, 32'sd1884077, 32'sd1404934, 32'sd1979577, 32'sd1918189, 32'sd1205655, -32'sd541686, 32'sd63609, -32'sd1245772, 32'sd297999, 32'sd1206687, 32'sd996932, -32'sd1737323, -32'sd1499215, 32'sd368078, -32'sd3082375, -32'sd773318, 32'sd322941, 32'sd1945416, 32'sd1945301, 32'sd478424, 32'sd1114459, 32'sd8382, -32'sd1143316, 32'sd1135103, -32'sd536644, 32'sd1310222, -32'sd1387725, 32'sd1903637, 32'sd1223147, -32'sd1472949, -32'sd698643, 32'sd1814914, -32'sd878687, 32'sd1109835, 32'sd1580336, 32'sd111188, -32'sd460339, -32'sd100606, 32'sd47169, -32'sd3842757, -32'sd1126611, -32'sd315354, -32'sd566307, 32'sd880838, 32'sd94477, 32'sd0, 32'sd1002382, -32'sd1387080, -32'sd180750, 32'sd201513, -32'sd1893994, -32'sd279914, -32'sd1046498, -32'sd447898, -32'sd1410106, 32'sd1938379, -32'sd619499, -32'sd818762, 32'sd394852, -32'sd661899, 32'sd1036325, 32'sd1546300, -32'sd226741, -32'sd485874, -32'sd277471, -32'sd998919, -32'sd724046, -32'sd977921, 32'sd183402, 32'sd1463475, -32'sd1737243, -32'sd332938, 32'sd0, 32'sd0, 32'sd0, 32'sd423854, -32'sd888196, 32'sd1657750, -32'sd1431550, -32'sd1072844, 32'sd1139054, -32'sd770075, 32'sd150921, 32'sd582593, -32'sd104172, 32'sd635241, -32'sd599095, -32'sd3273063, -32'sd2325480, -32'sd1311077, -32'sd1404432, -32'sd1838382, -32'sd91708, -32'sd371737, -32'sd152024, -32'sd1087184, -32'sd983040, -32'sd500414, 32'sd510454, 32'sd747962, 32'sd0, 32'sd0, 32'sd0, 32'sd1513184, 32'sd169465, 32'sd410545, 32'sd411173, 32'sd416991, 32'sd1164347, -32'sd691360, -32'sd1179976, 32'sd1414051, 32'sd173422, -32'sd104974, 32'sd420049, -32'sd839888, 32'sd59484, -32'sd11260, -32'sd898905, -32'sd1881955, -32'sd2395080, 32'sd152919, 32'sd79614, -32'sd797816, -32'sd1416198, -32'sd773423, 32'sd566972, 32'sd931104, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd346735, -32'sd116177, 32'sd25658, -32'sd4514, -32'sd132054, 32'sd523357, 32'sd582445, 32'sd843995, 32'sd589401, 32'sd360500, 32'sd1173256, 32'sd1094408, 32'sd1297174, -32'sd1180588, 32'sd502080, 32'sd191287, -32'sd469575, -32'sd1221992, -32'sd79306, -32'sd998402, -32'sd163968, 32'sd739183, 32'sd543348, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1200580, 32'sd1153105, -32'sd547921, 32'sd748082, -32'sd214441, 32'sd677206, -32'sd1248301, -32'sd1000630, -32'sd1360092, -32'sd312666, 32'sd722165, 32'sd141346, 32'sd212702, -32'sd312841, 32'sd575347, 32'sd994500, -32'sd545766, -32'sd1874384, -32'sd1041244, 32'sd628680, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd466339, 32'sd262774, 32'sd1613909, 32'sd1413168, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd74766, -32'sd777880, -32'sd166650, -32'sd418837, -32'sd1440947, 32'sd1376008, 32'sd1641833, -32'sd389569, 32'sd401260, -32'sd520438, 32'sd810683, -32'sd765018, 32'sd1559021, 32'sd295746, 32'sd969016, -32'sd529948, 32'sd69840, 32'sd1400241, 32'sd1073969, 32'sd1073817, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd755605, -32'sd797124, 32'sd357898, 32'sd1052940, -32'sd136340, -32'sd629830, -32'sd118736, 32'sd53970, 32'sd486393, 32'sd815033, 32'sd1307571, 32'sd439634, 32'sd29896, -32'sd544708, -32'sd609646, 32'sd524572, -32'sd928156, -32'sd1153195, 32'sd625190, -32'sd531570, 32'sd555974, 32'sd632059, 32'sd285790, 32'sd97384, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd117315, -32'sd488377, 32'sd1632788, -32'sd221824, 32'sd206760, -32'sd1064725, 32'sd607614, 32'sd68477, 32'sd721944, 32'sd1138057, -32'sd347497, 32'sd1930848, -32'sd942661, -32'sd1041308, 32'sd1512703, 32'sd385354, -32'sd430720, -32'sd75802, -32'sd71570, -32'sd421158, -32'sd2309991, -32'sd287486, 32'sd595118, 32'sd741269, 32'sd1226235, 32'sd0, 32'sd0, 32'sd729831, 32'sd602383, -32'sd2046956, -32'sd111153, 32'sd67184, 32'sd1465381, 32'sd2057251, 32'sd455092, 32'sd952104, -32'sd2336826, 32'sd503908, 32'sd738989, 32'sd2174862, 32'sd2105500, 32'sd1328378, 32'sd218487, -32'sd156014, 32'sd1010972, 32'sd1392529, -32'sd330588, -32'sd548410, -32'sd638480, -32'sd302876, 32'sd593271, -32'sd1668835, 32'sd648449, 32'sd427507, 32'sd0, 32'sd934290, -32'sd561575, 32'sd1396138, 32'sd1201457, 32'sd73622, 32'sd1676618, -32'sd232560, 32'sd619291, -32'sd597024, -32'sd771762, -32'sd203913, 32'sd2055555, 32'sd1961525, 32'sd1699306, 32'sd1409339, 32'sd1880738, -32'sd1602715, -32'sd1145925, -32'sd1850418, -32'sd691164, -32'sd610406, 32'sd60644, -32'sd1853984, -32'sd1007144, -32'sd6662, 32'sd56589, 32'sd582789, 32'sd0, 32'sd123271, -32'sd382956, 32'sd1352111, -32'sd836923, -32'sd1415211, 32'sd390550, -32'sd1425760, -32'sd467773, 32'sd667040, 32'sd2086157, 32'sd295115, 32'sd1289358, 32'sd1981025, 32'sd283221, 32'sd2588831, 32'sd2065953, 32'sd145551, -32'sd224351, -32'sd680421, -32'sd481108, 32'sd1795659, 32'sd379228, -32'sd1059238, 32'sd526757, 32'sd56101, -32'sd244476, -32'sd627207, 32'sd1304328, 32'sd231143, 32'sd79706, 32'sd1802826, 32'sd1897460, 32'sd566580, 32'sd160616, 32'sd586277, -32'sd669885, 32'sd1110390, 32'sd1240683, 32'sd2349304, 32'sd1253660, 32'sd2160324, 32'sd1705403, 32'sd997860, 32'sd3066278, 32'sd829825, -32'sd322838, -32'sd38544, -32'sd393188, -32'sd977957, -32'sd1059836, -32'sd870965, -32'sd23710, 32'sd1046807, 32'sd1020168, -32'sd32277, 32'sd1039135, -32'sd864863, 32'sd1266660, 32'sd888036, -32'sd1410942, -32'sd201695, -32'sd557843, 32'sd638016, -32'sd1410846, -32'sd368211, 32'sd723629, 32'sd1527033, 32'sd406828, 32'sd1068081, 32'sd2767566, 32'sd802374, 32'sd2467643, 32'sd3269699, -32'sd715687, 32'sd658234, -32'sd289495, 32'sd338286, -32'sd710115, 32'sd730241, 32'sd321123, -32'sd3880, 32'sd1600511, 32'sd901918, 32'sd812275, -32'sd1997691, 32'sd1239029, -32'sd104663, 32'sd66991, 32'sd1392532, -32'sd955666, 32'sd81685, -32'sd937016, 32'sd103998, 32'sd602036, -32'sd2516584, -32'sd636907, -32'sd1356001, -32'sd569105, 32'sd1099284, 32'sd1500821, 32'sd1975905, 32'sd2708367, 32'sd1094914, -32'sd802642, -32'sd1716815, -32'sd550288, 32'sd1192138, -32'sd1227938, 32'sd743324, -32'sd929896, 32'sd1065467, -32'sd912229, 32'sd172212, 32'sd1461995, 32'sd2549950, 32'sd788428, 32'sd1878693, 32'sd629366, 32'sd947039, -32'sd73771, -32'sd1373954, -32'sd948971, -32'sd1516766, -32'sd1631406, -32'sd2257896, -32'sd3560963, -32'sd3126413, 32'sd1607147, 32'sd3248594, 32'sd1689969, -32'sd937526, -32'sd1602435, 32'sd689648, -32'sd1249082, 32'sd554234, 32'sd50075, 32'sd485931, -32'sd1198208, -32'sd1648739, -32'sd1287731, -32'sd285775, -32'sd448009, 32'sd489156, 32'sd796561, -32'sd311786, -32'sd859157, 32'sd1166258, -32'sd402672, -32'sd568536, -32'sd1205993, -32'sd1896414, -32'sd1211474, -32'sd2650791, -32'sd5086507, -32'sd963089, -32'sd410475, 32'sd2217587, 32'sd1641553, -32'sd471720, -32'sd551815, -32'sd406312, -32'sd1584814, -32'sd376323, -32'sd1730026, -32'sd1260513, -32'sd675456, -32'sd51509, 32'sd1065639, 32'sd585145, 32'sd379821, -32'sd1371310, -32'sd1479478, -32'sd1236445, 32'sd49337, 32'sd508547, 32'sd317718, -32'sd332550, -32'sd821471, -32'sd1660751, -32'sd1093804, -32'sd4223696, -32'sd4957650, -32'sd2962140, -32'sd1334380, 32'sd1803583, 32'sd1201954, -32'sd1521911, -32'sd909219, -32'sd938734, -32'sd2186859, 32'sd544975, -32'sd1292033, -32'sd253717, -32'sd1112960, -32'sd347487, 32'sd488854, 32'sd908870, -32'sd1705298, 32'sd205764, -32'sd2494959, -32'sd893443, -32'sd734048, -32'sd1610880, -32'sd970527, 32'sd240819, 32'sd370769, -32'sd375687, -32'sd1753188, -32'sd2210072, -32'sd4139207, -32'sd3076323, 32'sd540395, 32'sd1745377, -32'sd393320, -32'sd629103, -32'sd163638, -32'sd1250806, -32'sd2608374, -32'sd430093, 32'sd503319, -32'sd896914, 32'sd459634, 32'sd1793578, 32'sd1088511, -32'sd893213, 32'sd386077, -32'sd929778, -32'sd579701, -32'sd569956, -32'sd843750, -32'sd261208, -32'sd1574744, -32'sd939411, -32'sd484008, -32'sd2645454, -32'sd1307283, -32'sd3014677, -32'sd1417359, -32'sd1392690, 32'sd445781, 32'sd1076884, 32'sd1332304, -32'sd2240173, -32'sd793198, -32'sd1908503, -32'sd814687, -32'sd1601854, 32'sd76500, -32'sd204814, 32'sd902007, 32'sd2565689, 32'sd515674, 32'sd738320, -32'sd394712, 32'sd1016391, -32'sd1738500, 32'sd18317, -32'sd1417579, -32'sd905408, -32'sd1137939, 32'sd484414, -32'sd820090, -32'sd1144244, -32'sd1212179, -32'sd2099197, -32'sd2061594, -32'sd1038351, -32'sd1960422, -32'sd593207, -32'sd1928222, -32'sd1936290, -32'sd1298049, -32'sd173009, -32'sd1463845, -32'sd1325573, -32'sd596406, 32'sd345696, 32'sd1172191, -32'sd37460, 32'sd903138, 32'sd906977, 32'sd586166, -32'sd2188886, -32'sd876371, -32'sd851072, 32'sd572730, -32'sd2112509, -32'sd1142630, -32'sd385630, 32'sd312434, 32'sd730588, 32'sd2224215, -32'sd1679021, -32'sd3444562, -32'sd2339123, -32'sd652651, -32'sd1299866, -32'sd727196, -32'sd442736, 32'sd198702, 32'sd434393, 32'sd78122, -32'sd1152361, 32'sd254015, -32'sd1449989, -32'sd1605564, 32'sd221675, 32'sd0, -32'sd710398, 32'sd136918, -32'sd1089346, 32'sd336998, -32'sd1868825, -32'sd1297154, -32'sd423939, -32'sd940401, -32'sd318769, 32'sd2301694, 32'sd773707, -32'sd608999, -32'sd2739293, -32'sd1568025, -32'sd2422955, -32'sd1326457, -32'sd679264, -32'sd792693, 32'sd641099, -32'sd1437174, -32'sd2011456, -32'sd1601823, -32'sd1411651, -32'sd1448486, 32'sd1479240, -32'sd128949, 32'sd572944, 32'sd29957, 32'sd21343, -32'sd829004, -32'sd2129623, -32'sd870719, -32'sd902074, 32'sd42242, 32'sd57869, -32'sd342394, 32'sd184826, 32'sd1895062, 32'sd995326, 32'sd2142601, 32'sd104073, -32'sd2482014, -32'sd2029911, -32'sd1578551, -32'sd411977, -32'sd1966899, 32'sd35256, -32'sd66394, -32'sd2028323, -32'sd1574161, -32'sd1265712, -32'sd22514, -32'sd107059, 32'sd997111, -32'sd147734, 32'sd288424, -32'sd125798, 32'sd1237285, -32'sd975432, -32'sd165865, -32'sd1959074, 32'sd872469, 32'sd2582453, 32'sd281250, -32'sd184411, 32'sd326242, 32'sd1260794, -32'sd599195, 32'sd250539, -32'sd2826965, -32'sd128964, -32'sd89333, -32'sd415777, -32'sd1544595, -32'sd466953, 32'sd2723352, -32'sd222008, 32'sd4650, -32'sd1566137, -32'sd1064161, 32'sd1714759, 32'sd1536552, 32'sd939147, 32'sd0, -32'sd436424, -32'sd790324, 32'sd1216467, -32'sd1137369, 32'sd848164, 32'sd1462773, 32'sd688627, 32'sd2456198, -32'sd1071250, 32'sd2358368, 32'sd3153651, 32'sd2826071, 32'sd1983335, 32'sd2086614, 32'sd2127307, 32'sd938259, -32'sd750230, -32'sd158271, -32'sd361401, 32'sd2161503, 32'sd1078101, -32'sd1192972, 32'sd430766, -32'sd644370, -32'sd662517, -32'sd902958, -32'sd418448, 32'sd132918, -32'sd1509381, -32'sd834560, -32'sd433687, -32'sd1174328, 32'sd1339357, 32'sd63702, -32'sd761544, 32'sd1161858, 32'sd951629, 32'sd867045, 32'sd2650973, 32'sd2267838, 32'sd1599835, 32'sd2700419, 32'sd3403889, 32'sd1227213, 32'sd465232, 32'sd974252, 32'sd461085, 32'sd361012, -32'sd68908, -32'sd1056897, 32'sd1257320, -32'sd1893543, -32'sd436448, 32'sd484788, 32'sd522923, 32'sd319384, -32'sd243521, 32'sd641627, 32'sd334404, -32'sd761264, 32'sd1408053, -32'sd249492, 32'sd261021, 32'sd260584, 32'sd948371, -32'sd772929, 32'sd973126, -32'sd336350, 32'sd1466514, 32'sd2470778, 32'sd1313307, 32'sd1121232, 32'sd1379795, 32'sd1466528, -32'sd111743, -32'sd750651, -32'sd417345, 32'sd1376250, 32'sd1347269, 32'sd679436, 32'sd73038, -32'sd1195401, 32'sd691268, 32'sd0, 32'sd370206, -32'sd825346, -32'sd1490920, 32'sd134688, 32'sd103573, -32'sd591588, 32'sd594061, 32'sd1072439, 32'sd1722222, -32'sd700589, 32'sd796149, 32'sd513277, -32'sd447412, 32'sd2082995, 32'sd787823, 32'sd151528, -32'sd298134, -32'sd131608, -32'sd75532, -32'sd646840, -32'sd1862181, 32'sd1523312, 32'sd1640848, 32'sd1174066, 32'sd1711803, -32'sd2538866, 32'sd0, 32'sd0, 32'sd0, 32'sd207055, 32'sd373432, 32'sd716659, -32'sd942379, -32'sd1545588, -32'sd679813, 32'sd416736, -32'sd121131, -32'sd191654, 32'sd391183, -32'sd336010, -32'sd1023146, 32'sd1055681, -32'sd411466, -32'sd1498338, 32'sd260739, 32'sd1154849, 32'sd1475982, -32'sd536458, -32'sd554745, 32'sd207487, -32'sd250978, -32'sd268652, -32'sd181655, 32'sd654326, 32'sd0, 32'sd0, 32'sd0, 32'sd680878, 32'sd744878, 32'sd1926780, -32'sd157318, 32'sd1557045, 32'sd903107, 32'sd1887196, 32'sd815264, 32'sd2389032, 32'sd246794, 32'sd1122102, 32'sd220508, 32'sd532524, -32'sd50685, -32'sd423886, 32'sd575830, 32'sd2146827, 32'sd611761, 32'sd1353459, 32'sd1724319, 32'sd1337975, 32'sd139742, 32'sd335565, 32'sd429851, 32'sd935021, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1034396, 32'sd222585, -32'sd990869, 32'sd998632, -32'sd71356, 32'sd1339491, -32'sd515404, -32'sd1815774, -32'sd1907209, 32'sd529098, -32'sd38380, 32'sd632122, -32'sd352460, 32'sd635210, 32'sd974464, 32'sd805918, -32'sd751919, -32'sd1531860, -32'sd2060740, 32'sd619841, -32'sd1252116, 32'sd34693, 32'sd29314, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd768870, 32'sd623217, 32'sd194713, 32'sd778414, -32'sd493833, 32'sd1173693, 32'sd511664, 32'sd1473459, 32'sd826244, 32'sd1210334, 32'sd1910006, 32'sd385827, 32'sd1409489, -32'sd323499, -32'sd576790, 32'sd876670, 32'sd84612, -32'sd1339273, -32'sd622413, 32'sd737653, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd373671, 32'sd388291, -32'sd171359, -32'sd723735, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1526784, 32'sd1733459, 32'sd368823, -32'sd168146, 32'sd702950, 32'sd1095927, -32'sd1115183, -32'sd119880, -32'sd468581, 32'sd549371, -32'sd1415984, -32'sd874333, 32'sd1360877, -32'sd132167, 32'sd325584, 32'sd1501414, 32'sd430572, 32'sd1445410, 32'sd1068085, 32'sd386223, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1486179, 32'sd1087546, 32'sd1228058, 32'sd1827065, 32'sd7996, 32'sd39988, -32'sd1079058, 32'sd441385, -32'sd36339, -32'sd1313138, 32'sd1088119, 32'sd438550, -32'sd1421631, -32'sd1290287, -32'sd196981, -32'sd1480496, 32'sd1224240, -32'sd236903, 32'sd1780798, 32'sd929650, 32'sd582937, 32'sd965479, -32'sd490778, 32'sd1488349, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd266131, 32'sd262037, 32'sd579453, -32'sd1425059, 32'sd139141, 32'sd370602, 32'sd543185, -32'sd663450, -32'sd2615780, 32'sd479888, 32'sd598172, 32'sd124350, -32'sd882271, -32'sd1667294, -32'sd674271, -32'sd434413, 32'sd1390563, -32'sd228697, -32'sd583281, -32'sd1431255, -32'sd370473, -32'sd1828492, -32'sd3519, -32'sd965615, 32'sd610351, 32'sd0, 32'sd0, 32'sd540320, -32'sd22987, 32'sd1365289, -32'sd81223, 32'sd292777, 32'sd212961, 32'sd1017127, -32'sd2098643, 32'sd45988, -32'sd1467194, -32'sd685283, -32'sd596267, -32'sd1158137, -32'sd1349620, -32'sd1713019, -32'sd1948310, -32'sd1791641, 32'sd807954, -32'sd1219735, -32'sd2277052, -32'sd1768646, -32'sd1236836, -32'sd1912051, -32'sd931341, -32'sd2342610, 32'sd804905, 32'sd1110373, 32'sd0, 32'sd14668, 32'sd488409, -32'sd929798, -32'sd455453, 32'sd897957, -32'sd409461, 32'sd682396, -32'sd405620, 32'sd197099, -32'sd1184155, -32'sd1414851, -32'sd2490589, -32'sd3142866, -32'sd4033505, -32'sd4053436, -32'sd3892860, -32'sd3286518, -32'sd597608, 32'sd1745675, 32'sd2781263, -32'sd1890578, -32'sd1328584, -32'sd1695329, -32'sd1771689, -32'sd175107, 32'sd1755228, 32'sd358890, 32'sd0, 32'sd1153119, -32'sd449150, -32'sd1270374, -32'sd108676, -32'sd1012027, -32'sd3128263, -32'sd790989, -32'sd1905385, -32'sd1308443, 32'sd99945, -32'sd480818, -32'sd3369003, -32'sd4294394, -32'sd3446880, -32'sd2637947, -32'sd4049052, -32'sd602598, 32'sd1389773, 32'sd2894828, 32'sd1964094, 32'sd143397, -32'sd74206, 32'sd572136, 32'sd1014681, 32'sd1024834, 32'sd1281722, -32'sd1829342, 32'sd670816, -32'sd537911, -32'sd563300, 32'sd291228, -32'sd274095, 32'sd109698, -32'sd1746265, -32'sd2369537, -32'sd313689, -32'sd506180, 32'sd486983, -32'sd1530898, -32'sd932759, 32'sd532841, -32'sd96459, 32'sd2336259, 32'sd599293, 32'sd2389189, 32'sd1266429, 32'sd2956565, 32'sd3246604, 32'sd2603581, -32'sd826171, 32'sd1280990, 32'sd136437, -32'sd889300, 32'sd2149318, 32'sd718031, 32'sd148226, 32'sd731396, -32'sd124481, -32'sd1267906, -32'sd2348802, -32'sd2070022, 32'sd238880, -32'sd2304850, -32'sd2426329, -32'sd337413, -32'sd216705, 32'sd910002, 32'sd1597727, 32'sd2497268, 32'sd3711682, 32'sd2893784, 32'sd3864908, 32'sd2135421, 32'sd3084560, 32'sd2932306, 32'sd2841865, 32'sd1955738, 32'sd1685831, -32'sd236073, 32'sd437763, -32'sd56644, -32'sd58902, -32'sd892096, 32'sd121820, -32'sd1068927, -32'sd1071626, 32'sd66135, -32'sd350292, -32'sd1106468, -32'sd1242104, -32'sd603146, -32'sd1250060, -32'sd1423531, 32'sd891291, 32'sd1558579, 32'sd3358195, 32'sd4695833, 32'sd3073445, 32'sd2177268, 32'sd2814408, 32'sd644550, 32'sd3276736, 32'sd4131242, 32'sd9553, 32'sd303808, 32'sd1275860, -32'sd803699, 32'sd2130635, 32'sd669121, -32'sd154524, 32'sd837599, 32'sd1303055, -32'sd568321, -32'sd206088, -32'sd471429, -32'sd552694, 32'sd188661, 32'sd848161, -32'sd971249, -32'sd1175343, 32'sd1006683, 32'sd4052067, 32'sd933317, 32'sd2353783, 32'sd2954696, 32'sd131882, 32'sd2325220, 32'sd994373, -32'sd491212, 32'sd132539, -32'sd195779, -32'sd1301901, -32'sd581380, -32'sd400872, -32'sd2324938, 32'sd948939, 32'sd1560761, 32'sd1270006, 32'sd269826, -32'sd347925, 32'sd100298, -32'sd254548, -32'sd2224397, 32'sd1992850, 32'sd1363420, -32'sd196963, -32'sd1099163, -32'sd1193724, 32'sd2139352, -32'sd926755, 32'sd1938674, 32'sd1339106, 32'sd1630954, 32'sd195335, 32'sd1120517, -32'sd903385, -32'sd1815884, -32'sd990922, -32'sd2239304, -32'sd1800851, -32'sd3200612, -32'sd1224247, -32'sd1657325, -32'sd1483309, 32'sd620887, 32'sd97652, 32'sd2022791, 32'sd233263, 32'sd181955, 32'sd315216, 32'sd489468, 32'sd559178, 32'sd1066647, -32'sd541371, -32'sd1573990, 32'sd618205, 32'sd323301, -32'sd879880, -32'sd767943, -32'sd463754, 32'sd1104951, -32'sd248155, -32'sd595273, -32'sd1381266, -32'sd2722829, 32'sd794118, -32'sd1455943, -32'sd874682, -32'sd619674, -32'sd669690, -32'sd553333, -32'sd187982, -32'sd2360546, -32'sd248508, -32'sd1025310, 32'sd418751, 32'sd215249, 32'sd228808, 32'sd720391, 32'sd92620, -32'sd720305, -32'sd569233, -32'sd996880, -32'sd483147, -32'sd2608290, -32'sd937439, -32'sd420788, -32'sd1095322, 32'sd1034505, -32'sd653278, 32'sd26192, -32'sd2696398, -32'sd2816627, -32'sd1416317, -32'sd11547, -32'sd1154943, -32'sd1918550, -32'sd922058, -32'sd1278579, -32'sd2216488, -32'sd3189251, -32'sd580728, 32'sd300549, 32'sd1124271, 32'sd49003, 32'sd733116, -32'sd766326, 32'sd2430503, -32'sd1262747, 32'sd867397, -32'sd310233, -32'sd1134243, 32'sd210495, -32'sd1501276, -32'sd209481, -32'sd566819, 32'sd652145, 32'sd967859, 32'sd1031473, -32'sd5192, -32'sd2339166, 32'sd151858, -32'sd3110572, 32'sd1084528, -32'sd1343595, -32'sd1362193, -32'sd508523, 32'sd2143966, -32'sd420819, -32'sd1168241, -32'sd3728, 32'sd973654, -32'sd82793, -32'sd1369085, 32'sd3817, 32'sd3391593, 32'sd3248888, 32'sd644884, -32'sd872518, -32'sd720328, -32'sd1209189, 32'sd1544705, -32'sd305792, 32'sd1920447, 32'sd532488, 32'sd748911, -32'sd2035894, -32'sd1471216, -32'sd562021, -32'sd1249532, -32'sd471960, 32'sd325910, 32'sd875685, -32'sd838943, -32'sd1059411, -32'sd183453, 32'sd966793, 32'sd1551895, 32'sd430699, 32'sd134120, 32'sd509713, -32'sd219220, 32'sd5855, 32'sd46452, 32'sd1191755, 32'sd1392718, 32'sd704664, 32'sd981226, -32'sd1259845, -32'sd1331637, 32'sd194534, 32'sd590180, -32'sd505902, -32'sd2015344, -32'sd2264637, -32'sd1359809, -32'sd218133, -32'sd981187, -32'sd657667, -32'sd1271084, -32'sd198094, 32'sd227803, -32'sd1055570, -32'sd320268, 32'sd1502734, 32'sd468205, 32'sd535077, 32'sd0, 32'sd389767, -32'sd745616, 32'sd1761083, -32'sd1946834, 32'sd1674635, 32'sd3225697, 32'sd1744816, 32'sd1199605, 32'sd1359094, 32'sd1170491, -32'sd462312, -32'sd1288889, -32'sd1263479, -32'sd401920, 32'sd202571, -32'sd2382920, -32'sd1963363, 32'sd795299, 32'sd495, -32'sd171128, -32'sd882775, 32'sd393002, 32'sd29780, -32'sd2855930, -32'sd1032846, -32'sd172247, 32'sd115071, 32'sd517497, 32'sd777363, -32'sd656702, 32'sd1115908, -32'sd460112, 32'sd827767, 32'sd1277479, 32'sd3048589, 32'sd1798229, -32'sd119763, -32'sd641625, 32'sd391686, 32'sd661540, -32'sd1410283, 32'sd1746111, -32'sd234864, 32'sd754345, 32'sd204494, -32'sd1662676, 32'sd675610, 32'sd638348, -32'sd1987401, -32'sd1076734, 32'sd859249, -32'sd671505, -32'sd331322, 32'sd1688033, -32'sd1253344, 32'sd369739, -32'sd151603, -32'sd1618895, 32'sd198486, 32'sd830327, -32'sd362683, 32'sd1217568, 32'sd1368307, 32'sd270993, -32'sd134969, 32'sd662493, -32'sd884181, -32'sd215515, -32'sd2286166, 32'sd1313782, -32'sd199663, -32'sd934406, -32'sd139317, 32'sd544892, 32'sd2091983, 32'sd667736, -32'sd933798, 32'sd950028, 32'sd3042501, -32'sd1671535, 32'sd450776, 32'sd1689323, -32'sd973129, 32'sd0, 32'sd268915, 32'sd432151, 32'sd276049, 32'sd61202, 32'sd2532933, 32'sd607010, 32'sd385730, -32'sd1161619, -32'sd1192573, -32'sd932973, -32'sd1852585, -32'sd2576838, -32'sd1803263, -32'sd238306, 32'sd335456, 32'sd335974, 32'sd1739751, 32'sd344166, 32'sd1110483, 32'sd1656063, -32'sd1050422, 32'sd189415, 32'sd1731306, -32'sd1817400, 32'sd1492522, 32'sd1496296, 32'sd846855, 32'sd522276, -32'sd908962, -32'sd2050274, 32'sd534290, -32'sd684363, 32'sd305434, 32'sd188219, -32'sd2020348, -32'sd2087518, -32'sd1241019, -32'sd2564941, -32'sd454451, -32'sd800176, -32'sd435317, 32'sd446836, -32'sd197850, 32'sd1273455, 32'sd673670, -32'sd184708, 32'sd1888723, 32'sd1157712, 32'sd755319, -32'sd522470, 32'sd79486, 32'sd896156, 32'sd869465, -32'sd238030, 32'sd249370, -32'sd494316, -32'sd1253714, 32'sd1173782, -32'sd116382, 32'sd585665, -32'sd1046891, -32'sd1677201, -32'sd919232, -32'sd1024553, 32'sd957748, 32'sd787112, -32'sd606913, 32'sd150101, 32'sd874987, 32'sd1198088, 32'sd1348707, -32'sd389560, 32'sd2573369, 32'sd1177084, -32'sd34423, 32'sd2440396, 32'sd1617558, -32'sd1537419, 32'sd157652, 32'sd557490, 32'sd1366368, -32'sd1006596, -32'sd280576, 32'sd0, 32'sd433853, 32'sd371359, 32'sd630241, -32'sd161253, 32'sd700159, -32'sd468885, 32'sd874348, -32'sd1067059, -32'sd692023, -32'sd434702, 32'sd2781251, 32'sd1810723, 32'sd369081, -32'sd165755, -32'sd252798, -32'sd510650, 32'sd1413140, -32'sd875851, 32'sd555305, 32'sd2477556, 32'sd360970, -32'sd548807, -32'sd616255, -32'sd1334646, -32'sd561549, -32'sd102230, 32'sd0, 32'sd0, 32'sd0, 32'sd222231, -32'sd996100, -32'sd145731, -32'sd533943, -32'sd187958, -32'sd332526, 32'sd594550, 32'sd156969, 32'sd1242729, 32'sd875464, 32'sd2697933, 32'sd415318, -32'sd23253, 32'sd885940, 32'sd54383, 32'sd1076933, -32'sd160562, 32'sd844140, -32'sd2148461, -32'sd1602005, -32'sd714852, -32'sd463694, -32'sd815436, 32'sd27443, 32'sd863546, 32'sd0, 32'sd0, 32'sd0, 32'sd67288, -32'sd425854, -32'sd1634743, -32'sd1320636, 32'sd2176310, 32'sd526249, 32'sd559190, -32'sd408746, 32'sd402750, 32'sd1681908, 32'sd1689130, 32'sd121494, -32'sd1230335, 32'sd721605, 32'sd1495087, 32'sd1683375, -32'sd1720010, 32'sd39571, 32'sd23180, 32'sd813567, -32'sd57889, -32'sd544566, -32'sd1408753, 32'sd70999, -32'sd959745, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1462623, -32'sd1984676, 32'sd223060, 32'sd1390987, 32'sd107347, 32'sd2947479, 32'sd456485, 32'sd9478, 32'sd1313074, 32'sd1280172, 32'sd2066881, 32'sd722170, 32'sd3574420, 32'sd288795, 32'sd1251081, 32'sd1490025, 32'sd1446353, 32'sd471398, -32'sd1173106, -32'sd1807618, -32'sd137288, 32'sd1273119, 32'sd753581, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1598288, 32'sd107224, 32'sd1042576, 32'sd1416211, 32'sd1864633, 32'sd939631, 32'sd2251459, 32'sd398868, 32'sd673114, 32'sd1440022, 32'sd302748, 32'sd1106933, 32'sd1613830, 32'sd241107, -32'sd1153845, 32'sd129583, 32'sd912510, 32'sd759975, 32'sd1159771, 32'sd1108775, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1307657, -32'sd505847, -32'sd89882, -32'sd25812, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd137655, -32'sd1348323, 32'sd119988, -32'sd274668, -32'sd1053594, -32'sd382849, -32'sd1565103, 32'sd447956, -32'sd544510, 32'sd604844, -32'sd95959, -32'sd431357, 32'sd1631269, 32'sd1368284, -32'sd1288698, 32'sd87988, 32'sd531106, 32'sd966839, 32'sd1191415, 32'sd519753, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd335140, 32'sd250413, 32'sd1393749, -32'sd109779, 32'sd759903, 32'sd781182, -32'sd1015694, -32'sd644795, 32'sd728018, -32'sd764806, -32'sd1400552, 32'sd2200975, 32'sd724128, 32'sd853479, 32'sd1296564, -32'sd1043688, -32'sd58505, 32'sd445677, 32'sd1668160, 32'sd2139865, 32'sd658623, -32'sd804299, 32'sd1223366, 32'sd112599, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd311363, -32'sd357376, -32'sd1211398, -32'sd64394, 32'sd693474, -32'sd1042706, -32'sd755680, 32'sd1487825, 32'sd962366, 32'sd262805, 32'sd2345505, 32'sd4692642, 32'sd1900865, 32'sd1834981, 32'sd716283, 32'sd413547, -32'sd186198, -32'sd318366, 32'sd511549, -32'sd26969, -32'sd163132, -32'sd491493, 32'sd312796, -32'sd965232, -32'sd346741, 32'sd0, 32'sd0, 32'sd143592, 32'sd384427, -32'sd1082994, 32'sd1019791, 32'sd218877, -32'sd508910, -32'sd2414991, -32'sd1940332, 32'sd212106, 32'sd2285782, 32'sd933816, 32'sd1313970, 32'sd1228416, 32'sd578498, -32'sd1208924, -32'sd271185, 32'sd548585, 32'sd526491, 32'sd1619798, 32'sd996184, -32'sd1215576, 32'sd140914, 32'sd1684697, -32'sd114625, 32'sd502076, 32'sd169221, -32'sd182818, 32'sd0, 32'sd259567, -32'sd831696, -32'sd492809, 32'sd286308, -32'sd1957505, 32'sd88394, -32'sd876613, 32'sd251170, 32'sd1604394, 32'sd2076139, 32'sd803748, 32'sd1979535, 32'sd1536983, 32'sd3434878, 32'sd260679, 32'sd3149937, 32'sd1904709, 32'sd2706563, 32'sd1567610, -32'sd310954, -32'sd846541, 32'sd202960, -32'sd242110, 32'sd229269, 32'sd1607321, 32'sd433667, 32'sd29917, 32'sd0, 32'sd538258, -32'sd320730, -32'sd4402, -32'sd42769, -32'sd2057835, -32'sd1925754, 32'sd331405, -32'sd869083, 32'sd419941, -32'sd1301327, 32'sd1739253, 32'sd476277, 32'sd1729561, 32'sd2088307, -32'sd157532, 32'sd1391695, 32'sd174507, 32'sd599396, -32'sd515751, -32'sd213223, -32'sd1852264, 32'sd273253, -32'sd1106694, -32'sd1618960, -32'sd769661, 32'sd864449, 32'sd860833, 32'sd324140, 32'sd1287845, -32'sd903298, -32'sd628836, -32'sd401966, -32'sd1096759, -32'sd1433499, -32'sd1289334, 32'sd833989, -32'sd11289, 32'sd1262122, 32'sd975113, 32'sd721901, 32'sd789610, 32'sd233047, -32'sd199507, -32'sd971405, -32'sd1458663, -32'sd1908087, -32'sd1194960, -32'sd1449385, -32'sd1740821, -32'sd2741799, -32'sd1512049, -32'sd1978292, -32'sd702922, -32'sd21178, -32'sd940908, 32'sd876758, -32'sd131117, 32'sd737792, -32'sd279913, -32'sd1714230, -32'sd514840, 32'sd364183, -32'sd64057, 32'sd1883976, 32'sd1918523, 32'sd1617617, 32'sd1969681, 32'sd1389515, 32'sd28553, -32'sd260300, -32'sd2910811, -32'sd2634927, -32'sd451894, -32'sd2183880, -32'sd2988564, -32'sd1244275, -32'sd1584091, -32'sd1790021, -32'sd1231960, -32'sd1364116, -32'sd1170211, -32'sd73531, 32'sd1171701, 32'sd605341, 32'sd1265294, 32'sd70567, -32'sd1059044, -32'sd1201576, -32'sd344092, 32'sd1859088, 32'sd2063882, 32'sd2062426, 32'sd1245515, 32'sd602200, 32'sd921839, -32'sd687227, -32'sd756677, -32'sd1851841, -32'sd1509493, -32'sd4156960, -32'sd2245931, -32'sd128495, -32'sd1361010, -32'sd2756705, -32'sd440947, -32'sd1587929, -32'sd1777546, 32'sd1507897, -32'sd834925, 32'sd1078425, 32'sd1292488, 32'sd144148, 32'sd1211436, 32'sd1442440, -32'sd1977469, -32'sd2887666, -32'sd312131, -32'sd279836, -32'sd617032, 32'sd1346662, 32'sd199481, 32'sd7962, -32'sd7493, -32'sd1412469, -32'sd436375, -32'sd785319, -32'sd1827604, -32'sd2566408, -32'sd393334, -32'sd855354, 32'sd729729, 32'sd385680, 32'sd372521, 32'sd825538, 32'sd976343, 32'sd1668444, -32'sd576974, 32'sd504721, -32'sd491959, -32'sd447703, 32'sd56957, 32'sd182555, 32'sd362840, -32'sd1447227, -32'sd1561056, -32'sd783573, -32'sd727363, -32'sd1716696, -32'sd2000062, -32'sd1282277, -32'sd2321422, -32'sd3442797, -32'sd170443, 32'sd1104699, 32'sd1442974, 32'sd880699, -32'sd637102, 32'sd1551571, 32'sd1881655, 32'sd219446, 32'sd1401026, 32'sd1035898, 32'sd4222299, 32'sd1605242, 32'sd789285, 32'sd1245160, 32'sd1597829, 32'sd380082, -32'sd998235, -32'sd214655, 32'sd999086, -32'sd154988, -32'sd139848, -32'sd1045591, -32'sd547356, -32'sd1183390, -32'sd1670477, -32'sd1499167, -32'sd1088208, -32'sd1859442, -32'sd668036, 32'sd116245, 32'sd2308907, 32'sd553793, -32'sd1555344, -32'sd1018726, 32'sd1144436, -32'sd1146278, 32'sd276837, -32'sd699173, 32'sd2202015, 32'sd2058698, 32'sd785774, -32'sd735695, -32'sd11636, 32'sd287969, 32'sd230729, 32'sd519177, -32'sd947215, -32'sd2196380, 32'sd641321, -32'sd585546, 32'sd782531, -32'sd2252959, 32'sd742893, 32'sd799574, -32'sd649338, -32'sd2085070, -32'sd1189223, 32'sd2803176, -32'sd23915, -32'sd2344750, -32'sd2078495, -32'sd2547634, 32'sd268866, 32'sd303764, 32'sd127087, 32'sd224031, -32'sd139242, 32'sd1016015, 32'sd248751, -32'sd1966, 32'sd1222288, 32'sd777479, -32'sd675486, 32'sd712005, 32'sd952988, 32'sd1105713, 32'sd2402706, 32'sd148063, 32'sd178436, 32'sd272293, 32'sd154518, 32'sd1876112, -32'sd1000547, 32'sd336723, -32'sd1530599, 32'sd224124, -32'sd2094962, -32'sd2427796, -32'sd2568662, -32'sd1294721, -32'sd1043988, -32'sd574628, 32'sd21964, 32'sd1460854, 32'sd1270349, 32'sd1446092, 32'sd218359, -32'sd1192549, 32'sd953545, 32'sd1209537, -32'sd1162452, 32'sd578274, -32'sd1860689, 32'sd95902, 32'sd846231, 32'sd477262, -32'sd603695, -32'sd79950, 32'sd1019905, -32'sd333048, -32'sd968522, -32'sd1077502, 32'sd1383598, 32'sd368310, -32'sd2534793, -32'sd3426942, -32'sd1434603, -32'sd275961, 32'sd1686273, -32'sd847769, -32'sd594920, -32'sd231396, -32'sd482502, -32'sd1309660, -32'sd1405236, -32'sd333294, 32'sd674786, 32'sd507674, 32'sd960428, -32'sd1082506, -32'sd1825956, -32'sd666441, 32'sd1378570, 32'sd470390, -32'sd1298074, -32'sd2254475, -32'sd1296266, -32'sd848546, -32'sd3135360, -32'sd1031137, 32'sd1071373, 32'sd1982069, -32'sd1570549, -32'sd3780810, -32'sd1483734, 32'sd19384, 32'sd210114, -32'sd817449, 32'sd37609, -32'sd343207, -32'sd187991, -32'sd1430799, 32'sd252675, 32'sd685509, -32'sd322870, 32'sd0, -32'sd25501, 32'sd55548, -32'sd2412600, 32'sd1029597, -32'sd34140, 32'sd616145, -32'sd1452549, -32'sd436473, -32'sd1193478, -32'sd1942199, -32'sd1068922, -32'sd1322589, -32'sd908901, 32'sd2650903, 32'sd929814, -32'sd202706, 32'sd436944, -32'sd597947, 32'sd367570, 32'sd606488, -32'sd338661, 32'sd180635, -32'sd89283, -32'sd1135992, -32'sd432043, -32'sd756150, 32'sd389989, 32'sd605233, 32'sd840470, 32'sd657023, -32'sd1372235, -32'sd689901, 32'sd1206749, 32'sd1271550, -32'sd1444017, -32'sd936025, 32'sd281852, 32'sd181673, -32'sd3085254, -32'sd880332, 32'sd473427, 32'sd3273180, 32'sd84184, 32'sd697883, -32'sd280222, 32'sd630544, -32'sd1553594, -32'sd425507, -32'sd529687, 32'sd763651, -32'sd99000, 32'sd2329249, -32'sd523730, -32'sd1217708, -32'sd268167, 32'sd528628, 32'sd1183614, -32'sd1986135, -32'sd1172480, -32'sd1940566, 32'sd1405147, 32'sd1487073, 32'sd985688, 32'sd410614, -32'sd193075, -32'sd300875, 32'sd729793, 32'sd743846, 32'sd3522937, 32'sd3476833, 32'sd775514, -32'sd716715, -32'sd651844, -32'sd1544493, -32'sd1167320, 32'sd645087, -32'sd1102190, 32'sd348228, -32'sd252891, -32'sd368035, 32'sd388835, -32'sd1990875, -32'sd115680, 32'sd0, 32'sd170038, -32'sd381206, -32'sd927646, -32'sd43513, 32'sd2107896, 32'sd678312, -32'sd1253871, -32'sd2555876, -32'sd764590, -32'sd1405549, 32'sd1811122, 32'sd2752876, 32'sd3171555, 32'sd925896, 32'sd2794909, 32'sd716067, -32'sd1702017, 32'sd289143, -32'sd5347, -32'sd1283222, -32'sd1913369, -32'sd80156, -32'sd484461, 32'sd134395, -32'sd1595434, -32'sd1533765, 32'sd129356, -32'sd58952, -32'sd1211369, 32'sd900001, 32'sd769621, 32'sd421316, 32'sd785217, 32'sd1959604, -32'sd1101740, -32'sd1932869, -32'sd2532859, -32'sd41366, 32'sd840135, 32'sd2162711, 32'sd1889126, 32'sd1504134, 32'sd2533463, -32'sd278460, -32'sd58398, 32'sd207386, -32'sd472187, 32'sd518760, 32'sd510586, 32'sd52708, -32'sd441391, 32'sd1012677, -32'sd1767472, 32'sd718568, 32'sd456720, 32'sd1858549, 32'sd1198800, -32'sd2155607, -32'sd728587, 32'sd132666, -32'sd1447026, 32'sd902166, 32'sd1075791, 32'sd529233, 32'sd460872, 32'sd795206, 32'sd159261, -32'sd1061794, -32'sd131644, 32'sd1531173, 32'sd1872957, 32'sd2064511, 32'sd325447, 32'sd1138619, -32'sd1264277, 32'sd633115, -32'sd183186, 32'sd1150232, -32'sd232364, 32'sd1965148, -32'sd1784813, -32'sd300282, 32'sd430646, 32'sd0, 32'sd6295, 32'sd585104, -32'sd578381, -32'sd788563, 32'sd1024898, 32'sd1019236, -32'sd164982, 32'sd256375, 32'sd685944, 32'sd473024, -32'sd460604, -32'sd810501, -32'sd764172, 32'sd1045522, 32'sd1535967, 32'sd1829102, 32'sd1682127, -32'sd2448408, -32'sd1269775, 32'sd1688098, -32'sd414395, 32'sd1177962, -32'sd731201, 32'sd501600, -32'sd1021777, -32'sd400700, 32'sd0, 32'sd0, 32'sd0, -32'sd112158, -32'sd357374, -32'sd1767982, -32'sd440285, -32'sd2998, -32'sd690814, 32'sd587416, -32'sd440883, -32'sd1298750, 32'sd1535366, -32'sd277782, 32'sd334939, -32'sd1457998, -32'sd769318, 32'sd1005515, 32'sd1763526, 32'sd1819585, 32'sd793881, 32'sd1461271, -32'sd856427, -32'sd180185, 32'sd594609, 32'sd1160267, 32'sd272832, -32'sd844124, 32'sd0, 32'sd0, 32'sd0, -32'sd842359, 32'sd1765057, 32'sd101921, 32'sd249761, 32'sd965263, 32'sd1780198, -32'sd1675399, -32'sd1840709, -32'sd2537317, -32'sd130235, -32'sd164812, -32'sd173618, -32'sd173026, -32'sd946865, 32'sd359954, 32'sd1640753, 32'sd1682971, -32'sd544789, 32'sd930694, 32'sd790793, 32'sd222767, 32'sd786920, 32'sd1277125, 32'sd810912, 32'sd435101, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd905738, 32'sd472360, 32'sd315306, 32'sd309033, 32'sd1201024, 32'sd2074872, 32'sd230848, 32'sd481026, 32'sd912114, -32'sd1778164, -32'sd1178439, 32'sd795039, 32'sd1756800, 32'sd132877, -32'sd2278568, -32'sd58017, -32'sd988054, 32'sd620667, -32'sd2111167, -32'sd1232336, 32'sd286440, 32'sd1284047, 32'sd70874, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd219940, 32'sd697875, 32'sd1439029, -32'sd1049398, 32'sd832126, -32'sd275510, 32'sd763554, 32'sd1034593, 32'sd720284, 32'sd872227, -32'sd666921, 32'sd769329, 32'sd613828, 32'sd873006, -32'sd633897, 32'sd238668, -32'sd457895, -32'sd1050033, -32'sd997416, 32'sd799866, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd602898, -32'sd1083024, 32'sd424221, -32'sd1053810, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1157151, 32'sd486324, -32'sd506013, -32'sd686522, -32'sd626817, 32'sd236907, 32'sd854668, -32'sd331152, -32'sd34213, 32'sd275032, 32'sd1109224, -32'sd693276, -32'sd1377725, 32'sd483422, -32'sd1202489, 32'sd547688, -32'sd388577, 32'sd49997, -32'sd1134340, 32'sd248939, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd34342, -32'sd350989, 32'sd1909626, -32'sd27062, -32'sd399775, -32'sd1106136, 32'sd885135, 32'sd1486566, 32'sd790237, 32'sd429851, -32'sd257703, -32'sd418988, -32'sd1019120, -32'sd1071597, -32'sd1508304, -32'sd992789, 32'sd82799, -32'sd458771, 32'sd570669, -32'sd476292, -32'sd174300, 32'sd657632, -32'sd775328, 32'sd486136, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd347043, -32'sd175923, -32'sd461952, -32'sd1027185, -32'sd1227908, 32'sd675293, -32'sd228174, -32'sd743388, -32'sd1765050, 32'sd177496, -32'sd560456, -32'sd70201, 32'sd2478619, -32'sd265757, -32'sd2806035, -32'sd838747, -32'sd1882938, -32'sd1292204, -32'sd1240631, 32'sd1022433, -32'sd383036, 32'sd319253, -32'sd4248, -32'sd811845, 32'sd1058831, 32'sd0, 32'sd0, -32'sd111546, -32'sd390823, 32'sd228121, -32'sd2905646, 32'sd343671, 32'sd83731, -32'sd507638, -32'sd237542, -32'sd2511299, -32'sd1407867, 32'sd47155, -32'sd18034, -32'sd1006034, -32'sd1868115, -32'sd2466856, -32'sd378319, -32'sd1021732, 32'sd878888, -32'sd908332, -32'sd248060, 32'sd2071052, 32'sd2286084, 32'sd497390, -32'sd696275, 32'sd139797, 32'sd598100, 32'sd896393, 32'sd0, 32'sd413824, -32'sd786853, 32'sd630149, 32'sd1278663, 32'sd212859, 32'sd978434, 32'sd1655748, 32'sd1503723, -32'sd540708, 32'sd665594, 32'sd725944, 32'sd1128785, 32'sd427318, -32'sd610488, -32'sd1825345, -32'sd1528310, -32'sd466136, -32'sd773748, -32'sd1215056, -32'sd1609549, 32'sd192189, 32'sd1050428, 32'sd435095, -32'sd1132645, 32'sd1678147, -32'sd694346, -32'sd1248804, 32'sd0, -32'sd45249, -32'sd1973152, 32'sd789050, 32'sd1583475, 32'sd589655, -32'sd302534, 32'sd1063447, 32'sd768829, -32'sd2367392, -32'sd731369, 32'sd330258, -32'sd625770, -32'sd578505, -32'sd805944, 32'sd539914, 32'sd1164097, 32'sd840342, -32'sd469600, 32'sd780100, 32'sd1068894, -32'sd43224, -32'sd112394, 32'sd2557857, 32'sd886502, -32'sd185163, 32'sd1549626, -32'sd38773, 32'sd427831, -32'sd442696, -32'sd973151, 32'sd259752, -32'sd490985, 32'sd60109, -32'sd1440270, -32'sd1905423, -32'sd1660494, -32'sd3333721, 32'sd136709, -32'sd511031, -32'sd988449, -32'sd731709, 32'sd1303578, 32'sd1027524, 32'sd1635339, 32'sd912547, -32'sd1094772, 32'sd2631378, 32'sd143719, 32'sd806431, 32'sd593120, 32'sd2462525, 32'sd991475, 32'sd1006705, -32'sd821173, -32'sd266892, 32'sd1024679, 32'sd184961, 32'sd80658, 32'sd1660133, -32'sd2341203, -32'sd625228, -32'sd1263219, -32'sd1039186, -32'sd1816772, 32'sd583196, 32'sd864172, 32'sd1400, 32'sd2187187, 32'sd1722401, -32'sd340856, -32'sd331772, -32'sd2631605, -32'sd1859556, 32'sd250123, -32'sd881509, 32'sd865146, 32'sd131128, 32'sd662126, -32'sd859422, 32'sd2166107, 32'sd1574394, 32'sd213125, 32'sd1227497, 32'sd682101, 32'sd116894, 32'sd6653, -32'sd1340156, -32'sd2798536, -32'sd445322, -32'sd146903, -32'sd2334832, -32'sd2016256, -32'sd900514, 32'sd607643, 32'sd985662, 32'sd3045597, 32'sd577965, -32'sd1621375, -32'sd906333, -32'sd1190822, -32'sd732327, -32'sd1492866, 32'sd1387092, 32'sd1031071, 32'sd302774, 32'sd215795, -32'sd886969, 32'sd949813, 32'sd530368, -32'sd14830, -32'sd486016, -32'sd263010, -32'sd201707, -32'sd1068873, 32'sd911451, -32'sd2314704, 32'sd904975, -32'sd925601, -32'sd1902878, -32'sd2425900, -32'sd577363, 32'sd445598, 32'sd2237709, 32'sd1052862, -32'sd2843150, -32'sd3262318, -32'sd3334334, -32'sd2599623, -32'sd1741858, -32'sd1830618, 32'sd1407406, 32'sd1102626, 32'sd94340, 32'sd1996270, 32'sd1931785, -32'sd456895, 32'sd1292490, -32'sd1164918, 32'sd409992, -32'sd590862, -32'sd1050443, 32'sd1812446, 32'sd212589, -32'sd1082922, -32'sd156500, -32'sd2011181, -32'sd1495342, -32'sd1212, 32'sd2462615, 32'sd2625262, -32'sd315816, -32'sd1042285, -32'sd4260192, -32'sd2500714, -32'sd2286184, -32'sd218480, 32'sd513011, -32'sd1103817, 32'sd364494, 32'sd1956166, 32'sd2035064, 32'sd1195145, 32'sd2292473, 32'sd817637, 32'sd539257, -32'sd1654858, -32'sd2081772, 32'sd654776, -32'sd1170044, 32'sd1136501, 32'sd961425, 32'sd541266, -32'sd278581, -32'sd1650018, -32'sd1591040, 32'sd1579442, 32'sd1086731, 32'sd2311615, -32'sd2036657, -32'sd2239433, -32'sd1451870, -32'sd1994567, -32'sd335598, 32'sd3260493, 32'sd214248, 32'sd683316, 32'sd2412437, 32'sd3437582, 32'sd3249964, 32'sd1645390, 32'sd1544345, 32'sd1522463, -32'sd1896750, -32'sd1155570, 32'sd126182, -32'sd23392, -32'sd121999, -32'sd546026, -32'sd1388750, -32'sd809448, -32'sd2401917, -32'sd675516, 32'sd1068656, 32'sd1088524, 32'sd1670170, -32'sd1277396, -32'sd391565, 32'sd761250, 32'sd65395, 32'sd2190464, 32'sd4927156, 32'sd1194937, 32'sd832398, 32'sd145764, 32'sd833213, 32'sd1726530, 32'sd2122475, 32'sd716413, 32'sd1216614, -32'sd461989, -32'sd1793624, -32'sd1951010, 32'sd567279, 32'sd745437, 32'sd623464, -32'sd123699, -32'sd795782, -32'sd201422, -32'sd778487, -32'sd3098171, 32'sd905457, -32'sd658656, -32'sd367466, -32'sd1274915, -32'sd537141, 32'sd541610, 32'sd4625823, 32'sd3295862, 32'sd3129770, 32'sd2677812, 32'sd1139514, -32'sd375071, 32'sd235123, 32'sd1305637, 32'sd375558, -32'sd1058241, -32'sd608360, -32'sd2074426, 32'sd676544, -32'sd644227, -32'sd440281, 32'sd467646, 32'sd1018496, -32'sd821439, 32'sd367082, -32'sd1347000, -32'sd1290233, -32'sd840926, 32'sd139635, 32'sd711123, -32'sd1325016, -32'sd291548, 32'sd1392572, 32'sd1525583, 32'sd2092882, 32'sd4824255, 32'sd2992617, 32'sd2548792, 32'sd524694, 32'sd654446, -32'sd2428420, -32'sd2391261, -32'sd365374, 32'sd525295, 32'sd698164, -32'sd697154, -32'sd1218802, 32'sd1058329, 32'sd935001, 32'sd8088, 32'sd1102365, -32'sd512161, 32'sd481207, 32'sd1204099, -32'sd553817, -32'sd1070625, 32'sd538735, 32'sd651205, -32'sd302462, 32'sd959362, 32'sd572341, 32'sd3379443, 32'sd3688595, 32'sd1837721, 32'sd309899, -32'sd173379, -32'sd962291, -32'sd1803878, -32'sd2068386, -32'sd71780, 32'sd346202, -32'sd975552, 32'sd1267248, 32'sd1279830, -32'sd1325284, 32'sd288238, 32'sd1367923, 32'sd0, -32'sd399700, -32'sd1629414, -32'sd146692, 32'sd493991, -32'sd2814081, -32'sd2319666, 32'sd347038, 32'sd339968, -32'sd3115460, -32'sd429469, 32'sd1244091, 32'sd1559529, 32'sd2690706, 32'sd766286, -32'sd277966, -32'sd957636, -32'sd2209339, -32'sd2367947, -32'sd600533, -32'sd1994848, -32'sd274996, 32'sd60283, -32'sd1054099, -32'sd2465650, -32'sd96712, -32'sd1181486, -32'sd1737626, 32'sd44468, 32'sd839813, -32'sd1149041, -32'sd2206527, -32'sd1237726, -32'sd1992122, -32'sd1813082, -32'sd138608, -32'sd1441010, 32'sd227908, -32'sd263480, 32'sd1645267, -32'sd603459, 32'sd409783, 32'sd1628965, 32'sd1102308, -32'sd2082610, -32'sd3134294, -32'sd1789414, -32'sd722273, -32'sd1700028, -32'sd1619810, -32'sd1665206, -32'sd834783, -32'sd1110597, 32'sd66035, 32'sd599443, 32'sd1119454, 32'sd197414, -32'sd781648, 32'sd1463273, -32'sd371103, 32'sd64238, -32'sd1104909, -32'sd958479, -32'sd356772, -32'sd1466183, 32'sd380084, 32'sd267280, -32'sd1340756, -32'sd822518, 32'sd970016, 32'sd3964787, -32'sd437708, -32'sd1689359, -32'sd315494, 32'sd142803, 32'sd935572, -32'sd1148320, 32'sd737268, -32'sd457677, -32'sd2514836, -32'sd376291, -32'sd567973, 32'sd1327559, 32'sd146721, 32'sd0, 32'sd786440, 32'sd1746231, -32'sd946625, 32'sd327794, 32'sd86066, -32'sd443454, 32'sd666376, -32'sd828806, -32'sd1896227, -32'sd520757, -32'sd2407166, 32'sd163795, 32'sd2119096, 32'sd3382191, 32'sd1332298, -32'sd1102977, 32'sd68516, -32'sd87537, -32'sd844582, -32'sd514209, 32'sd72146, -32'sd818528, -32'sd140937, -32'sd612349, 32'sd1172849, 32'sd1372732, -32'sd683873, 32'sd16393, 32'sd32958, -32'sd136173, 32'sd1206340, -32'sd241273, -32'sd986137, 32'sd1029499, 32'sd17359, -32'sd1898733, 32'sd264915, -32'sd262327, -32'sd313514, 32'sd678604, 32'sd621755, 32'sd238548, -32'sd374793, -32'sd2176942, -32'sd3985583, -32'sd533568, -32'sd1894297, -32'sd622344, -32'sd1058935, -32'sd882319, 32'sd898576, -32'sd1766606, -32'sd886224, 32'sd71568, 32'sd223053, 32'sd1454721, 32'sd81874, -32'sd545887, -32'sd1807347, 32'sd3072, -32'sd579051, 32'sd2819562, 32'sd1606924, -32'sd501642, -32'sd1148454, 32'sd515171, 32'sd89155, -32'sd163244, -32'sd801229, 32'sd1546489, -32'sd3075180, -32'sd5059838, -32'sd6069623, -32'sd1740852, -32'sd109323, -32'sd986700, -32'sd462698, -32'sd774024, -32'sd564964, -32'sd104777, -32'sd30064, -32'sd601852, 32'sd348944, 32'sd0, 32'sd58370, -32'sd362319, 32'sd648663, -32'sd2013333, 32'sd1433126, 32'sd360720, 32'sd785390, 32'sd2792127, -32'sd546032, 32'sd1177332, 32'sd1269307, -32'sd1399897, -32'sd1494557, 32'sd149161, -32'sd4163833, -32'sd3743347, -32'sd4026727, -32'sd197511, -32'sd2806072, -32'sd1406924, -32'sd756350, -32'sd1400022, 32'sd301358, 32'sd546395, 32'sd303927, 32'sd100627, 32'sd0, 32'sd0, 32'sd0, 32'sd1420079, -32'sd2402828, -32'sd939208, 32'sd581352, -32'sd123405, -32'sd930142, 32'sd1240003, 32'sd633694, 32'sd951303, -32'sd513464, 32'sd179794, 32'sd402343, 32'sd2806648, 32'sd908379, -32'sd1277513, -32'sd3900720, 32'sd244961, -32'sd770177, -32'sd546525, 32'sd914036, 32'sd1187456, 32'sd1555959, 32'sd832927, 32'sd29558, 32'sd811904, 32'sd0, 32'sd0, 32'sd0, 32'sd924973, -32'sd1832528, -32'sd327138, 32'sd513902, -32'sd185015, 32'sd943112, 32'sd358313, -32'sd348581, -32'sd346633, 32'sd764909, -32'sd1012976, 32'sd401163, 32'sd177458, -32'sd387101, -32'sd583137, -32'sd1920820, 32'sd1497749, 32'sd471590, -32'sd1072517, -32'sd2259921, 32'sd470889, 32'sd511635, -32'sd1081665, 32'sd657344, -32'sd21884, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd630351, 32'sd478921, 32'sd1020582, -32'sd439539, -32'sd70625, 32'sd458098, 32'sd383308, 32'sd1170598, 32'sd2067607, 32'sd1794403, 32'sd2005601, 32'sd1072554, -32'sd295497, 32'sd344805, 32'sd912224, 32'sd2414037, 32'sd43045, 32'sd718726, -32'sd699686, 32'sd633206, 32'sd87048, 32'sd924019, 32'sd867501, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd511654, 32'sd916342, 32'sd180529, 32'sd59304, 32'sd416429, -32'sd43843, 32'sd389636, 32'sd160685, 32'sd1000112, 32'sd182801, 32'sd1022298, 32'sd1023679, 32'sd2301305, 32'sd154071, 32'sd2277261, -32'sd35348, -32'sd466738, 32'sd244579, 32'sd194405, 32'sd94898, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1340798, 32'sd993668, 32'sd1351688, -32'sd468219, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd132098, 32'sd901119, -32'sd531107, 32'sd560848, 32'sd3807, 32'sd1419432, -32'sd855464, -32'sd806471, -32'sd281040, 32'sd148654, -32'sd316159, -32'sd149220, 32'sd1677447, 32'sd1689423, 32'sd1551205, 32'sd250768, 32'sd1635923, 32'sd2209046, 32'sd1160177, 32'sd719766, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1333675, 32'sd824275, -32'sd1609875, 32'sd229981, 32'sd636868, 32'sd1268749, 32'sd464396, -32'sd803566, 32'sd424455, -32'sd172708, -32'sd740410, -32'sd1254477, 32'sd1736035, 32'sd1276187, 32'sd761461, 32'sd1094936, -32'sd425171, -32'sd1015864, 32'sd433069, 32'sd2513985, 32'sd1455953, 32'sd1456638, 32'sd2218556, 32'sd1189290, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd322592, 32'sd1357615, 32'sd1085406, 32'sd542697, -32'sd843732, -32'sd7348, 32'sd1591487, 32'sd1771177, 32'sd333692, 32'sd1914736, 32'sd863525, 32'sd472441, 32'sd244420, 32'sd592581, 32'sd539227, -32'sd75061, 32'sd458921, -32'sd1187827, -32'sd1616879, -32'sd222727, -32'sd81008, 32'sd34815, 32'sd1949666, 32'sd352703, 32'sd34031, 32'sd0, 32'sd0, 32'sd823892, -32'sd280751, 32'sd426185, 32'sd1179245, 32'sd411318, 32'sd380314, -32'sd301844, 32'sd1340967, -32'sd884663, -32'sd622730, 32'sd1698797, 32'sd1393541, 32'sd87649, 32'sd286719, 32'sd51047, 32'sd68190, -32'sd658178, -32'sd97630, 32'sd1235282, -32'sd37787, -32'sd599735, -32'sd1093354, -32'sd1376650, -32'sd665260, 32'sd27273, 32'sd734860, 32'sd1250237, 32'sd0, 32'sd1264324, -32'sd291286, -32'sd881814, 32'sd336151, -32'sd1048386, 32'sd2138202, 32'sd1724415, 32'sd1892168, 32'sd299693, 32'sd3292036, 32'sd3526135, 32'sd2121909, 32'sd1013352, -32'sd946095, -32'sd2141492, 32'sd91874, -32'sd1256472, -32'sd298867, 32'sd805109, 32'sd1223629, 32'sd351137, -32'sd1231851, -32'sd655160, -32'sd2845366, -32'sd1708949, -32'sd354401, -32'sd55862, 32'sd0, 32'sd945151, -32'sd229777, -32'sd226419, -32'sd1295395, 32'sd606185, 32'sd384003, -32'sd56550, 32'sd1667165, 32'sd3715490, 32'sd3192690, 32'sd3540386, 32'sd1066582, 32'sd1651639, 32'sd890782, 32'sd2239323, 32'sd2066921, 32'sd427375, -32'sd703448, 32'sd941071, -32'sd379191, 32'sd399973, 32'sd652674, -32'sd157518, 32'sd167483, -32'sd60127, 32'sd752261, -32'sd1437400, 32'sd2166887, 32'sd340318, -32'sd354264, 32'sd1074881, -32'sd16499, -32'sd797211, 32'sd1109912, 32'sd2298985, -32'sd943026, 32'sd1109418, 32'sd1972248, 32'sd2529065, 32'sd2711870, 32'sd2482125, 32'sd2750063, 32'sd548404, 32'sd1548057, 32'sd1241168, 32'sd489491, 32'sd2788249, 32'sd1831369, 32'sd541178, -32'sd1082885, -32'sd249833, 32'sd2094186, 32'sd1550485, 32'sd2442808, -32'sd312618, 32'sd769494, 32'sd1195738, -32'sd1851865, 32'sd1413441, -32'sd444138, -32'sd314862, -32'sd1168443, 32'sd331168, -32'sd619212, -32'sd1613410, -32'sd1070988, 32'sd836524, -32'sd635675, 32'sd413100, 32'sd2092846, 32'sd1122608, 32'sd619783, 32'sd309725, 32'sd722785, 32'sd1305116, 32'sd46706, 32'sd538554, 32'sd144224, 32'sd799252, 32'sd483656, -32'sd546147, 32'sd1257908, -32'sd877459, 32'sd572270, -32'sd1924079, -32'sd1330754, 32'sd200342, 32'sd351799, -32'sd357883, -32'sd1913992, 32'sd1655800, -32'sd2242589, -32'sd2993122, -32'sd4220646, -32'sd1991816, -32'sd2962330, -32'sd3324924, -32'sd3348739, -32'sd1071749, -32'sd317863, 32'sd196345, 32'sd1119009, 32'sd1611602, 32'sd883468, -32'sd287870, 32'sd1926023, 32'sd1120589, -32'sd2002768, 32'sd348789, 32'sd523315, 32'sd962266, -32'sd533110, 32'sd315079, -32'sd394237, -32'sd815007, 32'sd843899, -32'sd1418389, -32'sd883547, -32'sd1397588, -32'sd2328941, -32'sd3095689, -32'sd5356843, -32'sd5541261, -32'sd3315053, -32'sd5649523, -32'sd3934369, -32'sd3262961, -32'sd355665, 32'sd1229257, 32'sd1130416, 32'sd1334982, 32'sd530040, -32'sd313429, 32'sd90357, -32'sd1016607, 32'sd840025, -32'sd321833, 32'sd2169448, 32'sd344693, -32'sd447718, -32'sd127041, -32'sd336859, -32'sd816532, -32'sd605682, -32'sd1596281, -32'sd2382476, -32'sd3753427, -32'sd5333534, -32'sd4366056, -32'sd5565312, -32'sd6070275, -32'sd7041733, -32'sd4726502, -32'sd3159139, -32'sd2656663, -32'sd714042, -32'sd152938, 32'sd825543, -32'sd939726, -32'sd453392, 32'sd69630, -32'sd584667, -32'sd473693, 32'sd462497, -32'sd240561, -32'sd790264, -32'sd883149, 32'sd745177, -32'sd438311, -32'sd1770342, -32'sd913798, -32'sd2783351, -32'sd4774384, -32'sd3657906, -32'sd4326716, -32'sd4427089, -32'sd3982265, -32'sd2584934, -32'sd3797133, -32'sd2246435, -32'sd288492, -32'sd1277268, 32'sd976591, -32'sd1451841, -32'sd1294054, -32'sd446392, -32'sd839272, 32'sd154491, 32'sd368502, -32'sd3412869, 32'sd1392911, 32'sd304121, -32'sd161702, -32'sd1772462, 32'sd659544, 32'sd1394722, 32'sd100813, -32'sd131445, -32'sd2105931, -32'sd1865110, -32'sd2822689, -32'sd4891107, -32'sd4417191, -32'sd2869265, -32'sd795032, -32'sd2010365, -32'sd1914605, -32'sd655632, 32'sd3466643, 32'sd791451, 32'sd245242, -32'sd1948733, -32'sd2768147, -32'sd125810, -32'sd43046, -32'sd332866, -32'sd914908, -32'sd2127166, -32'sd720574, 32'sd95120, -32'sd304306, 32'sd459479, 32'sd102001, 32'sd380399, -32'sd111341, -32'sd164780, -32'sd1425416, -32'sd842454, -32'sd584883, 32'sd1213163, -32'sd765994, 32'sd1803649, 32'sd3007791, 32'sd2392626, 32'sd589386, 32'sd2914520, 32'sd3641896, 32'sd324249, -32'sd55680, -32'sd1878312, -32'sd1382771, 32'sd548922, 32'sd204674, 32'sd259405, -32'sd261118, 32'sd707847, -32'sd743237, 32'sd1474192, 32'sd413161, 32'sd529764, -32'sd1173533, -32'sd269231, -32'sd1529345, -32'sd131574, 32'sd5273, -32'sd922957, 32'sd1742583, 32'sd2645601, 32'sd3136001, 32'sd2889618, 32'sd2036869, 32'sd1363691, 32'sd906369, 32'sd505030, 32'sd1677924, -32'sd532265, -32'sd251175, -32'sd683393, 32'sd1135839, 32'sd471656, -32'sd1139761, -32'sd255708, -32'sd412898, -32'sd1081258, 32'sd1883019, 32'sd706602, -32'sd484139, -32'sd727479, 32'sd1739610, 32'sd954356, -32'sd315620, 32'sd956846, -32'sd580635, 32'sd1223508, 32'sd2397328, 32'sd2973223, 32'sd3151712, 32'sd2847926, 32'sd3196252, 32'sd492051, 32'sd1871797, 32'sd217595, -32'sd239364, -32'sd225095, -32'sd546470, 32'sd313724, -32'sd671345, 32'sd71782, 32'sd891952, -32'sd552427, -32'sd717491, -32'sd540660, -32'sd160971, -32'sd872056, -32'sd592657, -32'sd807910, 32'sd2815348, 32'sd0, 32'sd140480, -32'sd325644, -32'sd23648, 32'sd225751, 32'sd2369932, 32'sd3403048, 32'sd1670769, 32'sd724224, -32'sd315404, -32'sd1744030, -32'sd1029134, 32'sd2450187, 32'sd1498024, 32'sd924253, -32'sd40526, -32'sd811889, -32'sd671550, -32'sd2546491, 32'sd970394, 32'sd118204, -32'sd1386156, -32'sd1340438, 32'sd687269, 32'sd1665729, -32'sd426303, -32'sd188646, -32'sd418495, 32'sd538229, 32'sd1661180, -32'sd99173, 32'sd2123113, 32'sd509629, 32'sd2455881, 32'sd1254022, 32'sd194103, -32'sd1618800, -32'sd1647581, -32'sd2158619, -32'sd948150, 32'sd1804659, 32'sd2298486, -32'sd1451138, 32'sd1151526, -32'sd1050725, 32'sd1172290, -32'sd616436, 32'sd1149952, 32'sd1027627, 32'sd640686, -32'sd893786, 32'sd2131648, 32'sd30152, -32'sd1995478, 32'sd266039, -32'sd589428, 32'sd1293904, 32'sd1277200, 32'sd593678, 32'sd950601, -32'sd897714, 32'sd1084024, -32'sd1842882, -32'sd1513910, -32'sd1461267, -32'sd1267747, -32'sd1393200, 32'sd973202, -32'sd126791, 32'sd2027216, -32'sd870715, -32'sd1503151, 32'sd1175000, 32'sd759346, 32'sd318499, 32'sd1412285, 32'sd1731059, -32'sd501840, 32'sd1079259, 32'sd253043, -32'sd982429, 32'sd2277411, 32'sd1657784, 32'sd721139, 32'sd0, 32'sd84015, 32'sd1244998, -32'sd163089, -32'sd999102, 32'sd33490, 32'sd982056, 32'sd104668, 32'sd118484, -32'sd2026525, 32'sd1475749, -32'sd334428, 32'sd379585, -32'sd1180540, -32'sd168629, 32'sd950820, -32'sd403093, 32'sd322829, 32'sd1346305, -32'sd721426, 32'sd724219, -32'sd345740, 32'sd512371, 32'sd758004, 32'sd586704, 32'sd918349, 32'sd1533677, 32'sd236948, 32'sd38324, 32'sd351650, 32'sd1627224, 32'sd326735, 32'sd172567, -32'sd323514, 32'sd106633, -32'sd293871, 32'sd223777, -32'sd1384920, 32'sd119621, -32'sd1712405, 32'sd1220535, 32'sd1072206, 32'sd1767376, 32'sd495087, -32'sd906841, -32'sd609727, 32'sd149281, 32'sd2623945, -32'sd324096, 32'sd1669693, 32'sd101031, 32'sd98482, 32'sd914772, 32'sd2178333, 32'sd111978, 32'sd32834, -32'sd863529, 32'sd573097, 32'sd2017158, 32'sd1180878, 32'sd463703, 32'sd1594886, 32'sd816881, 32'sd12832, 32'sd1024929, -32'sd210472, -32'sd493034, 32'sd32967, -32'sd542052, 32'sd282316, -32'sd1924334, -32'sd1376761, -32'sd196748, 32'sd1117263, 32'sd397631, -32'sd730143, 32'sd1078242, 32'sd125490, -32'sd2454548, -32'sd1169381, 32'sd181927, 32'sd332654, 32'sd1284819, 32'sd1584153, 32'sd0, 32'sd1054662, -32'sd239593, 32'sd498782, 32'sd106169, 32'sd550141, -32'sd1001893, 32'sd1564516, 32'sd606961, -32'sd10447, -32'sd664899, -32'sd802, -32'sd1161738, -32'sd204839, -32'sd501516, -32'sd1196801, -32'sd1939685, -32'sd3076397, -32'sd2100920, -32'sd1322667, -32'sd629119, 32'sd312322, -32'sd908418, -32'sd666346, 32'sd522787, 32'sd1327448, -32'sd389518, 32'sd0, 32'sd0, 32'sd0, -32'sd1496244, 32'sd338452, 32'sd694287, 32'sd305794, -32'sd1031116, 32'sd383651, 32'sd2574265, 32'sd1027772, 32'sd927096, 32'sd2025774, 32'sd778767, -32'sd420087, 32'sd2559580, -32'sd952533, -32'sd2028025, -32'sd804194, -32'sd409889, 32'sd587011, -32'sd361330, 32'sd60922, 32'sd1718196, -32'sd615916, 32'sd1350278, 32'sd251826, -32'sd82711, 32'sd0, 32'sd0, 32'sd0, 32'sd424639, 32'sd1137674, 32'sd212734, -32'sd721487, 32'sd983445, 32'sd504356, -32'sd251143, -32'sd377443, 32'sd951388, -32'sd140935, 32'sd2129576, -32'sd1636614, 32'sd514520, 32'sd1768242, -32'sd1796796, 32'sd817380, -32'sd3045387, -32'sd1173410, -32'sd1235564, 32'sd245118, 32'sd682854, 32'sd35921, -32'sd1454998, 32'sd809897, 32'sd625235, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1110759, 32'sd22263, 32'sd630765, -32'sd233660, -32'sd1100148, -32'sd1027136, 32'sd482684, 32'sd1429230, 32'sd1924603, 32'sd423890, 32'sd1064948, 32'sd932993, -32'sd798282, 32'sd773287, -32'sd109606, 32'sd1900767, -32'sd166490, -32'sd160880, -32'sd1348029, -32'sd568888, 32'sd1789277, -32'sd188673, 32'sd2062279, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2437007, 32'sd655007, 32'sd1835695, 32'sd1558274, 32'sd2487788, 32'sd1027170, 32'sd545803, 32'sd1805401, 32'sd2973698, 32'sd1831822, 32'sd1357894, 32'sd2068926, 32'sd1061744, 32'sd982424, 32'sd490685, -32'sd447906, 32'sd769531, 32'sd525432, -32'sd944709, 32'sd2773592, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd625037, -32'sd691637, 32'sd277785, -32'sd613359, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd303998, 32'sd793684, 32'sd36852, 32'sd13636, 32'sd939326, 32'sd1633167, 32'sd729666, 32'sd1660980, 32'sd1138789, -32'sd887888, -32'sd211612, 32'sd411947, 32'sd1305457, -32'sd579422, 32'sd779322, 32'sd803433, 32'sd476404, -32'sd110335, 32'sd639614, -32'sd122914, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd952592, -32'sd708326, -32'sd1328403, -32'sd746770, 32'sd1509996, 32'sd418844, 32'sd187176, -32'sd337177, -32'sd121922, 32'sd177931, 32'sd1983690, 32'sd1535755, 32'sd1407827, 32'sd1253721, 32'sd1132478, -32'sd706516, -32'sd504359, 32'sd356172, 32'sd818677, -32'sd583386, -32'sd1186861, 32'sd1424378, -32'sd455024, 32'sd363895, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd709282, 32'sd357647, 32'sd242893, 32'sd660988, -32'sd101802, -32'sd1624141, -32'sd2229846, 32'sd1425782, 32'sd490857, -32'sd400754, 32'sd1506129, 32'sd314414, 32'sd58345, 32'sd755687, 32'sd3471096, 32'sd1042190, 32'sd1169729, 32'sd253688, -32'sd217825, -32'sd259950, -32'sd211373, -32'sd1430530, -32'sd930030, 32'sd1128653, 32'sd1991026, 32'sd0, 32'sd0, -32'sd82848, 32'sd632484, -32'sd1136303, 32'sd621499, -32'sd393399, -32'sd2020075, -32'sd947532, -32'sd1478290, -32'sd1415205, -32'sd3355196, -32'sd2771601, -32'sd487353, -32'sd1159400, -32'sd104503, 32'sd1188540, 32'sd1256647, -32'sd1143109, 32'sd748937, 32'sd775843, -32'sd1077041, -32'sd1275994, -32'sd1279524, -32'sd710611, -32'sd243280, -32'sd128937, -32'sd951798, 32'sd83577, 32'sd0, 32'sd527550, -32'sd390797, -32'sd796901, 32'sd650108, -32'sd2485077, -32'sd1451232, -32'sd2651474, -32'sd1186169, -32'sd36662, -32'sd1273994, -32'sd1042690, -32'sd2622892, 32'sd1138454, 32'sd1681833, -32'sd267037, 32'sd14762, -32'sd631192, 32'sd737099, 32'sd21769, -32'sd2527937, -32'sd67167, 32'sd128394, -32'sd721012, 32'sd18808, -32'sd74688, 32'sd662112, 32'sd627123, 32'sd0, 32'sd454607, 32'sd786259, -32'sd1555287, -32'sd222584, 32'sd1088804, 32'sd735194, -32'sd1418591, -32'sd2808186, -32'sd955390, 32'sd223541, -32'sd2735313, -32'sd2859494, -32'sd417140, -32'sd1669995, -32'sd1246114, -32'sd750346, 32'sd1825094, 32'sd137722, 32'sd1401062, 32'sd939773, 32'sd730427, 32'sd1181619, -32'sd212838, 32'sd849956, -32'sd1898488, 32'sd240877, 32'sd509420, 32'sd1169688, -32'sd228989, -32'sd408766, -32'sd1081493, -32'sd1025100, 32'sd1058358, 32'sd1056229, -32'sd170259, -32'sd2197648, -32'sd981656, -32'sd1261570, -32'sd1914235, -32'sd1024605, -32'sd69503, 32'sd343399, 32'sd654470, 32'sd1122833, 32'sd687978, 32'sd2573303, 32'sd378209, 32'sd2279608, -32'sd663713, 32'sd293946, 32'sd996501, 32'sd96693, -32'sd2149269, 32'sd1375976, -32'sd1111298, 32'sd773134, 32'sd1165447, 32'sd219494, 32'sd331826, 32'sd205554, 32'sd566633, 32'sd450868, -32'sd863583, -32'sd2843960, -32'sd1971721, -32'sd1542808, 32'sd798264, 32'sd355833, -32'sd993621, 32'sd1751754, 32'sd907885, 32'sd2196593, 32'sd1962277, 32'sd2402886, 32'sd3101205, 32'sd3410091, 32'sd1913130, 32'sd3057596, 32'sd2425505, -32'sd1764925, 32'sd28785, 32'sd375319, 32'sd1414658, -32'sd245824, -32'sd1561322, 32'sd442694, 32'sd300336, -32'sd938751, -32'sd884864, 32'sd208043, 32'sd362398, -32'sd726957, -32'sd131700, -32'sd1300788, -32'sd614609, 32'sd3380342, 32'sd253016, 32'sd797674, 32'sd2139587, 32'sd635825, 32'sd1608884, 32'sd2208662, 32'sd481953, 32'sd2694290, 32'sd2750809, 32'sd1238432, 32'sd1746596, 32'sd115470, 32'sd746643, -32'sd877538, -32'sd113295, 32'sd310378, -32'sd1322611, -32'sd129008, -32'sd2147961, 32'sd242225, -32'sd1109764, -32'sd1398389, -32'sd1286130, -32'sd351059, -32'sd501987, 32'sd1134533, -32'sd503529, 32'sd738631, 32'sd1442329, 32'sd2125871, 32'sd630633, 32'sd2484049, 32'sd54358, 32'sd1318575, -32'sd518564, 32'sd731249, 32'sd1522907, 32'sd1340619, 32'sd620124, 32'sd862628, 32'sd411780, 32'sd1505904, 32'sd833850, 32'sd1044536, 32'sd1953595, -32'sd473577, -32'sd1139364, -32'sd1523553, -32'sd2045976, -32'sd5482, 32'sd132774, -32'sd521947, 32'sd342592, 32'sd443742, 32'sd789054, -32'sd1954577, -32'sd83259, 32'sd464065, 32'sd1676243, -32'sd432719, -32'sd1473189, -32'sd964175, 32'sd1060366, 32'sd1295722, -32'sd1044981, -32'sd856895, 32'sd30397, 32'sd2205334, -32'sd227158, -32'sd215670, 32'sd978565, 32'sd1286023, -32'sd525686, 32'sd305523, 32'sd1272615, -32'sd2341201, -32'sd1966395, 32'sd131095, -32'sd1102230, -32'sd1765388, -32'sd250166, 32'sd242691, -32'sd444371, -32'sd1790700, 32'sd351152, 32'sd1118118, 32'sd247712, 32'sd876820, -32'sd553860, 32'sd2021086, -32'sd171443, -32'sd1290083, 32'sd328601, 32'sd1781153, 32'sd1448170, -32'sd40196, 32'sd497132, -32'sd913649, 32'sd1427365, 32'sd399597, 32'sd1538454, 32'sd747113, 32'sd1262867, -32'sd1093951, -32'sd1556421, 32'sd1122646, 32'sd304939, -32'sd98126, -32'sd228657, 32'sd1600630, 32'sd438153, 32'sd998609, 32'sd1515064, 32'sd1393312, -32'sd382043, -32'sd1321073, -32'sd303136, -32'sd1823285, -32'sd1677917, -32'sd744593, 32'sd593888, 32'sd1250768, 32'sd664511, 32'sd153, -32'sd481392, -32'sd1059693, 32'sd1636579, 32'sd476909, 32'sd755317, -32'sd90708, 32'sd604734, -32'sd735385, 32'sd2922077, 32'sd413353, -32'sd1447601, -32'sd770422, 32'sd938533, 32'sd1402593, 32'sd2424245, 32'sd366324, 32'sd1049153, -32'sd966005, -32'sd980418, -32'sd2630758, 32'sd535094, -32'sd1099808, -32'sd1205775, 32'sd71085, 32'sd717388, -32'sd1001630, 32'sd963450, 32'sd1206921, -32'sd1622393, -32'sd1233019, -32'sd222867, -32'sd289190, 32'sd184905, -32'sd1774367, -32'sd2451980, 32'sd629773, 32'sd3567123, 32'sd1782014, -32'sd339619, 32'sd103933, -32'sd344063, 32'sd1723840, 32'sd1672003, 32'sd172848, -32'sd2381071, -32'sd3893131, -32'sd128383, -32'sd1483630, -32'sd528308, 32'sd1457258, -32'sd166806, -32'sd637132, -32'sd587979, 32'sd723181, -32'sd8130, 32'sd2941557, 32'sd220674, -32'sd448014, -32'sd301246, 32'sd402203, 32'sd733586, 32'sd82960, -32'sd1536527, -32'sd94993, 32'sd1686569, 32'sd479442, -32'sd1372655, -32'sd499320, -32'sd538187, 32'sd895298, 32'sd1497365, -32'sd852124, -32'sd4663381, -32'sd2574452, -32'sd379885, 32'sd370698, -32'sd150947, 32'sd308213, -32'sd905836, 32'sd466544, -32'sd542241, 32'sd825889, -32'sd1354396, -32'sd375570, 32'sd1734884, 32'sd1580474, 32'sd816368, 32'sd0, -32'sd611659, -32'sd573447, -32'sd4420, -32'sd10191, -32'sd97135, 32'sd1295027, 32'sd1782857, -32'sd122416, 32'sd1682116, 32'sd823304, -32'sd1268034, -32'sd844589, -32'sd1995487, -32'sd1517760, -32'sd995784, 32'sd1682545, -32'sd28868, -32'sd291983, 32'sd519409, 32'sd121528, -32'sd1279969, -32'sd2066158, 32'sd558950, 32'sd450117, 32'sd118134, -32'sd153948, 32'sd804129, -32'sd768890, 32'sd591235, -32'sd503829, -32'sd2286422, 32'sd773495, 32'sd491355, 32'sd619538, -32'sd661719, 32'sd1678468, 32'sd2412263, 32'sd1276943, -32'sd1836261, -32'sd3129171, -32'sd3124524, -32'sd461212, 32'sd1760522, -32'sd316356, 32'sd51137, -32'sd2024384, -32'sd1976430, 32'sd522889, -32'sd1543176, -32'sd241167, -32'sd1362373, 32'sd1049977, -32'sd593218, -32'sd672958, 32'sd792445, 32'sd1595988, 32'sd999145, 32'sd246504, -32'sd2442928, -32'sd1489067, 32'sd1171268, 32'sd230408, 32'sd1630113, 32'sd2691341, 32'sd267272, 32'sd1996747, -32'sd654087, 32'sd90262, -32'sd1491995, -32'sd706717, -32'sd838796, -32'sd1264910, -32'sd869896, -32'sd1516794, -32'sd1919417, 32'sd244148, 32'sd510672, 32'sd559160, 32'sd499599, 32'sd502869, 32'sd1062705, 32'sd572556, -32'sd886554, 32'sd0, 32'sd1318610, -32'sd961828, -32'sd725711, -32'sd680636, 32'sd867964, -32'sd1792610, -32'sd1357653, 32'sd3867, -32'sd96026, 32'sd1271296, 32'sd103402, 32'sd695162, -32'sd646056, -32'sd1698533, -32'sd255841, -32'sd1069908, 32'sd685297, -32'sd360056, 32'sd66250, -32'sd167579, 32'sd1580176, -32'sd88182, 32'sd160540, -32'sd1090132, -32'sd745170, -32'sd939882, 32'sd2010077, 32'sd503685, -32'sd1762564, -32'sd168243, -32'sd818171, 32'sd788694, -32'sd279850, 32'sd390562, -32'sd874547, 32'sd501680, -32'sd119144, 32'sd1280869, 32'sd869187, -32'sd1029157, -32'sd996365, 32'sd10306, -32'sd89924, -32'sd32004, -32'sd1963395, -32'sd642262, -32'sd1271372, -32'sd1558738, -32'sd893279, -32'sd382323, 32'sd648642, -32'sd3190938, -32'sd2948569, -32'sd916562, 32'sd320541, -32'sd556081, -32'sd1008401, -32'sd1370946, 32'sd712121, -32'sd1967799, -32'sd1335729, 32'sd2719979, 32'sd1015502, 32'sd941078, -32'sd370734, -32'sd432929, -32'sd77559, 32'sd752448, 32'sd522327, 32'sd1119884, 32'sd1079741, -32'sd714058, -32'sd1179057, 32'sd1337676, 32'sd25177, -32'sd667095, -32'sd898871, -32'sd2021787, -32'sd203453, -32'sd1301411, -32'sd1272378, -32'sd831688, 32'sd1108159, 32'sd0, -32'sd67944, -32'sd979491, -32'sd1182583, -32'sd819149, -32'sd1666836, -32'sd468434, 32'sd1148926, -32'sd1297629, 32'sd1529080, 32'sd1263335, 32'sd1613286, 32'sd2326066, 32'sd1878486, 32'sd1433652, 32'sd1987512, -32'sd723591, 32'sd1712145, -32'sd577663, 32'sd105163, -32'sd1673893, -32'sd1450021, -32'sd1022082, 32'sd508757, 32'sd1493606, -32'sd151918, -32'sd626920, 32'sd0, 32'sd0, 32'sd0, 32'sd109336, 32'sd195546, -32'sd2475749, -32'sd1706688, 32'sd857065, -32'sd240417, 32'sd1751740, 32'sd49564, 32'sd1205352, 32'sd2481025, 32'sd5683420, 32'sd1254617, 32'sd1797874, 32'sd1307520, -32'sd1405180, 32'sd1571132, -32'sd1115078, 32'sd626141, 32'sd1448094, 32'sd390917, -32'sd330115, 32'sd415758, 32'sd182685, -32'sd1116354, 32'sd973395, 32'sd0, 32'sd0, 32'sd0, 32'sd823361, 32'sd1013580, 32'sd763081, -32'sd1686649, 32'sd1373777, -32'sd1281967, -32'sd1494039, 32'sd1237723, 32'sd393238, 32'sd330857, 32'sd80770, -32'sd1214319, -32'sd793577, -32'sd1010023, -32'sd667453, 32'sd637431, 32'sd1224786, 32'sd446086, 32'sd755139, -32'sd722757, -32'sd434144, -32'sd1133207, 32'sd183132, 32'sd75553, 32'sd414721, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd661356, -32'sd1810226, 32'sd808588, -32'sd327959, 32'sd154046, -32'sd1196075, -32'sd1834511, -32'sd158661, -32'sd961653, -32'sd499094, -32'sd1170381, 32'sd133673, -32'sd512309, -32'sd745056, -32'sd2083, -32'sd598512, 32'sd439039, 32'sd349234, 32'sd1084936, 32'sd1502525, 32'sd1253168, -32'sd1581278, -32'sd253242, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd612207, 32'sd1337368, 32'sd116710, 32'sd240869, -32'sd903974, -32'sd346201, 32'sd1315515, 32'sd288718, 32'sd272858, 32'sd2139941, 32'sd1514370, 32'sd430811, -32'sd1334887, -32'sd270079, -32'sd428864, 32'sd943440, 32'sd1938689, 32'sd1801722, -32'sd259056, 32'sd517390, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1207884, 32'sd984904, -32'sd691282, -32'sd141319, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd855732, 32'sd564472, -32'sd275863, 32'sd407952, 32'sd1331072, 32'sd402372, 32'sd132749, -32'sd1079485, 32'sd492966, 32'sd1406919, 32'sd584429, 32'sd14851, -32'sd310202, 32'sd1193399, 32'sd1894827, 32'sd1221256, 32'sd954347, 32'sd1082488, 32'sd1009631, 32'sd758663, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1875057, 32'sd1264730, 32'sd1407176, -32'sd189651, 32'sd452662, 32'sd698915, 32'sd1173761, 32'sd2030203, 32'sd981392, 32'sd354032, 32'sd2180428, 32'sd654738, 32'sd540679, 32'sd61692, -32'sd981813, -32'sd439292, -32'sd1297196, 32'sd1773903, 32'sd2425677, 32'sd79878, 32'sd17210, 32'sd1721419, 32'sd1588456, 32'sd1514112, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd534953, -32'sd422986, -32'sd270646, 32'sd1808621, 32'sd898177, 32'sd881867, 32'sd727633, -32'sd208787, -32'sd696003, -32'sd1129767, 32'sd867358, 32'sd554200, 32'sd652053, -32'sd1298890, 32'sd184632, -32'sd1907249, -32'sd2437842, -32'sd2321304, 32'sd714018, -32'sd327432, -32'sd453315, -32'sd55479, 32'sd1596018, 32'sd205193, -32'sd838099, 32'sd0, 32'sd0, 32'sd701010, 32'sd449995, -32'sd100619, -32'sd1301993, -32'sd960896, 32'sd301959, 32'sd443509, -32'sd620551, 32'sd194406, -32'sd766708, 32'sd1234871, 32'sd548987, -32'sd574443, -32'sd897400, -32'sd473694, -32'sd1793424, -32'sd1542652, 32'sd889506, -32'sd34233, 32'sd1109091, 32'sd1866240, -32'sd111685, 32'sd718558, -32'sd49026, -32'sd1681354, -32'sd173922, 32'sd1862074, 32'sd0, 32'sd969592, -32'sd242081, 32'sd216766, 32'sd370365, 32'sd1244507, -32'sd603730, -32'sd639081, 32'sd1514007, -32'sd1223323, -32'sd1928728, -32'sd2179333, -32'sd2126048, -32'sd3000909, -32'sd604457, -32'sd2729387, -32'sd2432807, 32'sd906283, -32'sd1163090, 32'sd1547329, 32'sd1019780, 32'sd1141373, -32'sd1755831, -32'sd727844, -32'sd1075657, -32'sd244542, -32'sd486913, -32'sd298172, 32'sd0, 32'sd846555, 32'sd993455, -32'sd86111, 32'sd1663791, 32'sd406889, 32'sd614251, -32'sd467502, 32'sd931534, -32'sd1546392, -32'sd695026, -32'sd1877303, -32'sd593806, -32'sd272501, -32'sd461639, -32'sd925224, 32'sd248388, -32'sd992187, 32'sd321359, -32'sd40148, -32'sd344449, 32'sd1420810, 32'sd1211808, -32'sd82420, -32'sd1136636, 32'sd376895, -32'sd349357, 32'sd1514477, 32'sd2006226, 32'sd386355, 32'sd860456, 32'sd736914, 32'sd113732, -32'sd234442, 32'sd1056657, 32'sd417732, -32'sd904847, -32'sd2566549, -32'sd1847742, -32'sd1226777, 32'sd196224, 32'sd1147941, -32'sd1011429, -32'sd1999179, 32'sd1219310, 32'sd1196823, 32'sd1550503, 32'sd891223, -32'sd976185, 32'sd988840, 32'sd55788, -32'sd1077228, 32'sd1255182, 32'sd1174764, 32'sd680922, 32'sd319387, 32'sd1198289, 32'sd413578, 32'sd731461, -32'sd167578, 32'sd124405, -32'sd1777665, 32'sd844385, 32'sd113951, -32'sd515208, -32'sd1259677, 32'sd1261114, -32'sd518072, 32'sd479451, -32'sd2071357, -32'sd528571, 32'sd261543, 32'sd35140, 32'sd2105697, 32'sd641830, -32'sd1328833, 32'sd1761252, -32'sd1004315, 32'sd64272, -32'sd783779, 32'sd396794, -32'sd215628, -32'sd1540815, 32'sd878320, 32'sd1269529, 32'sd1795236, 32'sd1096974, 32'sd201614, 32'sd1351447, -32'sd1474796, 32'sd53683, -32'sd1327858, -32'sd479828, 32'sd1366952, 32'sd2296756, 32'sd1346597, 32'sd144053, -32'sd119755, -32'sd77164, -32'sd549410, 32'sd137812, 32'sd358755, 32'sd213213, 32'sd1927616, 32'sd308117, 32'sd1478005, 32'sd691548, 32'sd348236, 32'sd149264, 32'sd480792, -32'sd1272550, 32'sd673146, 32'sd1544338, -32'sd270607, 32'sd2972943, 32'sd39268, 32'sd1248823, 32'sd454673, 32'sd528190, 32'sd1425295, -32'sd16507, 32'sd596770, 32'sd1641380, 32'sd1723583, 32'sd690657, 32'sd2256302, 32'sd997537, 32'sd491093, 32'sd1833368, -32'sd463545, 32'sd2333446, 32'sd208726, 32'sd1046920, 32'sd2476598, 32'sd1687673, -32'sd1388356, 32'sd1604926, 32'sd663162, 32'sd424409, 32'sd1588153, 32'sd141365, 32'sd1225061, 32'sd872902, 32'sd1388049, 32'sd928908, 32'sd770929, 32'sd773247, 32'sd2091886, 32'sd862847, 32'sd422261, 32'sd50004, 32'sd3700006, 32'sd394188, 32'sd2476954, 32'sd4009500, 32'sd3335784, 32'sd837668, -32'sd467294, 32'sd883064, 32'sd1866808, 32'sd2406905, 32'sd1867887, 32'sd2847994, 32'sd1202363, 32'sd1488228, -32'sd389075, -32'sd575384, 32'sd313467, 32'sd748602, 32'sd822502, -32'sd66966, 32'sd1687440, 32'sd1991799, 32'sd3069163, 32'sd1238011, 32'sd1547464, 32'sd1569073, 32'sd2427544, 32'sd2689402, 32'sd4493350, 32'sd2923615, 32'sd1421618, 32'sd264961, 32'sd1242684, 32'sd7191, -32'sd952016, -32'sd22323, -32'sd292757, 32'sd1889818, 32'sd2911096, 32'sd1491922, 32'sd1642829, 32'sd490097, -32'sd494705, 32'sd66817, -32'sd397085, 32'sd884293, -32'sd1129105, 32'sd1001041, -32'sd346984, 32'sd1740219, 32'sd3810917, 32'sd1854099, 32'sd1814054, 32'sd693580, 32'sd505020, 32'sd2413299, 32'sd1056541, 32'sd11799, -32'sd1236959, -32'sd2676754, -32'sd2974922, -32'sd2207384, -32'sd4311368, -32'sd1012303, -32'sd963942, -32'sd597501, 32'sd1685094, 32'sd2653509, 32'sd2662825, -32'sd544234, 32'sd1012051, 32'sd1346290, 32'sd421992, 32'sd759323, -32'sd922490, -32'sd326872, 32'sd1615840, 32'sd2240563, 32'sd547791, 32'sd1775911, 32'sd618926, 32'sd2760706, -32'sd20416, -32'sd445363, -32'sd1457030, -32'sd2446895, -32'sd2889111, -32'sd3053138, -32'sd346503, -32'sd3249608, -32'sd3320793, -32'sd884127, -32'sd1713006, 32'sd1198698, 32'sd2029171, 32'sd2794766, 32'sd1449325, -32'sd2490824, -32'sd2776608, -32'sd160997, 32'sd812650, 32'sd454554, 32'sd614439, -32'sd284445, 32'sd800163, 32'sd825302, -32'sd341514, 32'sd1661599, 32'sd268676, 32'sd572610, -32'sd1310849, -32'sd430971, -32'sd1607623, -32'sd2182273, -32'sd510871, -32'sd140435, -32'sd1004636, -32'sd2482954, -32'sd2289089, -32'sd2125706, -32'sd2088723, 32'sd490467, 32'sd1692099, 32'sd1518682, -32'sd628857, -32'sd600909, 32'sd510536, -32'sd861373, 32'sd930888, 32'sd759815, -32'sd922134, -32'sd391464, -32'sd1061093, -32'sd435883, 32'sd1357896, -32'sd547623, 32'sd1035250, -32'sd66249, -32'sd1336495, -32'sd809223, -32'sd3013960, -32'sd3261614, -32'sd2704423, -32'sd1273143, -32'sd1181722, -32'sd1719755, -32'sd1842539, -32'sd1112497, -32'sd1030073, 32'sd829039, 32'sd461573, 32'sd1287646, 32'sd1597459, -32'sd217511, -32'sd1206463, -32'sd154741, -32'sd278669, 32'sd0, 32'sd695703, -32'sd372837, 32'sd125098, 32'sd949255, 32'sd1166200, 32'sd16330, 32'sd1472443, 32'sd213944, 32'sd171208, -32'sd2203406, -32'sd3069847, -32'sd1561368, 32'sd150867, -32'sd1446682, -32'sd1265673, -32'sd3147607, -32'sd14457, -32'sd829608, 32'sd1293103, 32'sd82595, 32'sd648569, 32'sd2065267, 32'sd332845, -32'sd1297502, 32'sd917622, 32'sd19416, 32'sd313175, 32'sd672514, 32'sd93732, -32'sd1355217, -32'sd60219, -32'sd679596, -32'sd1454051, -32'sd507785, 32'sd1050743, 32'sd2030090, 32'sd1129855, -32'sd178423, -32'sd1630783, -32'sd1757042, 32'sd519613, -32'sd448941, -32'sd263323, -32'sd1623849, 32'sd1348450, 32'sd1307357, -32'sd811484, -32'sd253049, 32'sd555962, 32'sd1491386, -32'sd492869, -32'sd480986, -32'sd110019, 32'sd406083, 32'sd224769, 32'sd867819, 32'sd626414, 32'sd258317, 32'sd1311848, 32'sd445670, 32'sd554249, -32'sd1178861, 32'sd1508757, 32'sd1150769, 32'sd950377, 32'sd1391954, -32'sd1020048, 32'sd1606230, -32'sd874153, -32'sd846373, 32'sd636454, 32'sd601552, 32'sd1727701, 32'sd431336, -32'sd1413357, 32'sd909944, -32'sd2319645, -32'sd695255, -32'sd492063, 32'sd379838, 32'sd759528, -32'sd1763067, 32'sd522401, 32'sd0, 32'sd964831, -32'sd1595560, -32'sd240704, -32'sd156319, -32'sd1218352, -32'sd588278, 32'sd1548945, 32'sd2847921, 32'sd1626885, 32'sd2298754, -32'sd1179518, -32'sd284743, 32'sd1408670, 32'sd114642, -32'sd1722711, 32'sd283203, -32'sd365794, 32'sd151812, -32'sd3018955, -32'sd2100373, 32'sd22192, 32'sd215639, -32'sd1346305, -32'sd752957, 32'sd2032990, -32'sd308739, 32'sd1082657, -32'sd594515, 32'sd64445, 32'sd371322, 32'sd1407759, -32'sd1040714, -32'sd1489578, 32'sd123075, 32'sd2868001, 32'sd1985023, -32'sd102825, -32'sd64442, -32'sd375890, 32'sd1115888, -32'sd1339292, -32'sd2012307, -32'sd607691, 32'sd498782, -32'sd1893452, -32'sd1249789, -32'sd2627217, -32'sd2119365, 32'sd150430, -32'sd1558476, 32'sd389759, 32'sd718599, 32'sd868238, -32'sd834614, -32'sd51462, 32'sd614969, -32'sd345966, -32'sd2136867, 32'sd1589862, 32'sd696929, 32'sd1174414, 32'sd442791, 32'sd1489115, 32'sd2295842, 32'sd1598088, 32'sd1208788, 32'sd294192, 32'sd143594, 32'sd705690, -32'sd1494662, -32'sd471150, -32'sd1995606, 32'sd1010326, -32'sd871460, -32'sd1692035, -32'sd2314539, -32'sd1397298, 32'sd1591740, 32'sd436411, 32'sd1182106, 32'sd1929200, -32'sd998771, 32'sd1293777, 32'sd0, 32'sd805361, 32'sd216960, -32'sd1687779, -32'sd1090742, -32'sd627684, -32'sd90169, -32'sd555546, 32'sd792023, -32'sd887546, 32'sd894055, -32'sd25862, -32'sd790850, 32'sd455135, -32'sd59889, 32'sd208885, 32'sd1711755, 32'sd198469, -32'sd104579, -32'sd1513493, -32'sd848783, -32'sd1802950, -32'sd720304, 32'sd682368, -32'sd432283, 32'sd443674, 32'sd231410, 32'sd0, 32'sd0, 32'sd0, -32'sd1246632, 32'sd39368, 32'sd1530128, 32'sd1875870, -32'sd120797, 32'sd83481, 32'sd775440, -32'sd169213, 32'sd2094448, 32'sd50614, 32'sd2176666, 32'sd807783, -32'sd89151, 32'sd226755, 32'sd1391635, 32'sd2207176, -32'sd664236, -32'sd533064, -32'sd111958, -32'sd974316, -32'sd49768, -32'sd609248, -32'sd444420, -32'sd1114084, 32'sd1660201, 32'sd0, 32'sd0, 32'sd0, 32'sd1315348, 32'sd719476, -32'sd694929, -32'sd628275, -32'sd371820, 32'sd67160, -32'sd991196, -32'sd412151, 32'sd522645, -32'sd634560, -32'sd2923318, -32'sd1638103, 32'sd496719, -32'sd492546, 32'sd3192773, -32'sd653206, -32'sd3244662, -32'sd1264210, -32'sd71669, -32'sd746824, 32'sd1148566, 32'sd856652, 32'sd70870, 32'sd1592554, 32'sd754137, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd866441, 32'sd874891, -32'sd427339, -32'sd182522, -32'sd1463557, 32'sd586868, 32'sd386518, -32'sd633062, 32'sd131375, -32'sd411186, 32'sd1920449, 32'sd1009567, 32'sd2175463, 32'sd1339581, -32'sd50163, -32'sd1669419, 32'sd869871, -32'sd753552, -32'sd425291, 32'sd1677649, -32'sd1041473, 32'sd1817003, 32'sd1978475, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd774822, 32'sd1102520, 32'sd458865, 32'sd33616, 32'sd2321601, 32'sd267083, 32'sd2276913, -32'sd305363, 32'sd1062010, 32'sd400208, 32'sd2007810, -32'sd121147, 32'sd2861059, 32'sd1243747, 32'sd665622, -32'sd944932, -32'sd43483, 32'sd1620967, 32'sd2517313, 32'sd981924, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1336679, 32'sd1605476, 32'sd801512, 32'sd316044, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd63405, 32'sd1308046, -32'sd1712435, -32'sd378363, -32'sd641844, -32'sd752557, 32'sd1367651, 32'sd1013442, 32'sd845160, 32'sd1888834, 32'sd213397, -32'sd447859, -32'sd968227, 32'sd786877, -32'sd641775, -32'sd852297, 32'sd861373, 32'sd1123615, -32'sd75293, 32'sd796869, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2087912, 32'sd175019, 32'sd475578, -32'sd1206153, 32'sd584584, 32'sd1092671, -32'sd1502296, -32'sd1484241, 32'sd1976081, 32'sd520620, -32'sd497558, 32'sd734892, 32'sd630198, -32'sd974870, 32'sd368002, -32'sd1058364, -32'sd206285, -32'sd608950, 32'sd784796, 32'sd2447508, 32'sd166110, 32'sd1206253, 32'sd842691, 32'sd1241885, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd576563, -32'sd92489, -32'sd213723, 32'sd1033390, 32'sd613574, 32'sd842953, -32'sd738240, -32'sd2673683, -32'sd1608024, 32'sd37015, -32'sd523449, -32'sd1109165, -32'sd911394, -32'sd1803171, -32'sd4027931, -32'sd1947361, -32'sd1292213, 32'sd1934733, 32'sd672574, -32'sd456135, 32'sd436186, -32'sd557941, 32'sd1286342, 32'sd115045, 32'sd497481, 32'sd0, 32'sd0, 32'sd1253743, 32'sd908676, 32'sd824992, -32'sd302647, -32'sd705146, -32'sd501605, -32'sd1684920, -32'sd12690, -32'sd381924, -32'sd2141995, 32'sd989556, 32'sd157941, -32'sd617623, -32'sd318449, -32'sd1910619, 32'sd1355491, 32'sd1113355, 32'sd925470, 32'sd2203926, 32'sd1977315, 32'sd1103640, 32'sd389113, 32'sd235305, 32'sd593491, -32'sd1259102, 32'sd2275387, 32'sd490221, 32'sd0, 32'sd1349673, -32'sd158502, 32'sd792307, -32'sd1016558, 32'sd865218, 32'sd708520, -32'sd655827, -32'sd214473, 32'sd1588208, -32'sd85512, -32'sd2068170, -32'sd2389877, -32'sd1515056, -32'sd3144026, -32'sd2474204, 32'sd64478, -32'sd588567, 32'sd2525177, 32'sd2000989, 32'sd2661308, 32'sd895210, 32'sd593100, 32'sd2447467, -32'sd933364, -32'sd1157388, -32'sd302002, 32'sd96704, 32'sd0, 32'sd319312, -32'sd11733, -32'sd1067142, 32'sd1828033, 32'sd208631, 32'sd2690705, 32'sd1966367, 32'sd1145843, 32'sd957491, -32'sd413740, 32'sd8517, -32'sd330175, -32'sd1620285, -32'sd3357311, -32'sd4444290, -32'sd1224723, 32'sd1539792, 32'sd1811867, 32'sd2366410, 32'sd1321517, 32'sd2529484, -32'sd672403, -32'sd647140, -32'sd1246806, -32'sd1888773, 32'sd51114, 32'sd691345, 32'sd2123636, 32'sd451941, 32'sd579177, 32'sd437104, 32'sd549056, -32'sd664517, 32'sd867556, 32'sd1395747, -32'sd1362548, 32'sd1839915, 32'sd514193, -32'sd1612279, -32'sd606915, -32'sd1672155, -32'sd3310607, -32'sd3259852, 32'sd1171511, 32'sd4505700, 32'sd3868566, 32'sd3492695, 32'sd879876, 32'sd1698887, 32'sd1708036, 32'sd958099, -32'sd44166, -32'sd1810719, -32'sd880860, 32'sd208354, 32'sd935080, 32'sd956951, -32'sd1407626, 32'sd708267, -32'sd1637968, -32'sd1008531, 32'sd459551, 32'sd737930, -32'sd1347195, 32'sd570792, 32'sd241624, -32'sd1212174, -32'sd1074376, -32'sd4199165, -32'sd5075548, -32'sd3570647, 32'sd1327838, 32'sd2683603, 32'sd4026384, 32'sd3129114, 32'sd764192, -32'sd809334, 32'sd887758, 32'sd1034902, -32'sd1435168, 32'sd265869, 32'sd1171940, 32'sd560123, 32'sd1549243, 32'sd603564, -32'sd519816, 32'sd524473, -32'sd715983, -32'sd2389192, -32'sd112195, -32'sd656236, -32'sd24702, -32'sd788161, -32'sd350215, 32'sd1012331, -32'sd188216, -32'sd5571572, -32'sd5197037, 32'sd724055, 32'sd2733995, 32'sd4423073, 32'sd2278129, 32'sd1390576, -32'sd829834, -32'sd481900, 32'sd1388366, -32'sd235402, -32'sd155547, 32'sd65713, -32'sd306339, 32'sd61112, 32'sd1332140, 32'sd170995, -32'sd184472, -32'sd895372, -32'sd1129106, 32'sd554986, 32'sd960556, -32'sd827396, 32'sd99620, 32'sd1606801, 32'sd256625, -32'sd928752, -32'sd2371411, -32'sd5051336, -32'sd3281570, 32'sd3033138, 32'sd3365016, 32'sd3398922, 32'sd940378, -32'sd628537, -32'sd1625651, -32'sd1930907, -32'sd306336, -32'sd160237, 32'sd279854, 32'sd1496673, -32'sd1582846, -32'sd685855, 32'sd1634534, 32'sd656746, -32'sd683557, -32'sd305843, -32'sd852748, -32'sd1109367, 32'sd677433, 32'sd90075, -32'sd1254330, 32'sd229588, 32'sd880570, -32'sd1410309, -32'sd2522518, -32'sd651395, 32'sd116514, 32'sd2444600, 32'sd2468883, 32'sd3282316, 32'sd2534460, 32'sd270532, -32'sd265254, -32'sd448663, 32'sd67442, -32'sd1596124, -32'sd453103, -32'sd662455, 32'sd44151, 32'sd1017769, -32'sd341036, 32'sd71434, 32'sd429423, -32'sd2060879, -32'sd482118, 32'sd1069179, -32'sd1740029, -32'sd1275975, 32'sd629831, 32'sd2245896, -32'sd712712, -32'sd2896421, -32'sd1638693, -32'sd1255628, 32'sd81300, 32'sd1678926, 32'sd989516, 32'sd680570, 32'sd1305124, -32'sd1040141, -32'sd2621288, -32'sd2179390, -32'sd974579, 32'sd208591, 32'sd1394471, 32'sd1178047, 32'sd230282, 32'sd964889, 32'sd655719, 32'sd391132, 32'sd181393, -32'sd280998, 32'sd454133, 32'sd489360, 32'sd1224318, 32'sd94753, 32'sd272287, 32'sd1079195, -32'sd1462783, -32'sd2026659, -32'sd1538777, -32'sd1530924, 32'sd847931, 32'sd859519, 32'sd1042853, 32'sd1418894, 32'sd155402, -32'sd28460, 32'sd119624, 32'sd449366, 32'sd862989, -32'sd1053793, 32'sd224672, 32'sd819608, 32'sd438233, -32'sd1204458, 32'sd1153497, 32'sd61361, 32'sd239323, 32'sd8398, 32'sd523126, 32'sd1046008, 32'sd399474, 32'sd447930, -32'sd979875, 32'sd274598, -32'sd433469, 32'sd949101, -32'sd1895197, 32'sd966088, 32'sd2465737, 32'sd477662, 32'sd1448447, 32'sd1490066, 32'sd1678037, 32'sd1529226, -32'sd243739, 32'sd903061, -32'sd903478, 32'sd446385, -32'sd530414, 32'sd721968, -32'sd43792, 32'sd319844, -32'sd1490181, -32'sd647468, 32'sd265523, 32'sd728569, -32'sd912777, -32'sd756591, -32'sd1429436, -32'sd392724, -32'sd1468573, -32'sd1748207, -32'sd1126703, 32'sd2417979, -32'sd1669902, 32'sd1207684, 32'sd983499, 32'sd218163, 32'sd257986, 32'sd210338, -32'sd98300, 32'sd1605310, -32'sd565073, -32'sd863214, -32'sd287243, 32'sd914793, -32'sd1136538, 32'sd354854, 32'sd679725, 32'sd1305644, 32'sd616377, 32'sd1360102, -32'sd220765, -32'sd123925, 32'sd556578, -32'sd793777, 32'sd382404, 32'sd376687, 32'sd319447, -32'sd868123, 32'sd1275680, -32'sd500582, 32'sd1798347, 32'sd1453184, 32'sd368356, -32'sd52705, 32'sd626140, 32'sd844040, 32'sd883882, 32'sd491657, 32'sd873270, 32'sd78031, -32'sd1101315, 32'sd206104, 32'sd1845838, -32'sd58939, 32'sd204472, 32'sd385570, 32'sd0, 32'sd366843, -32'sd2174324, -32'sd1025263, 32'sd212046, -32'sd573088, -32'sd451335, 32'sd995751, -32'sd447772, -32'sd840105, -32'sd1048817, 32'sd876795, 32'sd577665, 32'sd2850165, 32'sd2248204, -32'sd642977, 32'sd2280, 32'sd835236, 32'sd1834776, 32'sd2647957, 32'sd1678761, 32'sd1417495, 32'sd513323, -32'sd475915, 32'sd848362, 32'sd279570, 32'sd46656, 32'sd108254, -32'sd64192, 32'sd819394, 32'sd396416, -32'sd1551597, -32'sd57208, -32'sd1021327, -32'sd880955, -32'sd1142207, 32'sd140470, 32'sd1265651, -32'sd972841, -32'sd340414, -32'sd1172297, 32'sd2161326, 32'sd429176, -32'sd1457776, -32'sd160647, 32'sd1366481, 32'sd192359, -32'sd1321531, 32'sd66097, -32'sd1784715, -32'sd269095, -32'sd1024371, -32'sd2542883, -32'sd161835, 32'sd312359, 32'sd138735, 32'sd1524902, -32'sd1206738, 32'sd1396463, 32'sd765690, -32'sd1854194, -32'sd1693070, -32'sd572594, 32'sd1244788, -32'sd1796268, 32'sd1459486, -32'sd594815, 32'sd73960, -32'sd219528, -32'sd1127249, 32'sd104707, -32'sd535167, -32'sd249069, -32'sd877189, -32'sd383964, 32'sd417672, -32'sd584205, -32'sd345944, -32'sd989840, -32'sd1244464, 32'sd131108, 32'sd715390, 32'sd44319, 32'sd555209, 32'sd0, -32'sd182629, -32'sd255848, 32'sd2954442, 32'sd1168639, -32'sd1106661, -32'sd851894, -32'sd641549, 32'sd272438, -32'sd952098, -32'sd1578978, -32'sd642298, -32'sd451434, -32'sd804134, -32'sd681550, -32'sd588145, -32'sd1072176, -32'sd62062, 32'sd571051, -32'sd2112435, 32'sd868350, 32'sd2195029, 32'sd66156, 32'sd2393511, -32'sd611938, -32'sd931484, -32'sd241907, 32'sd836801, 32'sd266864, -32'sd6894, 32'sd325705, 32'sd793373, -32'sd273157, -32'sd177331, 32'sd1071853, -32'sd1448136, 32'sd236424, -32'sd1003783, -32'sd163038, 32'sd463235, 32'sd11994, -32'sd184175, -32'sd434407, -32'sd2162930, 32'sd571667, 32'sd637631, -32'sd1267898, -32'sd1453070, 32'sd806721, 32'sd1498274, 32'sd1326856, 32'sd1383101, 32'sd363478, -32'sd834074, 32'sd338768, 32'sd312172, 32'sd1049897, 32'sd1084894, -32'sd105310, 32'sd38244, -32'sd985699, 32'sd1912467, 32'sd1580556, -32'sd304925, -32'sd682330, -32'sd722007, 32'sd1404749, 32'sd283231, 32'sd914926, 32'sd3669247, 32'sd1724932, -32'sd985004, 32'sd68095, 32'sd1248407, 32'sd840811, -32'sd546734, 32'sd10064, 32'sd283298, -32'sd497982, -32'sd1990819, 32'sd529319, -32'sd1178960, 32'sd743446, 32'sd1519525, 32'sd0, 32'sd1805945, -32'sd711259, -32'sd1155983, 32'sd165078, 32'sd314871, 32'sd70214, 32'sd2172014, -32'sd131072, 32'sd1484678, 32'sd698851, -32'sd125044, 32'sd1401551, 32'sd2485055, 32'sd531866, 32'sd207657, 32'sd1124810, 32'sd557756, -32'sd1076514, -32'sd1288501, -32'sd260374, -32'sd581706, 32'sd271007, 32'sd883109, 32'sd242149, 32'sd893354, 32'sd1137914, 32'sd0, 32'sd0, 32'sd0, 32'sd843927, 32'sd1481100, -32'sd758603, 32'sd584054, -32'sd311227, 32'sd478181, -32'sd1013716, -32'sd269282, 32'sd649613, -32'sd997382, 32'sd975345, 32'sd1232837, -32'sd37739, -32'sd1185040, -32'sd602581, -32'sd781502, -32'sd403409, 32'sd871396, 32'sd2121528, -32'sd651156, 32'sd927135, 32'sd753901, -32'sd630843, 32'sd1326862, 32'sd442906, 32'sd0, 32'sd0, 32'sd0, 32'sd551268, 32'sd599050, -32'sd740077, 32'sd1268125, -32'sd471873, -32'sd862126, 32'sd81423, -32'sd242223, -32'sd1289629, -32'sd795366, 32'sd1843426, 32'sd2305402, 32'sd837704, -32'sd2634623, -32'sd1923076, -32'sd2084500, 32'sd317453, -32'sd890379, 32'sd2539120, -32'sd657628, 32'sd632458, -32'sd183403, -32'sd655192, -32'sd803861, -32'sd858350, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1586194, 32'sd795425, -32'sd1303681, 32'sd216904, -32'sd7331, 32'sd1105005, 32'sd322515, 32'sd603595, 32'sd351222, 32'sd1120081, -32'sd187347, -32'sd1337960, 32'sd13322, -32'sd785748, 32'sd202586, 32'sd829407, 32'sd1797871, 32'sd1627063, -32'sd845979, 32'sd2521844, 32'sd751517, -32'sd222059, 32'sd1250029, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1588527, 32'sd2488621, 32'sd933281, 32'sd3005973, 32'sd735300, -32'sd791280, -32'sd472655, -32'sd915426, 32'sd1046818, 32'sd1322034, 32'sd1238027, 32'sd636810, 32'sd990035, -32'sd155938, -32'sd1379898, 32'sd97724, -32'sd584881, 32'sd77024, 32'sd533701, 32'sd1451125, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd33852, -32'sd735680, 32'sd740226, -32'sd298626, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd447253, -32'sd1196526, 32'sd23037, -32'sd1981115, 32'sd441595, -32'sd40438, 32'sd144830, -32'sd346389, -32'sd144639, -32'sd873457, -32'sd534181, -32'sd2019710, -32'sd341291, 32'sd25340, 32'sd801384, -32'sd1203955, 32'sd252110, 32'sd939451, 32'sd770065, -32'sd146365, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd474529, 32'sd1236713, -32'sd308, 32'sd949904, -32'sd847116, 32'sd664647, -32'sd492326, -32'sd1495834, 32'sd242410, -32'sd1578819, -32'sd217715, -32'sd1068721, -32'sd477984, -32'sd3137773, -32'sd1967363, 32'sd450533, -32'sd2467604, -32'sd791816, -32'sd387349, 32'sd163805, -32'sd1172474, -32'sd912061, 32'sd106934, 32'sd1603445, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd243706, 32'sd228193, 32'sd40218, -32'sd1623588, 32'sd779618, 32'sd1812389, -32'sd1649696, -32'sd1587653, 32'sd287498, 32'sd1417059, -32'sd2152902, -32'sd1134939, -32'sd233149, -32'sd185489, -32'sd3130330, -32'sd2084938, -32'sd133382, -32'sd32172, -32'sd933102, 32'sd1444486, 32'sd790296, -32'sd541816, -32'sd407996, 32'sd1916173, -32'sd750042, 32'sd0, 32'sd0, -32'sd38530, 32'sd633954, -32'sd1002914, -32'sd2379238, 32'sd421240, 32'sd1793688, 32'sd297965, -32'sd318714, -32'sd1844176, -32'sd3043905, -32'sd982510, -32'sd1776754, -32'sd924554, 32'sd552828, 32'sd1186055, -32'sd1134785, -32'sd1540436, -32'sd2302862, -32'sd3006291, 32'sd784797, -32'sd813615, 32'sd1516494, 32'sd290210, -32'sd1040443, 32'sd1295152, 32'sd1095753, -32'sd582272, 32'sd0, 32'sd433034, 32'sd83646, 32'sd569037, -32'sd3399080, -32'sd3186723, -32'sd136755, 32'sd1026508, 32'sd841526, 32'sd854575, -32'sd380525, 32'sd791938, -32'sd328764, -32'sd1716485, -32'sd2114973, -32'sd53894, -32'sd1943166, -32'sd1175837, -32'sd1884173, -32'sd2297049, -32'sd325784, -32'sd865590, -32'sd421774, 32'sd1289078, 32'sd721339, -32'sd1295640, -32'sd435271, 32'sd372366, 32'sd0, 32'sd250614, -32'sd1479804, 32'sd1079200, -32'sd1256255, -32'sd411692, 32'sd624875, 32'sd1121441, -32'sd840444, 32'sd2502535, 32'sd1396978, 32'sd443069, -32'sd1346407, 32'sd1067100, 32'sd1611231, -32'sd842299, -32'sd379272, -32'sd292479, 32'sd116788, -32'sd166645, 32'sd1339507, 32'sd1670940, 32'sd143909, 32'sd564667, 32'sd1280187, -32'sd1120119, 32'sd421018, -32'sd744598, 32'sd175061, 32'sd1078690, -32'sd617660, 32'sd1887199, -32'sd623614, -32'sd3384, -32'sd873325, -32'sd618999, -32'sd246165, 32'sd572512, -32'sd1708219, -32'sd1345368, 32'sd426444, 32'sd1279648, -32'sd564960, -32'sd137999, -32'sd744193, -32'sd1650784, -32'sd371335, 32'sd45205, -32'sd121385, 32'sd1226018, -32'sd570506, -32'sd321960, -32'sd1776775, -32'sd458758, -32'sd768328, -32'sd190876, -32'sd531387, -32'sd165564, -32'sd540210, 32'sd12532, -32'sd1181792, -32'sd1233746, 32'sd648117, -32'sd1032719, 32'sd401357, -32'sd769834, -32'sd979977, 32'sd67990, -32'sd481294, 32'sd464795, 32'sd38843, -32'sd733367, -32'sd3577235, -32'sd2476069, -32'sd1751895, -32'sd180453, -32'sd1492762, 32'sd1442598, -32'sd872710, 32'sd477330, 32'sd18871, 32'sd433604, -32'sd375961, -32'sd941540, 32'sd546658, 32'sd1919953, 32'sd2187520, 32'sd534549, -32'sd140136, -32'sd98522, 32'sd493506, -32'sd1420394, 32'sd801833, 32'sd239462, -32'sd1229708, 32'sd873326, 32'sd1657916, -32'sd1659307, -32'sd744082, -32'sd2249624, -32'sd418810, 32'sd1392742, 32'sd795832, -32'sd1544628, -32'sd89393, 32'sd1627923, -32'sd1407678, -32'sd377636, -32'sd1074415, -32'sd925124, -32'sd246742, 32'sd660881, 32'sd1329698, 32'sd993944, -32'sd112817, -32'sd114683, -32'sd473776, 32'sd219418, 32'sd196282, -32'sd512681, -32'sd67575, -32'sd2058791, -32'sd1291205, -32'sd1067683, 32'sd1048521, 32'sd385820, -32'sd1408779, 32'sd111553, 32'sd750796, 32'sd589594, 32'sd538403, 32'sd1456110, 32'sd1242390, 32'sd939689, -32'sd234904, -32'sd2897533, -32'sd561166, 32'sd1738553, -32'sd261036, -32'sd908417, 32'sd1289959, -32'sd621468, 32'sd845669, -32'sd1426189, -32'sd850057, -32'sd1977977, -32'sd64730, -32'sd339948, -32'sd371668, -32'sd1725130, -32'sd311785, 32'sd268909, 32'sd581999, -32'sd709271, 32'sd1484882, 32'sd726214, -32'sd147845, 32'sd2246049, 32'sd2029560, 32'sd756569, -32'sd841860, 32'sd854347, -32'sd1006228, -32'sd3745480, -32'sd2723334, -32'sd13116, -32'sd387817, -32'sd5723, 32'sd1162692, 32'sd1087276, 32'sd22258, 32'sd754984, -32'sd1873061, -32'sd1109876, 32'sd1235028, -32'sd939736, 32'sd1135203, -32'sd861322, 32'sd1806784, 32'sd1270668, 32'sd1274981, 32'sd348937, -32'sd199844, 32'sd1037364, 32'sd1117245, 32'sd677199, -32'sd71311, 32'sd1783947, 32'sd1359426, -32'sd325752, -32'sd2191372, -32'sd2449562, -32'sd153545, -32'sd104120, 32'sd47596, -32'sd1081988, 32'sd10798, 32'sd80556, -32'sd1628142, 32'sd620528, -32'sd454764, 32'sd1602292, 32'sd221184, 32'sd416747, -32'sd711781, -32'sd1237876, 32'sd142091, -32'sd1201437, -32'sd1525400, -32'sd475086, 32'sd748486, -32'sd996061, -32'sd253126, 32'sd334902, 32'sd1077607, 32'sd89890, 32'sd1306426, 32'sd667274, -32'sd2699378, -32'sd3578675, 32'sd295157, -32'sd33045, -32'sd2546295, -32'sd269235, -32'sd269173, 32'sd105886, -32'sd1221071, 32'sd1337023, 32'sd834335, 32'sd919320, 32'sd798655, 32'sd2031506, 32'sd581312, 32'sd376797, 32'sd636810, -32'sd838788, -32'sd605914, -32'sd2507671, -32'sd2881940, -32'sd395711, 32'sd298812, 32'sd2084277, 32'sd2773778, 32'sd1068438, -32'sd55658, 32'sd462307, -32'sd142663, -32'sd2256162, -32'sd562590, 32'sd980924, 32'sd1841223, 32'sd281819, -32'sd706917, 32'sd222518, -32'sd722727, -32'sd646617, 32'sd899585, 32'sd763284, 32'sd901548, 32'sd1311153, 32'sd476778, -32'sd727027, -32'sd229498, -32'sd1104921, -32'sd1503225, -32'sd3047445, -32'sd1603587, 32'sd2597182, -32'sd556431, 32'sd3576287, 32'sd1227263, 32'sd2396509, 32'sd409854, -32'sd733196, 32'sd998666, -32'sd852515, -32'sd808447, 32'sd734477, -32'sd380244, 32'sd1156468, 32'sd284429, 32'sd219835, -32'sd1548849, -32'sd1031474, 32'sd476188, 32'sd1016966, 32'sd793724, 32'sd3093866, 32'sd2944916, -32'sd333663, -32'sd78579, -32'sd104760, 32'sd1011297, 32'sd108871, 32'sd711449, -32'sd140887, -32'sd613554, 32'sd922714, 32'sd2423722, 32'sd1143919, 32'sd2621833, -32'sd419275, 32'sd1418728, 32'sd109567, -32'sd2250646, 32'sd955532, -32'sd965545, 32'sd188822, 32'sd0, 32'sd586568, -32'sd95435, 32'sd30676, -32'sd688758, 32'sd521534, 32'sd1438489, 32'sd917861, 32'sd1364144, 32'sd894901, 32'sd1472701, 32'sd1853740, 32'sd435318, 32'sd804118, -32'sd386502, 32'sd601356, 32'sd609937, -32'sd295499, -32'sd614133, 32'sd1096485, -32'sd657274, -32'sd1209068, -32'sd1477159, -32'sd1990754, -32'sd3479525, 32'sd391021, 32'sd92081, -32'sd283294, 32'sd314376, -32'sd363722, -32'sd799403, -32'sd1384461, -32'sd1176258, -32'sd1255300, -32'sd1114480, 32'sd929251, 32'sd2612212, 32'sd2027655, 32'sd2550074, 32'sd3818715, 32'sd1737828, 32'sd1158544, -32'sd832194, 32'sd281901, 32'sd670631, 32'sd1834489, -32'sd2492402, -32'sd707337, -32'sd1233809, -32'sd959046, -32'sd3252518, -32'sd1018174, -32'sd3663237, -32'sd400449, -32'sd328075, -32'sd1095423, 32'sd491748, -32'sd665107, -32'sd884425, -32'sd1117186, -32'sd2382454, -32'sd1452939, -32'sd792231, 32'sd1299192, 32'sd1043253, 32'sd386745, 32'sd2551822, 32'sd3031783, 32'sd2020156, -32'sd1329551, -32'sd74440, -32'sd542322, -32'sd887316, 32'sd400557, -32'sd2397104, -32'sd1907604, -32'sd1003470, -32'sd1226295, -32'sd3173184, -32'sd1432372, -32'sd2144369, 32'sd87027, 32'sd170469, 32'sd1000861, 32'sd0, 32'sd591540, -32'sd1381603, -32'sd821181, 32'sd497092, -32'sd405116, -32'sd938903, -32'sd667652, -32'sd853227, -32'sd2009954, 32'sd113959, -32'sd1029447, -32'sd529091, -32'sd1665391, -32'sd2103180, -32'sd1007093, -32'sd855333, 32'sd152679, -32'sd638604, 32'sd876399, -32'sd1897459, -32'sd2163910, -32'sd1010854, -32'sd882861, -32'sd1502051, 32'sd1217711, -32'sd1844741, 32'sd705683, -32'sd241643, -32'sd690305, -32'sd337009, -32'sd608363, 32'sd32809, -32'sd491575, -32'sd14969, -32'sd5291, -32'sd2573354, -32'sd1154485, -32'sd3236581, -32'sd3593174, -32'sd1621142, -32'sd3745224, -32'sd3740519, -32'sd1800389, -32'sd881589, -32'sd790364, -32'sd131195, 32'sd436453, 32'sd30652, 32'sd412750, 32'sd1375862, 32'sd626356, 32'sd685853, 32'sd1175646, -32'sd828201, 32'sd724573, 32'sd862224, -32'sd57589, 32'sd312428, -32'sd922684, -32'sd700373, -32'sd453121, -32'sd819531, -32'sd1260578, 32'sd68557, -32'sd1773422, -32'sd1616081, -32'sd2443750, -32'sd2947573, -32'sd2982272, -32'sd2155403, -32'sd2917648, 32'sd605099, -32'sd2396921, 32'sd1243345, -32'sd174502, 32'sd1109901, 32'sd709265, 32'sd559330, -32'sd621738, 32'sd276324, 32'sd1712467, -32'sd746385, 32'sd166077, 32'sd0, 32'sd1124047, 32'sd510767, -32'sd1981922, -32'sd167471, -32'sd206068, 32'sd1197100, 32'sd1100893, -32'sd555757, -32'sd2456468, -32'sd2011814, -32'sd1552548, -32'sd2337423, -32'sd1943207, -32'sd570774, -32'sd1888417, -32'sd420643, -32'sd1036906, -32'sd908891, 32'sd507896, -32'sd1302089, 32'sd623388, 32'sd1377829, -32'sd17607, 32'sd119141, 32'sd283936, 32'sd119956, 32'sd0, 32'sd0, 32'sd0, -32'sd871070, -32'sd247386, -32'sd562315, 32'sd1982390, 32'sd29649, 32'sd1452370, -32'sd498774, -32'sd588125, -32'sd1608566, 32'sd523127, -32'sd3393663, -32'sd1199796, -32'sd638174, -32'sd1337343, -32'sd1057691, 32'sd555404, -32'sd914760, 32'sd591116, 32'sd561038, 32'sd1510585, -32'sd591352, 32'sd970268, -32'sd656641, -32'sd313073, 32'sd653330, 32'sd0, 32'sd0, 32'sd0, 32'sd638367, -32'sd297145, 32'sd1232444, 32'sd2204726, -32'sd739786, 32'sd663544, -32'sd488537, -32'sd2918148, 32'sd23800, 32'sd1731678, -32'sd1156882, -32'sd1107098, 32'sd199109, -32'sd3219558, -32'sd335390, 32'sd965111, 32'sd872501, -32'sd312834, -32'sd984082, -32'sd296410, 32'sd1514074, 32'sd1132094, 32'sd669488, 32'sd422963, -32'sd1167064, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1132526, 32'sd1206771, 32'sd1171934, 32'sd806456, 32'sd117149, -32'sd694132, 32'sd550592, -32'sd463119, -32'sd358886, -32'sd1778008, -32'sd1443078, -32'sd139757, -32'sd1507303, 32'sd730149, 32'sd1388738, -32'sd302245, -32'sd673522, -32'sd618913, -32'sd1253049, -32'sd913626, -32'sd348726, -32'sd277351, 32'sd617478, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd503359, 32'sd1042784, -32'sd273509, -32'sd278772, 32'sd154841, -32'sd637592, -32'sd455428, -32'sd226626, 32'sd343829, 32'sd30016, 32'sd218141, 32'sd258350, 32'sd277531, 32'sd998848, 32'sd1075441, 32'sd729961, 32'sd24387, -32'sd1212724, 32'sd1389689, 32'sd422439, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd952307, 32'sd932630, 32'sd405532, -32'sd950391, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1209019, 32'sd393942, -32'sd47883, 32'sd1781737, 32'sd1528755, -32'sd51009, -32'sd759754, 32'sd1315419, 32'sd236720, 32'sd396682, -32'sd836528, -32'sd178329, 32'sd1797762, 32'sd393315, -32'sd1287657, -32'sd138097, -32'sd690778, 32'sd337098, -32'sd203434, -32'sd166212, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15644, -32'sd12557, -32'sd22686, 32'sd1658084, 32'sd689004, 32'sd458552, 32'sd351997, 32'sd1034043, -32'sd1088448, 32'sd980768, 32'sd923520, -32'sd1151640, 32'sd4575, -32'sd1841323, 32'sd286950, -32'sd109400, 32'sd224334, -32'sd86949, 32'sd485790, -32'sd1145246, 32'sd855785, 32'sd200771, 32'sd730073, -32'sd587522, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd744488, 32'sd329500, -32'sd640216, -32'sd257447, 32'sd988161, -32'sd1377883, 32'sd524373, 32'sd640837, -32'sd1540284, 32'sd146833, 32'sd660911, -32'sd373976, 32'sd674, -32'sd1024364, -32'sd57061, 32'sd1419602, 32'sd2644972, -32'sd1482318, -32'sd1375522, -32'sd1873173, -32'sd2557290, -32'sd1746800, 32'sd333540, 32'sd637795, 32'sd856499, 32'sd0, 32'sd0, -32'sd369505, -32'sd323714, 32'sd620539, 32'sd1469936, 32'sd684486, 32'sd1694371, 32'sd919885, 32'sd279623, -32'sd1133878, -32'sd1164027, -32'sd1331306, -32'sd1387065, -32'sd1444227, -32'sd682627, 32'sd1227300, -32'sd576369, 32'sd1539938, 32'sd2008170, 32'sd291496, 32'sd280942, -32'sd539686, 32'sd674250, 32'sd381904, -32'sd1479049, 32'sd105730, 32'sd536730, -32'sd25028, 32'sd0, 32'sd320871, 32'sd249461, 32'sd187364, -32'sd726129, -32'sd140816, -32'sd1109682, 32'sd421821, 32'sd153240, -32'sd582431, -32'sd836336, 32'sd463559, -32'sd623010, 32'sd892172, 32'sd804820, -32'sd1635360, -32'sd1992136, 32'sd1074955, -32'sd306164, 32'sd1385, -32'sd578000, -32'sd1183247, -32'sd1034356, -32'sd1527977, -32'sd462775, 32'sd1683477, 32'sd1635335, -32'sd648362, 32'sd0, 32'sd416016, 32'sd21617, -32'sd1284637, -32'sd1522117, 32'sd222185, -32'sd588299, -32'sd288217, 32'sd826088, -32'sd1215124, 32'sd805670, 32'sd126510, -32'sd486924, -32'sd4386, -32'sd579687, -32'sd247633, -32'sd106355, 32'sd1030554, 32'sd392752, 32'sd918323, 32'sd2228226, 32'sd2269783, -32'sd69001, 32'sd436830, 32'sd862542, 32'sd978879, -32'sd1588465, 32'sd138761, 32'sd62007, 32'sd917492, -32'sd885826, -32'sd744203, -32'sd584131, 32'sd999589, -32'sd1350050, -32'sd1169547, 32'sd842632, -32'sd572312, -32'sd630411, -32'sd717072, -32'sd1971052, -32'sd17920, -32'sd511106, 32'sd1226179, 32'sd1753701, 32'sd2001257, 32'sd1544594, 32'sd2939531, 32'sd2405499, 32'sd1591311, 32'sd538419, 32'sd137744, 32'sd559933, 32'sd652643, -32'sd1332816, 32'sd287018, 32'sd48449, -32'sd1178257, 32'sd517325, 32'sd1023200, -32'sd97207, 32'sd303806, -32'sd3790, -32'sd43741, 32'sd971303, -32'sd169999, -32'sd614932, -32'sd725972, -32'sd459354, -32'sd1346107, -32'sd33346, 32'sd1655173, 32'sd3212735, 32'sd2201298, 32'sd1028644, 32'sd1532900, 32'sd1000306, 32'sd260515, 32'sd667338, -32'sd328797, 32'sd384229, -32'sd1393654, -32'sd710058, 32'sd491326, -32'sd558662, -32'sd835342, 32'sd489531, 32'sd1264756, -32'sd683331, -32'sd1550102, 32'sd681666, -32'sd770306, -32'sd120505, -32'sd117645, -32'sd1582770, 32'sd180116, 32'sd237976, 32'sd429896, -32'sd1072050, -32'sd2273087, -32'sd851894, 32'sd482629, -32'sd1254438, -32'sd342901, 32'sd142394, 32'sd1382759, -32'sd560201, 32'sd1410346, 32'sd423676, 32'sd817205, 32'sd139971, -32'sd845110, 32'sd62453, 32'sd77988, 32'sd266366, 32'sd932707, 32'sd145186, -32'sd362694, -32'sd1424790, -32'sd2615199, -32'sd2072317, -32'sd37923, -32'sd258706, -32'sd253130, 32'sd115530, -32'sd246021, -32'sd2836610, -32'sd2282100, -32'sd2995676, -32'sd4283915, -32'sd1582250, -32'sd2170108, 32'sd238686, -32'sd655463, -32'sd151604, -32'sd726444, -32'sd101449, 32'sd649053, 32'sd153519, 32'sd535146, 32'sd825011, -32'sd1129773, -32'sd926504, -32'sd1956162, -32'sd1313586, -32'sd713883, -32'sd912189, -32'sd774424, 32'sd954002, 32'sd1837633, 32'sd1085683, 32'sd1713243, -32'sd784629, -32'sd3730692, -32'sd653192, -32'sd1120659, -32'sd2610056, -32'sd842540, -32'sd1135447, 32'sd252720, 32'sd1628967, 32'sd2280279, 32'sd2164428, 32'sd3058711, 32'sd2533793, 32'sd1341008, -32'sd276402, 32'sd1710902, 32'sd907010, -32'sd1053314, -32'sd690890, -32'sd2316641, 32'sd709665, 32'sd1158435, 32'sd1412065, -32'sd648011, 32'sd992130, 32'sd2004671, 32'sd394667, -32'sd1823453, -32'sd1667482, -32'sd931532, -32'sd621352, -32'sd1300938, -32'sd1052796, -32'sd1061488, -32'sd178933, 32'sd96113, 32'sd1057698, 32'sd2953919, 32'sd1331216, 32'sd3060445, 32'sd291211, 32'sd1565346, 32'sd804004, 32'sd850994, 32'sd838327, -32'sd947567, 32'sd335350, -32'sd227374, 32'sd466703, -32'sd891388, -32'sd44950, -32'sd1235155, -32'sd7732, 32'sd966942, 32'sd792357, 32'sd985570, -32'sd93967, 32'sd50087, 32'sd616707, 32'sd96204, 32'sd133918, -32'sd417000, 32'sd1712454, 32'sd1096152, -32'sd596874, 32'sd42394, -32'sd1357857, 32'sd1086334, 32'sd851783, 32'sd272297, 32'sd65621, 32'sd837156, 32'sd128624, 32'sd1124511, -32'sd687900, -32'sd1687356, 32'sd537977, 32'sd570505, -32'sd649595, -32'sd487327, -32'sd417454, 32'sd1913586, 32'sd1542894, 32'sd1297097, 32'sd1098785, 32'sd1652536, 32'sd349595, 32'sd1509314, -32'sd1481638, -32'sd332969, 32'sd160517, -32'sd1428638, -32'sd706413, -32'sd505819, -32'sd2623795, -32'sd1164757, 32'sd198520, 32'sd705088, -32'sd86843, -32'sd1038580, -32'sd1061064, 32'sd249, -32'sd913311, -32'sd1773423, -32'sd392708, 32'sd1392876, 32'sd298806, 32'sd402961, 32'sd1515738, 32'sd1595177, 32'sd2801618, 32'sd2418157, 32'sd3346324, 32'sd1375969, 32'sd2786484, 32'sd54800, -32'sd1058819, -32'sd163557, -32'sd885178, -32'sd732192, -32'sd1735500, -32'sd3043511, -32'sd981382, -32'sd798165, 32'sd233474, -32'sd242550, 32'sd1490337, -32'sd666378, 32'sd850101, 32'sd1331879, -32'sd233042, 32'sd365938, -32'sd760456, -32'sd741933, 32'sd472599, -32'sd864757, -32'sd562487, 32'sd946395, 32'sd3773787, 32'sd2809460, 32'sd4326081, 32'sd2737769, 32'sd1816816, 32'sd213103, 32'sd786192, 32'sd248375, -32'sd1596395, -32'sd3081627, -32'sd2920235, -32'sd1608593, 32'sd140602, -32'sd999150, -32'sd443418, 32'sd407107, 32'sd258537, 32'sd704031, 32'sd0, -32'sd641524, -32'sd874209, -32'sd1786513, -32'sd1288071, -32'sd769496, 32'sd221456, -32'sd972705, -32'sd1062835, -32'sd1865009, 32'sd576686, 32'sd988479, 32'sd1415288, 32'sd2970343, 32'sd1164201, 32'sd2708702, -32'sd431571, -32'sd622673, -32'sd181526, -32'sd3826969, -32'sd586244, -32'sd1994988, -32'sd2047622, -32'sd2433199, 32'sd300825, 32'sd80147, 32'sd1010122, -32'sd825413, 32'sd523188, -32'sd197110, -32'sd1884266, -32'sd1137007, -32'sd1782305, -32'sd2495611, -32'sd1194407, -32'sd94306, -32'sd760061, -32'sd3702704, -32'sd1131802, -32'sd1422599, -32'sd1472202, 32'sd66369, -32'sd100834, 32'sd1931914, 32'sd1263327, -32'sd925569, -32'sd1594133, 32'sd6752, -32'sd1130776, 32'sd30604, -32'sd1071525, -32'sd1801774, -32'sd1680982, -32'sd289454, 32'sd218351, -32'sd436079, -32'sd152895, -32'sd45946, 32'sd83580, -32'sd505986, -32'sd1666148, -32'sd502635, -32'sd917565, -32'sd1453720, -32'sd1639448, -32'sd3040173, -32'sd2954285, -32'sd1078552, -32'sd428853, -32'sd1443446, -32'sd1508867, 32'sd1415295, 32'sd1785408, 32'sd1138983, 32'sd46402, -32'sd581870, -32'sd473159, 32'sd103443, -32'sd1871980, -32'sd2015689, 32'sd501163, 32'sd76644, 32'sd372062, -32'sd580942, 32'sd0, -32'sd791462, 32'sd918298, -32'sd260031, -32'sd721107, 32'sd1248928, 32'sd1569856, 32'sd211386, -32'sd192009, -32'sd2652452, -32'sd227485, -32'sd819111, -32'sd1850014, -32'sd1511332, -32'sd19800, -32'sd261340, -32'sd327421, 32'sd3568860, 32'sd1414221, 32'sd834788, 32'sd82980, 32'sd1135186, -32'sd1868118, -32'sd1042259, -32'sd1346918, -32'sd207152, -32'sd58187, 32'sd556986, 32'sd90055, 32'sd83879, 32'sd579174, -32'sd114312, 32'sd968407, -32'sd260884, 32'sd639844, 32'sd2017419, 32'sd618822, 32'sd225903, -32'sd882577, -32'sd1230635, -32'sd556513, -32'sd341379, 32'sd22690, 32'sd1350847, 32'sd92223, 32'sd2149103, -32'sd133938, -32'sd828907, -32'sd141322, -32'sd926214, -32'sd1104415, -32'sd1671707, -32'sd432310, -32'sd1544338, 32'sd192398, 32'sd7617, -32'sd253120, 32'sd450293, -32'sd426850, -32'sd516291, -32'sd186572, 32'sd18049, 32'sd1982312, 32'sd1934059, 32'sd272419, -32'sd40011, 32'sd908187, 32'sd44471, -32'sd906406, 32'sd748967, 32'sd2130571, 32'sd1359261, -32'sd1803203, 32'sd271040, -32'sd1763866, -32'sd456165, 32'sd66270, -32'sd2579401, -32'sd2090720, -32'sd642661, -32'sd540914, -32'sd772551, -32'sd272919, 32'sd926546, 32'sd0, 32'sd582308, 32'sd50755, -32'sd800717, -32'sd479268, -32'sd578667, -32'sd1224788, 32'sd1274701, 32'sd1969989, 32'sd1146214, -32'sd93933, 32'sd1704138, 32'sd1982949, 32'sd1986541, -32'sd70741, 32'sd874423, -32'sd893731, -32'sd751731, -32'sd330739, -32'sd341160, 32'sd741724, -32'sd907258, -32'sd161715, 32'sd67412, -32'sd524181, -32'sd844911, -32'sd576031, 32'sd0, 32'sd0, 32'sd0, 32'sd182477, -32'sd181814, -32'sd1442140, -32'sd857533, -32'sd381353, 32'sd507469, -32'sd676237, 32'sd1526119, 32'sd1745791, 32'sd1140986, 32'sd1358277, 32'sd2531708, -32'sd310040, 32'sd994887, 32'sd467881, -32'sd1545426, -32'sd1570212, -32'sd178550, 32'sd1092278, -32'sd657124, -32'sd401293, -32'sd549512, 32'sd871063, -32'sd172793, -32'sd40653, 32'sd0, 32'sd0, 32'sd0, 32'sd1784427, 32'sd689494, -32'sd1678171, -32'sd1510526, -32'sd67114, 32'sd917341, 32'sd328444, 32'sd1125858, -32'sd587686, 32'sd1035446, 32'sd2102717, 32'sd716126, 32'sd233978, -32'sd994966, -32'sd234501, 32'sd627375, 32'sd437233, 32'sd2246371, 32'sd19392, 32'sd1673283, 32'sd582685, 32'sd354538, 32'sd307224, -32'sd54249, 32'sd546300, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd380270, 32'sd1879578, 32'sd432149, 32'sd787763, 32'sd1036116, 32'sd1159324, 32'sd124238, 32'sd738411, -32'sd1123126, 32'sd2280443, 32'sd2581831, 32'sd2416251, 32'sd427383, 32'sd2004531, 32'sd1088875, 32'sd2032308, 32'sd1221860, 32'sd1349425, 32'sd359348, 32'sd304696, 32'sd1791516, -32'sd1399017, 32'sd18417, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd319959, 32'sd589645, -32'sd744928, 32'sd396019, -32'sd455330, 32'sd58579, 32'sd1333948, 32'sd1007130, -32'sd86373, 32'sd1110241, 32'sd1560870, 32'sd116194, 32'sd779092, 32'sd700478, 32'sd727292, 32'sd484043, 32'sd132003, -32'sd336846, -32'sd2045424, 32'sd247027, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd361924, -32'sd932046, -32'sd541203, -32'sd466958, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd94610, -32'sd380196, -32'sd418289, -32'sd144143, -32'sd564524, -32'sd161703, 32'sd429315, -32'sd1052420, -32'sd654275, -32'sd574734, -32'sd1366256, -32'sd201273, 32'sd586211, -32'sd422258, 32'sd349857, -32'sd61291, -32'sd52178, -32'sd388996, 32'sd179690, -32'sd468127, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd76756, 32'sd465039, -32'sd8479, -32'sd392548, 32'sd711315, 32'sd1041825, -32'sd813813, -32'sd1079100, 32'sd869554, -32'sd1154287, -32'sd1849596, 32'sd237156, 32'sd656996, -32'sd258461, -32'sd1545542, 32'sd126444, -32'sd925481, -32'sd2177296, -32'sd1176116, 32'sd187899, 32'sd349565, -32'sd980608, 32'sd397694, 32'sd703347, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd884911, -32'sd967973, 32'sd473559, -32'sd1337198, -32'sd459045, -32'sd81281, 32'sd526713, -32'sd1359542, 32'sd221500, 32'sd31898, -32'sd1114085, -32'sd1676779, -32'sd1301429, -32'sd973402, -32'sd1692583, -32'sd2936439, -32'sd1199854, -32'sd3115838, -32'sd801456, -32'sd1910126, -32'sd282240, 32'sd830934, 32'sd986963, 32'sd743104, -32'sd149945, 32'sd0, 32'sd0, 32'sd70848, -32'sd268254, 32'sd695959, 32'sd1205262, 32'sd207461, -32'sd851567, 32'sd969197, 32'sd470758, -32'sd526777, -32'sd235707, 32'sd772052, 32'sd1132599, 32'sd2219350, -32'sd1076367, -32'sd566219, -32'sd540315, -32'sd1266656, -32'sd2671399, -32'sd1243167, -32'sd2895592, -32'sd730152, -32'sd165824, -32'sd1034026, 32'sd141522, -32'sd687756, -32'sd293182, -32'sd472193, 32'sd0, -32'sd17520, 32'sd50660, 32'sd1076499, 32'sd1191840, 32'sd1096773, 32'sd143848, 32'sd1548227, -32'sd140492, -32'sd6488, 32'sd923136, 32'sd108930, 32'sd876249, -32'sd209998, -32'sd556818, 32'sd378520, -32'sd1644461, -32'sd3052986, -32'sd2240932, -32'sd2197465, -32'sd2356252, -32'sd3020750, -32'sd913020, 32'sd1580695, -32'sd1955024, 32'sd692262, -32'sd1084786, -32'sd722167, 32'sd0, 32'sd810314, 32'sd93392, 32'sd267710, 32'sd745452, 32'sd867806, 32'sd535554, 32'sd992080, 32'sd999757, 32'sd1525401, 32'sd1891237, 32'sd896779, -32'sd489390, 32'sd1023733, 32'sd940681, 32'sd1318099, -32'sd1198568, -32'sd326270, -32'sd285096, -32'sd1303226, -32'sd1263057, -32'sd283986, 32'sd1005403, -32'sd1101753, -32'sd1525721, -32'sd1935467, 32'sd1268803, -32'sd1381659, -32'sd280366, -32'sd1049000, 32'sd25112, 32'sd737428, 32'sd1834602, 32'sd832297, 32'sd1425231, 32'sd1095884, 32'sd1398808, 32'sd84528, 32'sd14902, -32'sd1088371, 32'sd1356782, 32'sd452521, 32'sd2735061, 32'sd70624, 32'sd781126, -32'sd1052132, -32'sd1015112, -32'sd958644, -32'sd770763, -32'sd1558452, -32'sd1687282, -32'sd2203457, -32'sd410391, 32'sd1141956, 32'sd855597, 32'sd382915, 32'sd653348, -32'sd791820, -32'sd955670, -32'sd338669, 32'sd1752538, 32'sd1635224, 32'sd5160, -32'sd2326008, 32'sd1962584, -32'sd464800, 32'sd745010, 32'sd673998, -32'sd672279, 32'sd2060785, 32'sd635744, -32'sd107602, -32'sd865292, 32'sd139734, -32'sd459908, -32'sd72964, -32'sd914484, -32'sd1410269, 32'sd102616, 32'sd182427, -32'sd865259, 32'sd1429819, -32'sd91642, -32'sd1396939, 32'sd1058935, -32'sd874304, 32'sd1155475, -32'sd137959, -32'sd123490, -32'sd286183, -32'sd1817151, 32'sd329156, 32'sd72274, 32'sd137070, -32'sd343401, -32'sd468957, 32'sd1798310, 32'sd3343190, 32'sd3802482, 32'sd1828372, -32'sd1158898, -32'sd1616740, -32'sd2074558, -32'sd366323, -32'sd1062952, 32'sd671245, 32'sd1646381, 32'sd1099047, -32'sd1696, -32'sd212619, 32'sd371083, 32'sd311288, 32'sd336439, -32'sd192197, -32'sd236541, 32'sd1268853, -32'sd1327935, -32'sd988432, -32'sd1618447, 32'sd694825, -32'sd733007, -32'sd2107223, -32'sd1329084, 32'sd2157783, 32'sd516100, 32'sd2176141, 32'sd1301103, -32'sd661146, -32'sd886224, -32'sd1600487, -32'sd840816, -32'sd1458753, 32'sd1422113, 32'sd1131119, -32'sd532308, 32'sd2238781, 32'sd1189565, -32'sd405251, 32'sd296096, 32'sd1285405, -32'sd708325, -32'sd1378542, 32'sd300363, 32'sd2262059, -32'sd313887, -32'sd1224554, -32'sd95203, 32'sd154525, 32'sd235394, -32'sd1528560, 32'sd1604790, 32'sd754422, -32'sd1378976, -32'sd435836, 32'sd152777, -32'sd965284, -32'sd1294061, -32'sd609668, -32'sd1382338, 32'sd70164, 32'sd1972539, 32'sd698700, -32'sd640411, 32'sd428805, -32'sd2237814, 32'sd830304, 32'sd541729, 32'sd188783, 32'sd493281, -32'sd433878, 32'sd229133, 32'sd357805, 32'sd818453, -32'sd284236, 32'sd1233111, -32'sd2048334, 32'sd231613, -32'sd286154, -32'sd331751, -32'sd2147039, -32'sd4367935, -32'sd1102537, 32'sd589359, 32'sd211817, 32'sd55675, 32'sd196110, 32'sd848304, 32'sd880835, 32'sd1985069, 32'sd313266, -32'sd1051390, 32'sd364796, -32'sd103644, 32'sd496713, -32'sd1175386, -32'sd447961, -32'sd285195, 32'sd1395425, 32'sd1258984, 32'sd1113974, -32'sd1427478, -32'sd1605683, 32'sd1745208, -32'sd892635, -32'sd561005, 32'sd178648, -32'sd2539949, -32'sd3427685, -32'sd2386838, 32'sd439956, 32'sd3266406, 32'sd2075188, 32'sd1504177, 32'sd2654962, 32'sd2986560, 32'sd506812, 32'sd125651, -32'sd475086, -32'sd1499130, -32'sd334066, -32'sd752891, 32'sd161695, -32'sd585397, -32'sd376332, -32'sd441013, -32'sd759515, 32'sd1677624, -32'sd2689194, -32'sd798247, -32'sd1613924, -32'sd1749708, 32'sd1415068, -32'sd361708, -32'sd2112370, -32'sd3852452, -32'sd854512, 32'sd1870534, 32'sd2123189, 32'sd3421502, 32'sd3317160, 32'sd2513804, 32'sd2364808, 32'sd280712, 32'sd844182, -32'sd40359, 32'sd848524, -32'sd2726026, -32'sd1207918, 32'sd190552, 32'sd184239, 32'sd2278080, 32'sd460376, -32'sd848567, 32'sd1076763, 32'sd871187, -32'sd835570, -32'sd1990998, 32'sd410706, -32'sd504050, -32'sd1963782, -32'sd2140313, -32'sd3003629, -32'sd1399946, -32'sd927822, 32'sd1629144, 32'sd3520528, 32'sd4399367, 32'sd1249734, 32'sd3948618, 32'sd2255326, -32'sd1245480, 32'sd346105, 32'sd2276759, -32'sd491152, -32'sd2064433, -32'sd716573, -32'sd1439296, 32'sd550150, 32'sd1125603, 32'sd1130980, 32'sd56460, -32'sd947656, 32'sd639247, 32'sd643369, 32'sd1873159, 32'sd921596, -32'sd981742, 32'sd1279897, -32'sd1678257, 32'sd350370, 32'sd576422, 32'sd1308, 32'sd3587826, 32'sd3992186, 32'sd1419848, 32'sd372059, 32'sd91413, -32'sd1222896, -32'sd143632, -32'sd88764, 32'sd775112, 32'sd735373, -32'sd508921, -32'sd1358733, 32'sd172982, -32'sd122125, -32'sd354657, -32'sd494191, 32'sd0, 32'sd977725, -32'sd957845, 32'sd902996, 32'sd1548458, 32'sd1662216, -32'sd491061, -32'sd384654, -32'sd170551, -32'sd2281021, -32'sd2039760, -32'sd1323947, 32'sd1778996, 32'sd283186, 32'sd82478, -32'sd346530, -32'sd2497770, -32'sd2072285, -32'sd2686991, -32'sd711555, 32'sd477016, -32'sd721827, -32'sd2797505, -32'sd1133985, 32'sd581451, 32'sd620027, 32'sd566449, 32'sd162559, -32'sd1153275, -32'sd173735, 32'sd1068346, -32'sd1495774, 32'sd1422788, 32'sd743618, -32'sd1184672, -32'sd942226, -32'sd2147378, -32'sd2146111, -32'sd2678944, -32'sd667579, -32'sd822480, -32'sd1295615, -32'sd1598283, -32'sd1785015, -32'sd600090, -32'sd2126134, -32'sd1226926, -32'sd1220142, -32'sd674926, -32'sd795168, -32'sd1067403, 32'sd247304, -32'sd1190699, -32'sd1372324, -32'sd1825676, -32'sd1309927, -32'sd45600, 32'sd669624, -32'sd536182, -32'sd1281847, 32'sd1583407, 32'sd430162, -32'sd1443133, -32'sd2350520, -32'sd948186, -32'sd322089, 32'sd561390, -32'sd2691739, -32'sd3257862, -32'sd2647130, -32'sd1263285, -32'sd1913962, 32'sd914979, -32'sd1397007, -32'sd617274, -32'sd243991, -32'sd1017094, 32'sd670256, -32'sd835090, 32'sd83985, -32'sd543381, 32'sd752000, -32'sd1514850, 32'sd171757, 32'sd0, 32'sd849114, -32'sd317096, 32'sd1266086, -32'sd406082, -32'sd378220, 32'sd455607, 32'sd792993, -32'sd386222, 32'sd25293, -32'sd2236417, -32'sd1713561, -32'sd978519, -32'sd1420185, 32'sd635454, -32'sd1590489, -32'sd1946251, 32'sd216993, 32'sd1133939, 32'sd7440, 32'sd547552, 32'sd401733, -32'sd371188, -32'sd312642, -32'sd1335526, -32'sd462216, -32'sd805421, -32'sd471778, -32'sd45017, 32'sd823251, -32'sd968947, 32'sd1133190, 32'sd1273605, 32'sd2022353, 32'sd1166506, 32'sd1045761, 32'sd255628, -32'sd774340, 32'sd1113104, -32'sd109560, -32'sd1655362, -32'sd1478862, -32'sd1652363, -32'sd1782347, -32'sd945502, -32'sd2981196, -32'sd64954, -32'sd453739, 32'sd565750, -32'sd1222112, -32'sd1102231, -32'sd1477274, -32'sd1995061, -32'sd48598, -32'sd902938, 32'sd1184815, -32'sd443659, 32'sd532469, -32'sd485573, -32'sd557987, 32'sd1835697, -32'sd104278, -32'sd573031, 32'sd899457, 32'sd645885, 32'sd549435, 32'sd124863, -32'sd1825734, -32'sd404160, -32'sd675604, 32'sd209290, -32'sd499580, -32'sd2014950, -32'sd710416, 32'sd1435995, -32'sd593981, -32'sd531527, -32'sd573020, 32'sd445006, -32'sd1506312, 32'sd823401, 32'sd397057, 32'sd730684, 32'sd781819, 32'sd0, -32'sd530508, 32'sd358021, 32'sd340522, 32'sd299855, 32'sd742392, 32'sd241376, 32'sd1411834, -32'sd598955, 32'sd448797, -32'sd955411, -32'sd943836, 32'sd545324, -32'sd894965, 32'sd739603, 32'sd972372, -32'sd472489, -32'sd505191, 32'sd495437, -32'sd630908, -32'sd1487349, -32'sd205872, -32'sd238062, -32'sd1793056, 32'sd1327241, -32'sd445887, 32'sd1302290, 32'sd0, 32'sd0, 32'sd0, -32'sd1152161, 32'sd404505, -32'sd1205886, 32'sd191355, 32'sd821978, -32'sd84119, -32'sd360188, -32'sd1030096, 32'sd754175, -32'sd831593, -32'sd2691571, -32'sd427295, 32'sd820437, -32'sd625715, 32'sd1712, 32'sd1381878, 32'sd2064753, 32'sd1267031, 32'sd1568620, 32'sd93021, 32'sd167251, -32'sd1992976, 32'sd153408, -32'sd1168672, 32'sd894168, 32'sd0, 32'sd0, 32'sd0, 32'sd1517777, 32'sd330770, 32'sd33061, 32'sd2195232, -32'sd572940, 32'sd2307980, 32'sd1727349, 32'sd860521, -32'sd619462, -32'sd619169, -32'sd705802, 32'sd1297558, 32'sd705193, -32'sd934712, -32'sd146797, -32'sd129848, -32'sd1324292, -32'sd747119, 32'sd842214, 32'sd1643116, -32'sd866236, 32'sd553218, -32'sd470365, -32'sd106041, 32'sd362473, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd535973, 32'sd1728987, 32'sd1554270, -32'sd234431, 32'sd2969019, 32'sd773057, 32'sd1839307, 32'sd872643, 32'sd1633276, 32'sd1431798, -32'sd338211, -32'sd139368, -32'sd2012289, -32'sd377180, 32'sd771267, -32'sd747144, -32'sd383056, 32'sd529330, 32'sd908995, 32'sd529346, -32'sd20707, -32'sd863134, 32'sd48262, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd730618, -32'sd381829, -32'sd613733, -32'sd153423, 32'sd93032, -32'sd773955, 32'sd1291779, -32'sd609358, 32'sd1022331, -32'sd87754, 32'sd1794794, -32'sd296862, -32'sd116922, 32'sd808896, 32'sd830403, -32'sd1484251, 32'sd826569, -32'sd777596, -32'sd1434722, -32'sd185066, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd83063, 32'sd1122243, 32'sd722612, 32'sd1798884, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd724494, -32'sd143304, -32'sd552929, -32'sd920983, -32'sd1053285, -32'sd647469, 32'sd712108, 32'sd1702931, -32'sd610479, -32'sd369129, -32'sd479304, 32'sd1294225, 32'sd636138, 32'sd783403, -32'sd830108, -32'sd273024, 32'sd1093572, 32'sd1131796, -32'sd1120009, 32'sd1369403, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1457694, -32'sd273068, -32'sd1565419, 32'sd183994, -32'sd205147, 32'sd765980, 32'sd475306, 32'sd46554, 32'sd2449350, 32'sd779349, 32'sd717685, 32'sd454813, 32'sd759059, 32'sd704733, 32'sd1971238, -32'sd118736, 32'sd972507, 32'sd2327427, 32'sd2081982, 32'sd565157, 32'sd219931, -32'sd962173, 32'sd1153419, 32'sd929545, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd981416, 32'sd365367, 32'sd1205360, 32'sd435010, 32'sd1179978, 32'sd778117, 32'sd160314, 32'sd1039405, -32'sd45009, 32'sd14127, 32'sd1209116, 32'sd337351, -32'sd327552, 32'sd2131059, 32'sd135714, 32'sd839232, 32'sd3902649, 32'sd2178664, -32'sd723314, 32'sd899102, 32'sd2328681, 32'sd285179, 32'sd894138, 32'sd546133, 32'sd218866, 32'sd0, 32'sd0, 32'sd200535, 32'sd775109, 32'sd1502869, 32'sd116223, -32'sd702873, 32'sd601181, -32'sd3473, 32'sd2207109, 32'sd1127292, 32'sd1378077, 32'sd250548, 32'sd179623, 32'sd1515910, -32'sd282432, 32'sd1592408, 32'sd2118809, 32'sd873882, 32'sd2424842, 32'sd1764808, 32'sd492390, 32'sd1352021, -32'sd345708, -32'sd2718263, 32'sd793580, 32'sd1315257, -32'sd492345, 32'sd586039, 32'sd0, 32'sd1298423, 32'sd1104026, 32'sd1286665, -32'sd724822, 32'sd2411508, -32'sd294897, 32'sd643069, 32'sd1882040, 32'sd2116641, 32'sd1892551, -32'sd693918, -32'sd1074430, -32'sd63835, -32'sd307702, 32'sd621130, 32'sd877473, 32'sd1133144, 32'sd3385044, 32'sd283024, 32'sd1488917, 32'sd208737, 32'sd92413, 32'sd1748674, 32'sd1065629, -32'sd929763, -32'sd1364603, 32'sd405002, 32'sd0, 32'sd385137, 32'sd311373, 32'sd932930, 32'sd330441, -32'sd743031, -32'sd121587, 32'sd1478030, 32'sd651575, 32'sd2639657, 32'sd3341358, 32'sd110242, 32'sd1492039, 32'sd1205067, 32'sd804753, 32'sd1489538, -32'sd643427, -32'sd556100, 32'sd1005773, 32'sd1812478, -32'sd849745, 32'sd918648, 32'sd667647, -32'sd463439, 32'sd579658, 32'sd714166, 32'sd810211, -32'sd1356612, 32'sd1512308, 32'sd1081562, 32'sd30675, 32'sd1363020, -32'sd178563, -32'sd1202974, -32'sd80972, 32'sd445883, -32'sd1003, 32'sd309981, 32'sd424334, 32'sd218605, 32'sd723495, 32'sd926580, 32'sd1241385, -32'sd590655, 32'sd198603, 32'sd814463, 32'sd1254501, 32'sd3002276, 32'sd945189, 32'sd2265418, 32'sd542253, 32'sd1998483, -32'sd920085, 32'sd1736359, 32'sd124237, 32'sd768320, 32'sd650984, 32'sd869841, 32'sd411117, -32'sd244530, -32'sd41880, -32'sd411351, -32'sd959473, 32'sd808220, -32'sd1110974, -32'sd775727, -32'sd1201467, -32'sd682472, 32'sd129618, -32'sd1577482, -32'sd1615785, -32'sd1311535, 32'sd1097278, 32'sd1795475, 32'sd195084, 32'sd3674814, 32'sd108321, 32'sd699232, -32'sd94749, 32'sd88401, -32'sd630440, 32'sd144727, 32'sd2228519, 32'sd1105837, -32'sd157838, -32'sd469969, -32'sd986281, 32'sd708297, 32'sd1362107, 32'sd96220, 32'sd773683, 32'sd399037, -32'sd482080, 32'sd25316, -32'sd1538145, -32'sd3638299, -32'sd2175846, -32'sd3372557, -32'sd4246872, -32'sd2779451, 32'sd796406, 32'sd3168728, 32'sd627833, 32'sd1509931, -32'sd552262, -32'sd1831973, 32'sd1087183, 32'sd430271, -32'sd2014121, -32'sd1014217, -32'sd63882, 32'sd535559, 32'sd877526, 32'sd173788, 32'sd634427, 32'sd858143, 32'sd1760978, -32'sd2676389, -32'sd1724275, -32'sd3162229, -32'sd884077, -32'sd1535061, -32'sd4449735, -32'sd5048791, -32'sd3835345, -32'sd5737860, -32'sd4457275, -32'sd2907841, 32'sd3628716, 32'sd2517013, 32'sd692365, 32'sd1592833, -32'sd557036, -32'sd749505, 32'sd164938, -32'sd1462194, -32'sd774289, 32'sd409630, 32'sd1457432, 32'sd737291, -32'sd250196, -32'sd752392, 32'sd535805, -32'sd155873, -32'sd1313976, -32'sd2462360, -32'sd2443862, -32'sd3701008, -32'sd4768471, -32'sd3962394, -32'sd3654993, -32'sd4207576, -32'sd2761086, -32'sd3886785, -32'sd3824126, -32'sd349788, 32'sd2421395, 32'sd1567049, 32'sd1573336, 32'sd974350, -32'sd161836, 32'sd475802, -32'sd473602, -32'sd48952, -32'sd655844, 32'sd882428, 32'sd237226, -32'sd117353, 32'sd818090, -32'sd13490, -32'sd942181, 32'sd368523, -32'sd1408169, -32'sd1718347, -32'sd3484274, -32'sd4108104, -32'sd3325142, -32'sd2572124, 32'sd461703, -32'sd261721, -32'sd1755355, -32'sd594237, -32'sd61803, 32'sd3431402, 32'sd3038632, 32'sd77847, 32'sd1916134, 32'sd92525, -32'sd1699568, 32'sd31172, -32'sd397928, 32'sd798315, -32'sd2224016, 32'sd118138, 32'sd317202, 32'sd92944, 32'sd1284334, -32'sd347846, -32'sd586909, -32'sd1732951, 32'sd593844, -32'sd900314, 32'sd301037, 32'sd50315, 32'sd734019, -32'sd671313, 32'sd833100, -32'sd409555, 32'sd102687, 32'sd497515, 32'sd781831, 32'sd1106002, 32'sd1701313, 32'sd1522092, 32'sd577069, 32'sd445745, -32'sd616787, -32'sd94306, -32'sd1267241, -32'sd1313844, -32'sd579850, 32'sd134342, -32'sd256530, 32'sd1145254, 32'sd904717, -32'sd649151, -32'sd278738, 32'sd204682, 32'sd1393535, 32'sd934713, 32'sd2543249, 32'sd853307, 32'sd322559, 32'sd1883605, 32'sd1517184, 32'sd66023, -32'sd626110, -32'sd274614, 32'sd1534287, 32'sd2659091, 32'sd3414906, 32'sd2956048, 32'sd2194007, -32'sd2203300, -32'sd1542548, -32'sd331240, 32'sd878420, -32'sd1168664, -32'sd508968, -32'sd773743, 32'sd256547, 32'sd1225611, 32'sd816710, 32'sd859796, -32'sd489515, 32'sd1440861, 32'sd291134, 32'sd1571148, 32'sd1601963, -32'sd1660042, -32'sd453334, 32'sd798333, 32'sd297606, -32'sd1703140, -32'sd1654308, -32'sd1361615, 32'sd178874, 32'sd2831848, 32'sd757299, 32'sd743772, 32'sd1585566, -32'sd1518979, -32'sd1907960, -32'sd2232514, -32'sd1009305, -32'sd589187, -32'sd800600, 32'sd192062, -32'sd566016, 32'sd984806, 32'sd1151598, 32'sd264519, -32'sd1007180, 32'sd384477, 32'sd912579, 32'sd923768, -32'sd754884, -32'sd835616, -32'sd4310048, -32'sd677023, -32'sd1000522, -32'sd363114, -32'sd2782823, -32'sd1334978, 32'sd41261, 32'sd3233547, 32'sd1059507, -32'sd641675, 32'sd1445387, -32'sd1488211, 32'sd396784, -32'sd173725, -32'sd1287393, -32'sd717591, 32'sd630655, 32'sd1019946, -32'sd663877, -32'sd381168, 32'sd0, 32'sd1814400, -32'sd59535, -32'sd179337, -32'sd457410, 32'sd141383, -32'sd2257001, -32'sd561968, -32'sd2850743, -32'sd2495255, -32'sd589211, 32'sd1140540, -32'sd1068465, -32'sd358995, 32'sd2176437, 32'sd2740438, 32'sd470428, 32'sd287379, -32'sd356619, 32'sd450825, -32'sd1281465, -32'sd103348, -32'sd718195, -32'sd469872, 32'sd926442, 32'sd1326139, 32'sd2349916, 32'sd776888, -32'sd600279, -32'sd816326, 32'sd886702, 32'sd1034797, -32'sd1621303, -32'sd978862, -32'sd1224133, -32'sd1039031, -32'sd1206460, -32'sd125022, -32'sd994871, 32'sd1737472, -32'sd447865, -32'sd654468, 32'sd905577, 32'sd119225, 32'sd1772619, 32'sd1475335, 32'sd1323530, 32'sd123714, -32'sd2067938, -32'sd1911727, -32'sd787407, 32'sd1518909, 32'sd1702751, 32'sd742532, 32'sd805471, 32'sd1091388, 32'sd1630581, 32'sd1012013, 32'sd479315, 32'sd1541563, 32'sd594551, -32'sd1201875, 32'sd451613, 32'sd2125348, 32'sd644017, 32'sd1387558, 32'sd1152634, 32'sd2699539, 32'sd1772048, -32'sd269854, -32'sd101241, 32'sd555257, 32'sd1540275, 32'sd917056, -32'sd1313496, 32'sd888281, -32'sd210729, -32'sd135334, -32'sd483920, -32'sd163615, 32'sd910384, 32'sd1586925, 32'sd2011472, 32'sd1128700, 32'sd0, -32'sd864807, 32'sd204823, -32'sd124458, -32'sd388186, 32'sd701147, -32'sd219537, 32'sd279003, 32'sd804292, -32'sd12984, 32'sd2377236, 32'sd804251, 32'sd3053887, -32'sd696397, -32'sd117878, -32'sd1186160, 32'sd2226240, 32'sd708603, -32'sd320672, -32'sd111960, -32'sd51563, 32'sd2035136, -32'sd1028557, -32'sd393388, -32'sd181431, 32'sd1166393, 32'sd2536811, 32'sd1029354, 32'sd410671, 32'sd1341874, 32'sd762110, 32'sd1571110, 32'sd819398, -32'sd1026457, 32'sd739504, 32'sd2394635, 32'sd823842, -32'sd50589, 32'sd2206940, 32'sd2294770, 32'sd268012, -32'sd294827, -32'sd391967, -32'sd2068272, 32'sd915182, 32'sd25342, 32'sd361601, 32'sd561250, -32'sd564955, 32'sd2146179, -32'sd1025059, 32'sd776894, 32'sd890123, 32'sd660455, 32'sd728274, 32'sd596449, 32'sd1939208, -32'sd422121, 32'sd697720, 32'sd690537, -32'sd1070543, 32'sd1508489, -32'sd474793, 32'sd1559783, 32'sd2089321, -32'sd442112, 32'sd335340, -32'sd1063079, 32'sd14565, -32'sd1046152, -32'sd911079, 32'sd1108481, 32'sd1327690, -32'sd858679, -32'sd199275, -32'sd847370, -32'sd451416, 32'sd17200, 32'sd715711, 32'sd1721083, 32'sd251690, -32'sd137464, -32'sd1108021, 32'sd1610410, 32'sd0, 32'sd795468, -32'sd974436, 32'sd624963, -32'sd298941, 32'sd1750880, -32'sd11345, 32'sd499565, -32'sd1489996, 32'sd1425625, -32'sd1720947, -32'sd255739, -32'sd1469436, 32'sd1672981, -32'sd833685, -32'sd727936, 32'sd973312, 32'sd269161, -32'sd1521685, 32'sd162971, -32'sd1092366, -32'sd496767, -32'sd67952, 32'sd160222, 32'sd953477, 32'sd1593730, -32'sd1153633, 32'sd0, 32'sd0, 32'sd0, 32'sd2236417, -32'sd390327, 32'sd1969283, 32'sd256482, -32'sd29237, -32'sd741258, 32'sd1525776, -32'sd752309, -32'sd1939544, -32'sd1793542, -32'sd710269, -32'sd63170, 32'sd438123, 32'sd1135816, -32'sd1407212, -32'sd431755, -32'sd2066439, -32'sd3917777, -32'sd1658454, -32'sd245888, -32'sd2080141, -32'sd112939, 32'sd1312203, -32'sd339788, 32'sd163010, 32'sd0, 32'sd0, 32'sd0, 32'sd935826, 32'sd318258, 32'sd2329839, 32'sd1098056, 32'sd604307, 32'sd2508161, 32'sd1703585, -32'sd295594, -32'sd2016067, 32'sd292182, -32'sd242595, 32'sd568609, 32'sd692983, -32'sd2441902, 32'sd153473, 32'sd1187498, -32'sd1181336, -32'sd1652458, -32'sd1010987, -32'sd103452, 32'sd232145, 32'sd769286, -32'sd253506, -32'sd337572, -32'sd61154, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1556570, -32'sd4466, -32'sd459624, 32'sd58023, 32'sd1789844, 32'sd1834592, -32'sd149999, 32'sd433149, 32'sd3371984, 32'sd823214, -32'sd673185, 32'sd2765663, 32'sd227481, 32'sd1106289, 32'sd2548299, 32'sd802938, -32'sd770987, 32'sd257517, -32'sd346865, -32'sd1565967, -32'sd730120, 32'sd819477, 32'sd1304118, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1359985, 32'sd790377, 32'sd1598829, 32'sd1950525, 32'sd1000967, 32'sd981168, 32'sd2356546, 32'sd967919, 32'sd1442898, 32'sd2100873, 32'sd2273331, 32'sd637845, 32'sd1294085, 32'sd2325526, 32'sd1049009, 32'sd247193, 32'sd736915, 32'sd127293, -32'sd155857, 32'sd884615, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd940827, 32'sd1330343, 32'sd1101478, 32'sd19520, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1638848, 32'sd741916, 32'sd1344196, 32'sd767862, -32'sd92591, -32'sd519812, 32'sd1649253, 32'sd1271297, 32'sd1999155, 32'sd1158508, 32'sd74145, -32'sd576430, 32'sd348961, 32'sd1129117, 32'sd961624, -32'sd216982, 32'sd1518881, -32'sd27203, 32'sd1320630, 32'sd539631, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd582083, 32'sd487030, 32'sd144341, 32'sd97811, 32'sd570937, 32'sd973375, 32'sd1528245, 32'sd1624056, 32'sd2737011, 32'sd1495793, -32'sd568641, -32'sd120280, 32'sd528433, -32'sd23982, 32'sd156056, -32'sd65734, 32'sd974480, 32'sd742169, -32'sd707864, 32'sd1504848, 32'sd740013, -32'sd1365621, 32'sd608735, 32'sd402853, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1333481, 32'sd867147, 32'sd686273, -32'sd88405, 32'sd2164457, 32'sd562004, -32'sd619859, 32'sd1064254, 32'sd1044250, -32'sd513635, -32'sd2833355, -32'sd308523, -32'sd487635, 32'sd477371, 32'sd1302921, 32'sd1397609, -32'sd1485435, -32'sd640679, -32'sd2731510, -32'sd757815, 32'sd878314, 32'sd609662, -32'sd424648, -32'sd629078, -32'sd117846, 32'sd0, 32'sd0, -32'sd123541, 32'sd229236, -32'sd474322, -32'sd558464, -32'sd440514, 32'sd538736, -32'sd2044651, -32'sd35872, 32'sd19888, -32'sd23498, -32'sd592179, -32'sd2149893, -32'sd1477315, -32'sd1318501, -32'sd1520284, 32'sd1927370, 32'sd724084, -32'sd1568276, -32'sd424762, -32'sd1473888, -32'sd1939653, -32'sd2911111, -32'sd1954481, 32'sd1069796, 32'sd558762, 32'sd104635, -32'sd288974, 32'sd0, 32'sd1214650, 32'sd1132152, 32'sd348174, 32'sd938965, -32'sd1880613, 32'sd151631, 32'sd1152074, 32'sd966764, 32'sd948953, 32'sd844588, 32'sd765254, 32'sd808575, -32'sd1234379, -32'sd2134455, -32'sd1959001, 32'sd878203, -32'sd30715, -32'sd1924824, -32'sd781755, -32'sd586783, -32'sd423660, 32'sd1590548, -32'sd329176, 32'sd888553, -32'sd551660, -32'sd1496903, 32'sd808361, 32'sd0, 32'sd298594, -32'sd903561, 32'sd532570, -32'sd539345, -32'sd1659829, 32'sd936450, 32'sd1442453, 32'sd2735875, 32'sd1555168, -32'sd1226288, -32'sd1055558, -32'sd665243, -32'sd1503205, 32'sd560763, -32'sd685706, -32'sd1381573, -32'sd856173, -32'sd614644, -32'sd1219375, -32'sd697583, 32'sd829999, 32'sd614486, -32'sd782614, -32'sd2880748, 32'sd182967, 32'sd19258, 32'sd962674, 32'sd569522, 32'sd1948531, -32'sd1090975, -32'sd300070, 32'sd924480, -32'sd318819, -32'sd295838, 32'sd1703857, 32'sd2893828, 32'sd1656823, -32'sd1307990, -32'sd1035229, -32'sd1450705, -32'sd410584, 32'sd26449, 32'sd238739, -32'sd2072516, 32'sd643463, -32'sd1345390, 32'sd1433468, 32'sd295443, -32'sd577851, -32'sd2534409, -32'sd2540638, -32'sd1390444, 32'sd270763, 32'sd409015, -32'sd54918, 32'sd1439406, 32'sd833465, -32'sd1100688, -32'sd448283, 32'sd1999345, -32'sd1368113, 32'sd1674345, 32'sd3208553, 32'sd126002, 32'sd2217741, -32'sd816078, -32'sd2359060, -32'sd1665655, 32'sd1483659, 32'sd17105, -32'sd766657, 32'sd992493, -32'sd794075, -32'sd1373254, 32'sd1283145, 32'sd1176623, 32'sd1571277, -32'sd1656202, -32'sd1401702, 32'sd980498, -32'sd420867, 32'sd108325, -32'sd278385, 32'sd1396699, -32'sd619155, -32'sd1773238, 32'sd357348, 32'sd2581059, 32'sd435967, -32'sd837623, 32'sd683773, 32'sd936028, 32'sd349209, 32'sd992516, -32'sd1712392, 32'sd466521, -32'sd364007, -32'sd881463, -32'sd23731, 32'sd2095722, 32'sd2028892, -32'sd1195942, -32'sd131335, 32'sd1733311, -32'sd824868, -32'sd416916, -32'sd1429082, -32'sd1023012, -32'sd1011337, -32'sd741333, 32'sd155977, 32'sd738320, 32'sd1221629, 32'sd531260, -32'sd229283, -32'sd537324, 32'sd265486, 32'sd720333, 32'sd733122, 32'sd1677626, 32'sd1374994, -32'sd138332, -32'sd29879, -32'sd1127022, -32'sd640193, -32'sd1590563, 32'sd291689, 32'sd717949, -32'sd99920, -32'sd1430764, -32'sd1648784, 32'sd219006, -32'sd1002916, -32'sd299396, -32'sd2745287, 32'sd155517, -32'sd1292432, 32'sd104797, -32'sd1531691, -32'sd435700, -32'sd1291795, 32'sd109743, 32'sd859487, 32'sd1098133, 32'sd1449503, 32'sd8905, 32'sd527928, 32'sd936244, 32'sd1207003, 32'sd327320, -32'sd1208302, -32'sd1359147, -32'sd927412, 32'sd309133, 32'sd1560645, 32'sd2222146, 32'sd346461, -32'sd750420, 32'sd192760, 32'sd630365, -32'sd710715, -32'sd18649, -32'sd2710523, -32'sd3044470, 32'sd1279887, 32'sd217591, -32'sd1663108, 32'sd1510308, -32'sd906303, 32'sd1110031, -32'sd671075, 32'sd1832026, -32'sd34391, -32'sd2678577, 32'sd384791, 32'sd1278397, 32'sd449655, -32'sd1479672, -32'sd548647, -32'sd3060579, 32'sd815683, 32'sd418941, 32'sd3477992, 32'sd318348, -32'sd672957, 32'sd114670, -32'sd780440, 32'sd265105, 32'sd745111, -32'sd236772, -32'sd3083903, -32'sd1573482, 32'sd1002817, -32'sd602344, -32'sd348894, 32'sd666039, -32'sd1187413, 32'sd834074, 32'sd1828829, 32'sd397314, 32'sd1312556, -32'sd485397, -32'sd809083, 32'sd329118, -32'sd1294389, -32'sd1191041, -32'sd298032, -32'sd152416, 32'sd2263605, 32'sd404023, 32'sd2660391, -32'sd1349752, -32'sd1193082, 32'sd1181732, 32'sd156731, 32'sd315362, 32'sd584985, 32'sd674838, -32'sd303327, -32'sd1671641, 32'sd982155, 32'sd149370, 32'sd506577, -32'sd185918, 32'sd77645, -32'sd848971, 32'sd846419, 32'sd2075314, 32'sd439242, 32'sd238949, -32'sd2328570, -32'sd664079, -32'sd899474, -32'sd2588472, -32'sd744598, 32'sd157307, 32'sd2981260, 32'sd2445436, -32'sd1171565, -32'sd2075189, 32'sd927765, 32'sd2159394, 32'sd2691168, 32'sd646706, -32'sd1376549, -32'sd1406052, 32'sd1899656, -32'sd643056, 32'sd180854, 32'sd921324, 32'sd787815, -32'sd42047, 32'sd507901, -32'sd616501, 32'sd153783, -32'sd642051, -32'sd2078894, -32'sd400186, -32'sd1232962, -32'sd1368180, -32'sd1944081, -32'sd1798812, 32'sd1446774, 32'sd1225177, 32'sd3319998, 32'sd2162483, -32'sd273539, -32'sd1524586, -32'sd2089760, 32'sd465774, 32'sd841773, 32'sd1299506, 32'sd201433, -32'sd384334, 32'sd2123839, 32'sd1326128, -32'sd720824, 32'sd644770, 32'sd329853, 32'sd1054148, 32'sd1303415, -32'sd764955, 32'sd1351192, -32'sd1528889, 32'sd694350, 32'sd210607, -32'sd1140338, -32'sd2367394, -32'sd4110842, -32'sd1763385, 32'sd2356753, 32'sd2041949, 32'sd1760618, 32'sd2273731, 32'sd559758, -32'sd57429, -32'sd949602, -32'sd1565900, 32'sd960326, 32'sd1190400, -32'sd1123600, 32'sd1964889, 32'sd3004646, 32'sd692923, 32'sd190452, -32'sd642856, -32'sd363315, 32'sd0, -32'sd1115846, 32'sd654864, 32'sd957034, 32'sd380102, -32'sd1147087, -32'sd1968027, -32'sd1343777, -32'sd5121618, -32'sd3174652, 32'sd1908667, 32'sd2255238, 32'sd4013959, 32'sd1116148, -32'sd374354, 32'sd693733, 32'sd444495, 32'sd1973664, 32'sd984175, 32'sd1899518, 32'sd699996, 32'sd52796, -32'sd742245, 32'sd676105, -32'sd696983, -32'sd465627, -32'sd925390, -32'sd311637, 32'sd427221, 32'sd246296, -32'sd171084, -32'sd282104, -32'sd1160644, -32'sd242491, -32'sd2430627, -32'sd2826401, -32'sd3431269, -32'sd314512, 32'sd2696430, 32'sd3125733, 32'sd4167277, 32'sd3640476, -32'sd560539, 32'sd462609, -32'sd688417, -32'sd97273, 32'sd1575074, -32'sd49183, -32'sd494482, 32'sd100673, -32'sd555266, -32'sd3344767, -32'sd160823, -32'sd567854, -32'sd704768, -32'sd392844, 32'sd987917, 32'sd230611, -32'sd1699362, -32'sd839761, 32'sd212219, -32'sd564011, -32'sd1327633, -32'sd2803721, -32'sd3508744, -32'sd1168460, 32'sd1854517, 32'sd961129, 32'sd1469888, 32'sd2786718, 32'sd80674, -32'sd890453, 32'sd1536391, 32'sd557135, -32'sd1032191, 32'sd587081, -32'sd369986, -32'sd450248, -32'sd2026422, -32'sd908764, -32'sd1488228, -32'sd566270, -32'sd216086, 32'sd54545, 32'sd0, 32'sd501344, -32'sd1207182, -32'sd379927, 32'sd42545, -32'sd2281064, -32'sd1363758, -32'sd3018792, -32'sd2856748, -32'sd2685358, -32'sd356360, 32'sd2458602, 32'sd1062445, 32'sd1760611, 32'sd747278, 32'sd1396774, 32'sd18379, 32'sd1160863, 32'sd364688, -32'sd1055307, 32'sd877448, -32'sd76638, -32'sd2650868, -32'sd2583144, 32'sd780470, 32'sd694488, 32'sd385892, 32'sd42804, 32'sd37301, -32'sd1130214, -32'sd167739, 32'sd186126, -32'sd995714, -32'sd1462295, -32'sd220349, -32'sd978667, -32'sd2509584, -32'sd2952244, -32'sd1191855, -32'sd1114724, 32'sd1074749, 32'sd3262665, 32'sd2907979, 32'sd1617161, 32'sd2296733, -32'sd439879, -32'sd1073525, 32'sd440813, -32'sd1881716, -32'sd1845726, -32'sd674550, 32'sd1436411, -32'sd1315547, 32'sd136955, -32'sd776408, 32'sd356845, -32'sd148944, -32'sd741624, 32'sd263506, -32'sd586893, -32'sd121786, 32'sd590453, -32'sd445645, -32'sd1915105, -32'sd1901435, -32'sd3056930, -32'sd2695645, -32'sd513473, 32'sd2431501, 32'sd764614, 32'sd1191674, 32'sd1001398, 32'sd1350506, 32'sd1438088, -32'sd1779762, -32'sd619930, -32'sd2053972, -32'sd2457089, -32'sd147202, 32'sd557094, -32'sd2647352, -32'sd899395, -32'sd1721506, 32'sd935136, 32'sd0, 32'sd266351, -32'sd364494, -32'sd670095, -32'sd1827050, -32'sd1171203, -32'sd1290058, -32'sd1629439, -32'sd1621334, -32'sd2013663, -32'sd2136976, -32'sd1071132, 32'sd739812, 32'sd1095606, 32'sd1947125, 32'sd1386593, 32'sd1965205, -32'sd27984, -32'sd1592965, -32'sd163222, -32'sd918512, 32'sd640194, -32'sd147450, 32'sd268047, 32'sd4611, 32'sd249492, 32'sd490598, 32'sd0, 32'sd0, 32'sd0, 32'sd202974, -32'sd819055, -32'sd723047, -32'sd274397, -32'sd1722701, -32'sd1146334, -32'sd1582126, -32'sd1340132, -32'sd1849419, -32'sd1319855, -32'sd1762635, -32'sd617462, 32'sd1851355, -32'sd485249, -32'sd434562, -32'sd1423139, -32'sd1579636, -32'sd792565, -32'sd75078, -32'sd1804426, -32'sd243169, 32'sd626885, -32'sd1126759, -32'sd1193608, -32'sd73548, 32'sd0, 32'sd0, 32'sd0, -32'sd55434, 32'sd222263, -32'sd315487, 32'sd521037, -32'sd1690144, 32'sd467938, -32'sd508134, -32'sd1213401, -32'sd2030675, -32'sd2004821, -32'sd1982777, -32'sd2821580, -32'sd793221, 32'sd38423, -32'sd1966193, -32'sd430166, -32'sd3254277, 32'sd199539, 32'sd862820, -32'sd1420833, -32'sd2195600, -32'sd14496, 32'sd650773, 32'sd588469, 32'sd961689, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1157716, -32'sd93863, -32'sd894955, 32'sd835270, 32'sd1316451, 32'sd1140842, -32'sd573037, -32'sd821341, 32'sd163810, -32'sd748458, -32'sd1866970, -32'sd1931842, -32'sd1432408, -32'sd102970, 32'sd621784, -32'sd544186, -32'sd1790761, 32'sd39966, -32'sd1871514, -32'sd1564201, -32'sd235417, 32'sd335740, 32'sd1017619, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd882131, 32'sd260807, 32'sd1439199, 32'sd1721779, 32'sd156676, -32'sd483849, -32'sd227695, 32'sd1163941, -32'sd1057229, 32'sd439956, -32'sd764334, -32'sd387573, 32'sd698183, 32'sd1139197, -32'sd401572, 32'sd3305138, 32'sd2169661, -32'sd975370, -32'sd746615, 32'sd1279271, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1666424, 32'sd345738, -32'sd32107, -32'sd31609, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1001084, 32'sd661033, -32'sd467424, -32'sd1365566, -32'sd753490, -32'sd1857254, 32'sd677978, -32'sd661307, 32'sd1523000, 32'sd145102, 32'sd1020650, -32'sd561145, 32'sd486231, 32'sd134909, -32'sd39491, 32'sd885523, 32'sd1509880, 32'sd1029538, 32'sd503293, -32'sd153038, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd89823, 32'sd808020, 32'sd1623038, -32'sd675398, -32'sd303470, -32'sd1868467, 32'sd935317, 32'sd698705, 32'sd1085964, -32'sd678984, 32'sd92194, 32'sd540184, -32'sd1204453, 32'sd630445, 32'sd103818, 32'sd595422, -32'sd594640, 32'sd403591, -32'sd1036128, -32'sd1580072, -32'sd991273, 32'sd595126, 32'sd1070792, 32'sd187787, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd826115, 32'sd267874, -32'sd839827, -32'sd1520358, 32'sd679346, -32'sd403540, 32'sd909424, -32'sd895895, 32'sd84583, 32'sd679397, 32'sd1219139, 32'sd474715, 32'sd1378058, 32'sd790398, -32'sd1794533, -32'sd264465, -32'sd1550154, -32'sd698251, 32'sd31126, 32'sd680186, 32'sd1543544, 32'sd541378, -32'sd322407, 32'sd877645, 32'sd36678, 32'sd0, 32'sd0, 32'sd310035, 32'sd903797, -32'sd971144, -32'sd398242, 32'sd120155, -32'sd911581, -32'sd1159213, -32'sd993902, -32'sd941846, -32'sd2885642, 32'sd104173, 32'sd880179, -32'sd450851, -32'sd2029795, -32'sd902241, -32'sd2273445, -32'sd1818278, -32'sd2777076, -32'sd76195, -32'sd591379, 32'sd2298482, 32'sd1542494, 32'sd1718216, 32'sd737632, 32'sd830987, 32'sd748416, 32'sd815834, 32'sd0, 32'sd481664, 32'sd784902, 32'sd431706, -32'sd1468460, -32'sd1140461, 32'sd2081406, 32'sd1061678, -32'sd376354, -32'sd914621, -32'sd1599605, -32'sd2142868, -32'sd146943, -32'sd1161531, 32'sd869176, -32'sd1195046, -32'sd2054551, -32'sd1328320, 32'sd495817, 32'sd72433, -32'sd140011, 32'sd674613, 32'sd2208377, 32'sd2855440, 32'sd1389084, 32'sd1176708, 32'sd183643, 32'sd1046883, 32'sd0, 32'sd1026868, -32'sd148404, -32'sd230360, 32'sd490636, 32'sd1083755, 32'sd101792, -32'sd1719494, 32'sd193111, -32'sd4157288, -32'sd1431706, 32'sd576975, -32'sd326285, -32'sd102139, 32'sd362375, -32'sd976346, -32'sd3381033, -32'sd1460986, 32'sd867165, -32'sd1319885, 32'sd851923, -32'sd434348, 32'sd108612, 32'sd2134402, 32'sd1325256, 32'sd807316, -32'sd1352944, 32'sd118077, 32'sd1024980, -32'sd68497, -32'sd31860, 32'sd401736, 32'sd18650, 32'sd2227643, -32'sd1918930, -32'sd331695, -32'sd376607, -32'sd2693574, -32'sd458696, 32'sd1240737, 32'sd1407092, 32'sd1657297, 32'sd452157, -32'sd1094045, -32'sd2488467, -32'sd412161, -32'sd274888, 32'sd55332, -32'sd2608839, -32'sd3110468, -32'sd299825, -32'sd299874, -32'sd465757, -32'sd637513, 32'sd143296, 32'sd607042, 32'sd1307937, -32'sd840457, -32'sd285959, 32'sd1119868, 32'sd1140763, -32'sd1363034, 32'sd119828, -32'sd740226, -32'sd2735682, -32'sd2574674, -32'sd329710, -32'sd1250647, 32'sd1444836, 32'sd1127961, 32'sd252790, -32'sd3217890, -32'sd3135076, -32'sd2578056, -32'sd593596, -32'sd1655601, -32'sd1338125, -32'sd204896, -32'sd266606, -32'sd784590, 32'sd432511, 32'sd1153611, 32'sd45878, 32'sd609687, -32'sd158409, 32'sd57571, -32'sd1465113, 32'sd903049, -32'sd757830, -32'sd993558, -32'sd949596, -32'sd897564, -32'sd2392082, -32'sd874287, -32'sd3358600, 32'sd1113397, 32'sd876324, 32'sd1847053, -32'sd284152, -32'sd3480267, -32'sd2068220, -32'sd71740, -32'sd130384, 32'sd893013, -32'sd579957, -32'sd1354078, -32'sd5542, -32'sd280503, -32'sd478530, -32'sd1177806, -32'sd99557, -32'sd939862, 32'sd1082743, 32'sd2217389, -32'sd238845, -32'sd1339766, -32'sd1068390, 32'sd468511, -32'sd2590666, -32'sd3665847, -32'sd2255061, 32'sd210511, -32'sd3350297, -32'sd1581273, 32'sd239288, -32'sd1420149, 32'sd1129488, -32'sd1270087, 32'sd570780, 32'sd1920077, 32'sd35804, 32'sd2164400, 32'sd280661, 32'sd579360, 32'sd1549827, 32'sd274883, 32'sd897931, -32'sd1163943, -32'sd1069781, 32'sd505230, 32'sd1678385, 32'sd1211761, -32'sd232787, 32'sd201836, 32'sd106557, -32'sd1363932, -32'sd2711916, -32'sd1327693, 32'sd42997, 32'sd522960, -32'sd677749, -32'sd976410, 32'sd1304942, 32'sd1254665, 32'sd860070, -32'sd530189, 32'sd2938126, 32'sd1945725, 32'sd3487461, 32'sd2307783, 32'sd274141, -32'sd586856, 32'sd1724963, 32'sd2917729, 32'sd1643620, -32'sd563077, 32'sd1295010, -32'sd1896562, -32'sd4524, 32'sd594689, -32'sd1171724, 32'sd259888, 32'sd416261, 32'sd390943, -32'sd2501532, 32'sd94884, 32'sd1053769, 32'sd1527589, -32'sd81120, 32'sd273732, -32'sd426389, 32'sd2340375, 32'sd4075578, 32'sd1277237, 32'sd26974, 32'sd1770570, 32'sd1619888, 32'sd2777902, 32'sd1275035, 32'sd1931608, 32'sd2547912, 32'sd1039981, 32'sd1339509, -32'sd646566, 32'sd1333726, 32'sd530440, 32'sd365394, -32'sd327503, 32'sd1338760, -32'sd130376, -32'sd420808, -32'sd1407732, -32'sd175206, -32'sd721795, 32'sd556598, 32'sd846678, 32'sd1785836, 32'sd2930971, 32'sd2239477, 32'sd3267794, 32'sd2323165, 32'sd544348, -32'sd235370, 32'sd982368, -32'sd665648, 32'sd1396277, 32'sd798479, 32'sd1614209, -32'sd216035, 32'sd294106, -32'sd606769, -32'sd211158, -32'sd395821, -32'sd81695, 32'sd1260626, 32'sd232972, -32'sd1324377, 32'sd1471743, 32'sd442429, -32'sd79833, -32'sd3019197, 32'sd62479, -32'sd25318, 32'sd2581570, 32'sd2566095, 32'sd2015468, 32'sd309345, 32'sd2175603, 32'sd719118, 32'sd487883, 32'sd1476977, 32'sd1276445, -32'sd54640, 32'sd719595, 32'sd1803152, 32'sd356684, -32'sd1384717, -32'sd2729323, -32'sd904293, -32'sd2354855, -32'sd442717, -32'sd400642, -32'sd51289, 32'sd944380, -32'sd759092, 32'sd165102, 32'sd942832, -32'sd937066, -32'sd1423868, 32'sd483292, 32'sd1993679, 32'sd1244108, 32'sd1176802, 32'sd525832, 32'sd1151983, -32'sd619333, 32'sd2251790, 32'sd1362680, -32'sd168392, 32'sd875313, -32'sd425576, -32'sd328163, -32'sd2450234, -32'sd111875, -32'sd1315402, -32'sd1379369, -32'sd576504, -32'sd156012, -32'sd1312865, -32'sd414128, 32'sd1109761, 32'sd600551, -32'sd264743, -32'sd72110, 32'sd1040908, -32'sd272745, -32'sd1549532, -32'sd1930611, 32'sd1017630, -32'sd665514, 32'sd563608, -32'sd939218, -32'sd44342, 32'sd524299, 32'sd346937, 32'sd438546, -32'sd1820119, 32'sd1470512, 32'sd121509, -32'sd1781151, -32'sd1305240, -32'sd1728893, -32'sd1515985, -32'sd2404388, -32'sd1703307, -32'sd1471890, 32'sd173679, 32'sd738394, 32'sd0, -32'sd34653, -32'sd1256878, -32'sd191455, 32'sd2029754, -32'sd1133822, -32'sd630221, -32'sd2015185, -32'sd161401, -32'sd1149340, 32'sd1177082, -32'sd212753, 32'sd932484, -32'sd455418, 32'sd607714, -32'sd913636, -32'sd1166215, -32'sd38677, -32'sd211758, -32'sd358294, -32'sd316689, -32'sd1946751, -32'sd1500092, -32'sd1402402, -32'sd1625756, -32'sd21965, 32'sd395241, -32'sd1579310, -32'sd718064, 32'sd614312, -32'sd1912066, -32'sd411005, 32'sd76535, -32'sd1358557, -32'sd1235219, -32'sd595945, -32'sd515738, -32'sd769993, 32'sd2010345, 32'sd2594766, 32'sd1472360, -32'sd1821079, -32'sd1587100, -32'sd1690435, -32'sd1002404, 32'sd996471, -32'sd1510730, -32'sd958640, -32'sd656110, -32'sd394452, -32'sd3384185, -32'sd3011714, -32'sd2551037, -32'sd737739, 32'sd1350556, 32'sd454754, 32'sd646833, 32'sd305932, -32'sd1310479, -32'sd2290302, -32'sd1954451, 32'sd1246034, -32'sd1407252, 32'sd530122, -32'sd992764, 32'sd538885, 32'sd1988027, 32'sd984980, 32'sd644781, -32'sd112702, -32'sd581008, -32'sd655154, -32'sd446082, 32'sd446932, 32'sd483836, -32'sd2160552, -32'sd2055592, -32'sd1437894, -32'sd2977596, -32'sd1625591, -32'sd1479451, -32'sd747602, 32'sd974230, -32'sd1422267, 32'sd0, -32'sd31411, 32'sd1500939, -32'sd2905075, -32'sd1063922, -32'sd2585739, -32'sd467163, -32'sd1245945, -32'sd1316190, 32'sd99245, 32'sd777496, 32'sd603654, -32'sd974480, 32'sd475859, -32'sd1113334, 32'sd1242282, -32'sd421069, 32'sd42802, -32'sd889814, -32'sd1090704, -32'sd2351397, -32'sd3336684, -32'sd1735054, -32'sd2941490, -32'sd1996847, 32'sd1013839, 32'sd1384657, 32'sd1055049, 32'sd1491639, -32'sd68158, 32'sd757270, -32'sd196530, -32'sd1410772, -32'sd668022, -32'sd1609885, 32'sd1158882, -32'sd900631, 32'sd1678391, -32'sd1704209, -32'sd1353240, -32'sd47385, 32'sd147332, -32'sd1522174, 32'sd23605, -32'sd1258472, -32'sd610285, -32'sd1723008, -32'sd3273005, -32'sd1287168, -32'sd1784689, -32'sd294358, -32'sd1045499, -32'sd143936, 32'sd757256, 32'sd595308, 32'sd1158473, -32'sd232515, 32'sd892321, 32'sd863662, 32'sd61083, -32'sd1572943, -32'sd1440715, 32'sd560776, -32'sd265112, 32'sd1149340, 32'sd931938, 32'sd540595, 32'sd311623, 32'sd878228, 32'sd495377, 32'sd786280, -32'sd2235880, -32'sd4146548, -32'sd4293848, -32'sd2923819, -32'sd873771, -32'sd2474486, -32'sd1477225, 32'sd463220, -32'sd1845195, -32'sd1407798, -32'sd399797, 32'sd156968, 32'sd884438, 32'sd0, -32'sd58550, 32'sd17783, -32'sd793443, -32'sd1645793, -32'sd694292, -32'sd1127847, -32'sd910737, 32'sd2885036, 32'sd64683, 32'sd159636, 32'sd82545, -32'sd957140, -32'sd1836088, -32'sd1290282, -32'sd3815755, -32'sd420158, -32'sd2757962, -32'sd1187776, -32'sd885000, -32'sd2071679, -32'sd1698486, -32'sd331135, 32'sd335336, -32'sd529913, 32'sd527584, -32'sd1252498, 32'sd0, 32'sd0, 32'sd0, -32'sd68753, -32'sd469619, 32'sd1120489, 32'sd427376, -32'sd610953, -32'sd365582, 32'sd1009309, 32'sd247386, -32'sd160780, 32'sd473600, -32'sd367883, -32'sd323608, 32'sd1078683, -32'sd1159672, 32'sd2166937, -32'sd1444151, -32'sd2541593, -32'sd461855, -32'sd1137465, 32'sd817635, 32'sd84728, -32'sd498627, -32'sd790570, -32'sd128803, 32'sd96611, 32'sd0, 32'sd0, 32'sd0, 32'sd558651, -32'sd1873997, 32'sd131865, -32'sd781178, -32'sd82683, 32'sd802294, 32'sd366066, 32'sd57789, -32'sd830188, 32'sd705911, -32'sd1973386, -32'sd617303, -32'sd1264389, -32'sd423842, -32'sd943511, -32'sd2571225, 32'sd273291, 32'sd841381, 32'sd502455, 32'sd8496, -32'sd2110240, -32'sd603248, -32'sd729689, -32'sd355168, -32'sd10972, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1041513, 32'sd1437330, -32'sd776651, -32'sd79449, -32'sd108323, 32'sd196760, -32'sd2043402, -32'sd1168841, 32'sd3161623, -32'sd198226, 32'sd1049942, 32'sd474322, -32'sd452277, -32'sd297115, -32'sd1314596, 32'sd868552, -32'sd31966, 32'sd748620, -32'sd665394, 32'sd313602, 32'sd493626, -32'sd495988, 32'sd68834, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd288284, 32'sd355756, -32'sd389893, -32'sd399110, -32'sd1049950, 32'sd203967, 32'sd409643, 32'sd658856, -32'sd767137, 32'sd1149721, 32'sd790542, 32'sd1111650, 32'sd211073, 32'sd208337, 32'sd935236, -32'sd1177761, -32'sd1342130, -32'sd815632, -32'sd278391, -32'sd255, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1213472, -32'sd1335802, 32'sd373747, -32'sd500499, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd188958, -32'sd640787, 32'sd766915, -32'sd1582915, -32'sd606791, 32'sd308875, 32'sd1295785, 32'sd65030, -32'sd728441, 32'sd496422, -32'sd451500, 32'sd240796, -32'sd232830, 32'sd218810, 32'sd331139, 32'sd768242, 32'sd944190, 32'sd1043895, 32'sd772522, 32'sd177836, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd758504, 32'sd797016, 32'sd172632, 32'sd26341, 32'sd46744, -32'sd335718, -32'sd1065088, -32'sd622532, 32'sd1332009, 32'sd1393602, -32'sd1345807, 32'sd296627, -32'sd1120038, 32'sd23678, -32'sd444262, 32'sd3054200, 32'sd1112091, 32'sd1749781, -32'sd78993, 32'sd1617952, 32'sd460929, -32'sd151733, 32'sd1016221, 32'sd562740, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd934718, 32'sd85989, 32'sd860795, -32'sd270153, 32'sd897767, 32'sd1074630, 32'sd42052, 32'sd2007660, 32'sd235532, -32'sd2116199, -32'sd1532626, -32'sd239507, -32'sd1174905, -32'sd1688002, -32'sd1338714, 32'sd2661836, 32'sd1306774, 32'sd2678866, -32'sd487684, -32'sd713862, -32'sd749840, -32'sd30160, 32'sd86754, -32'sd307382, -32'sd952412, 32'sd0, 32'sd0, 32'sd684660, 32'sd1286285, -32'sd602256, -32'sd1615466, 32'sd651060, -32'sd1215453, -32'sd352168, 32'sd584123, 32'sd207082, -32'sd1897172, 32'sd168799, 32'sd1057687, -32'sd287389, -32'sd1894239, -32'sd1627337, 32'sd339527, 32'sd2895176, 32'sd1865275, 32'sd1221215, -32'sd1724003, -32'sd2829888, -32'sd2335488, -32'sd1994488, 32'sd588474, 32'sd294579, -32'sd945290, -32'sd398485, 32'sd0, -32'sd170068, 32'sd1466675, -32'sd1101398, 32'sd202026, -32'sd898109, -32'sd2123416, -32'sd758814, -32'sd2470964, -32'sd2952003, -32'sd2653206, -32'sd1699443, -32'sd2180873, -32'sd636144, 32'sd636678, 32'sd2056025, 32'sd2280459, 32'sd1087574, 32'sd748206, 32'sd1024356, -32'sd144194, -32'sd2273037, -32'sd2227825, -32'sd1076304, 32'sd77968, 32'sd129241, 32'sd784594, 32'sd1021244, 32'sd0, -32'sd181160, 32'sd630417, -32'sd510151, -32'sd860498, -32'sd236717, -32'sd1264994, -32'sd1503641, -32'sd1002779, -32'sd4334786, -32'sd2919795, 32'sd312060, -32'sd184595, 32'sd968922, 32'sd2978319, 32'sd1420542, 32'sd967508, -32'sd1106648, -32'sd536758, -32'sd317215, -32'sd2291752, -32'sd2114827, 32'sd7488, 32'sd222866, -32'sd1646843, -32'sd819626, -32'sd164327, -32'sd249399, 32'sd268682, -32'sd114270, -32'sd750804, -32'sd276204, -32'sd515002, -32'sd865454, -32'sd3581924, -32'sd3905576, -32'sd3170436, -32'sd2815075, -32'sd756134, 32'sd2362305, 32'sd2427923, 32'sd2814476, 32'sd831350, -32'sd90875, -32'sd634383, -32'sd1409171, -32'sd1932950, -32'sd2359378, -32'sd2164605, -32'sd1581890, 32'sd2092236, -32'sd1437930, -32'sd320271, -32'sd571563, 32'sd1691334, 32'sd658547, 32'sd167637, -32'sd651795, -32'sd146711, -32'sd356163, -32'sd1743372, -32'sd1852167, -32'sd3583332, -32'sd3270908, -32'sd2425578, -32'sd2983946, -32'sd1034331, 32'sd1330596, 32'sd3430661, 32'sd929618, -32'sd1298386, -32'sd1987427, -32'sd2146162, -32'sd1312167, -32'sd1581099, -32'sd37039, -32'sd1833292, -32'sd64993, 32'sd350713, 32'sd571805, 32'sd1634915, 32'sd3696978, 32'sd423491, 32'sd1454136, -32'sd167928, -32'sd1148491, 32'sd1646622, -32'sd767739, -32'sd2384930, -32'sd3543734, -32'sd633937, -32'sd2639280, 32'sd36846, -32'sd675127, 32'sd736843, 32'sd3351289, 32'sd2161783, 32'sd934902, -32'sd1443708, -32'sd1737977, 32'sd41851, -32'sd168782, -32'sd1876414, 32'sd1740700, -32'sd1424991, 32'sd85952, 32'sd582670, 32'sd1137358, 32'sd1103454, 32'sd620486, 32'sd1068166, 32'sd1277087, -32'sd1117536, -32'sd186267, 32'sd1632987, 32'sd261660, -32'sd123741, -32'sd1650391, -32'sd2497098, -32'sd1397952, 32'sd1180443, -32'sd1316323, -32'sd789679, -32'sd710358, -32'sd280919, -32'sd60773, 32'sd231667, 32'sd326327, -32'sd1620366, -32'sd271871, 32'sd944743, 32'sd2527589, 32'sd1083745, 32'sd2900701, 32'sd346956, 32'sd1762074, 32'sd987713, 32'sd1431133, 32'sd1299463, -32'sd1272410, -32'sd179524, -32'sd43517, -32'sd12506, -32'sd846575, -32'sd694029, -32'sd1069192, -32'sd995375, -32'sd595958, -32'sd335454, -32'sd272352, -32'sd458838, -32'sd903444, -32'sd820416, 32'sd1298364, 32'sd346404, 32'sd72295, 32'sd930444, 32'sd306500, 32'sd247660, 32'sd558127, 32'sd308000, 32'sd241279, 32'sd869600, 32'sd478861, 32'sd1207751, 32'sd278411, -32'sd441531, 32'sd790604, 32'sd984768, 32'sd580313, 32'sd808803, -32'sd619675, -32'sd1794414, 32'sd33996, 32'sd546983, 32'sd930112, -32'sd351316, 32'sd424610, 32'sd860887, 32'sd3208586, 32'sd1847625, 32'sd741813, 32'sd1481157, 32'sd140083, -32'sd939153, 32'sd55325, -32'sd1930099, 32'sd562501, 32'sd1145445, 32'sd441845, 32'sd1412519, -32'sd205904, -32'sd590059, 32'sd1245155, 32'sd592461, -32'sd446146, -32'sd63053, -32'sd521852, -32'sd1422117, 32'sd938467, -32'sd1161549, -32'sd954687, -32'sd969836, 32'sd79461, 32'sd545566, 32'sd2720719, -32'sd42171, 32'sd1095181, 32'sd2502394, 32'sd134814, -32'sd77915, -32'sd1146936, -32'sd1699996, -32'sd749515, -32'sd3338208, 32'sd744168, -32'sd1784285, -32'sd1098939, 32'sd484131, -32'sd1196076, -32'sd1902142, -32'sd1127416, -32'sd3545, 32'sd640745, 32'sd2016450, 32'sd224205, -32'sd495007, 32'sd1220087, 32'sd259775, -32'sd1942978, -32'sd1972734, -32'sd248220, 32'sd380860, 32'sd2366503, 32'sd1189242, 32'sd1203924, 32'sd2279692, -32'sd601520, -32'sd2153949, -32'sd1068879, 32'sd265671, 32'sd641860, -32'sd2749049, -32'sd2942148, -32'sd1644599, 32'sd555498, 32'sd2975415, -32'sd187264, -32'sd131300, -32'sd909027, -32'sd352652, 32'sd1018296, 32'sd839982, 32'sd862386, -32'sd397528, 32'sd2268608, 32'sd1287638, 32'sd809478, 32'sd238919, 32'sd495523, 32'sd1378629, 32'sd2090449, 32'sd383834, 32'sd543458, -32'sd636200, -32'sd1118335, -32'sd1039056, 32'sd1355755, 32'sd1591939, -32'sd1420384, -32'sd1849967, -32'sd1805228, 32'sd346281, 32'sd1757681, -32'sd364968, -32'sd466162, -32'sd1173580, -32'sd825181, -32'sd189969, 32'sd249779, -32'sd25125, -32'sd1126370, 32'sd5696, 32'sd204188, 32'sd657186, -32'sd438235, -32'sd1561861, -32'sd2210600, 32'sd1139561, -32'sd516803, 32'sd1795820, -32'sd232074, 32'sd952825, -32'sd975142, 32'sd1124862, 32'sd673799, 32'sd1198060, -32'sd2500281, -32'sd2362757, -32'sd430447, -32'sd517483, 32'sd303303, -32'sd1172911, -32'sd622462, -32'sd592445, -32'sd336561, 32'sd985087, 32'sd139808, 32'sd0, 32'sd1380429, 32'sd523558, 32'sd64244, -32'sd182822, 32'sd217475, 32'sd810728, -32'sd935023, -32'sd921952, -32'sd2616805, 32'sd1443631, 32'sd1233525, -32'sd589712, -32'sd1311907, -32'sd830580, 32'sd2166793, 32'sd172705, -32'sd75933, -32'sd3174875, -32'sd1851000, 32'sd895301, 32'sd365815, 32'sd226771, -32'sd1745829, -32'sd992121, -32'sd763908, 32'sd2246198, -32'sd1031204, -32'sd546273, -32'sd168654, 32'sd898739, -32'sd1022882, 32'sd171156, -32'sd895220, 32'sd224525, 32'sd97726, -32'sd1181383, -32'sd1896916, -32'sd1799706, -32'sd2715222, 32'sd424796, -32'sd1001384, 32'sd674385, 32'sd2566770, 32'sd602854, -32'sd2638493, -32'sd2041556, -32'sd2264742, -32'sd280922, -32'sd459849, 32'sd139132, -32'sd251029, -32'sd525835, 32'sd356620, -32'sd309901, 32'sd1135097, 32'sd76105, 32'sd599028, 32'sd946780, -32'sd283420, -32'sd441174, 32'sd518277, -32'sd714619, -32'sd90888, -32'sd435520, -32'sd1920612, -32'sd496688, -32'sd340347, -32'sd672881, -32'sd622794, 32'sd456711, 32'sd2799206, -32'sd922918, -32'sd1030834, 32'sd1110175, -32'sd1655058, 32'sd181135, 32'sd614866, -32'sd1104693, 32'sd1126928, -32'sd186936, -32'sd827017, 32'sd193472, -32'sd478585, 32'sd0, 32'sd279277, -32'sd588469, 32'sd544191, -32'sd81559, 32'sd1579308, 32'sd1026977, -32'sd1555328, -32'sd2877655, -32'sd1121701, 32'sd60397, 32'sd607089, 32'sd1261030, 32'sd414963, -32'sd728726, 32'sd1241214, 32'sd2481872, 32'sd1266420, 32'sd2197167, 32'sd616167, -32'sd593706, 32'sd29040, 32'sd752565, -32'sd585121, 32'sd297072, -32'sd391428, 32'sd637062, -32'sd430034, 32'sd1347084, -32'sd292152, -32'sd684806, 32'sd1564674, -32'sd181610, -32'sd1653245, -32'sd1376873, -32'sd610277, -32'sd245880, 32'sd1896237, -32'sd336339, 32'sd1412087, 32'sd1359151, 32'sd1694797, 32'sd652694, 32'sd1667936, 32'sd534549, 32'sd1814418, -32'sd322280, -32'sd822408, 32'sd48580, -32'sd380894, -32'sd61832, 32'sd1403437, 32'sd939488, 32'sd591338, 32'sd279388, -32'sd247335, 32'sd1066231, 32'sd1185948, -32'sd798658, 32'sd1946316, 32'sd130194, -32'sd2883875, -32'sd3389602, -32'sd1579147, -32'sd802191, -32'sd97220, 32'sd981542, -32'sd624055, 32'sd1461946, 32'sd976732, 32'sd249092, -32'sd166138, 32'sd1374287, 32'sd2108199, 32'sd2122557, 32'sd217766, -32'sd954578, 32'sd411671, 32'sd779326, 32'sd1351812, -32'sd1077100, -32'sd1138789, 32'sd734773, 32'sd83036, 32'sd0, 32'sd713606, -32'sd591808, 32'sd1588726, 32'sd928008, -32'sd865749, -32'sd1792316, -32'sd2331838, 32'sd740905, -32'sd1050247, 32'sd152919, -32'sd575071, 32'sd705607, 32'sd2047038, 32'sd916203, -32'sd581686, 32'sd1767446, 32'sd958210, -32'sd258728, -32'sd1273711, 32'sd291006, 32'sd643227, 32'sd634714, 32'sd748794, -32'sd1267931, 32'sd1042387, 32'sd1634667, 32'sd0, 32'sd0, 32'sd0, -32'sd448962, 32'sd575562, 32'sd532227, -32'sd711961, -32'sd1393985, -32'sd3984129, -32'sd3390627, -32'sd1872090, 32'sd629172, 32'sd660131, 32'sd449972, -32'sd1889504, -32'sd613369, 32'sd122872, 32'sd2068661, -32'sd825640, 32'sd304713, 32'sd361447, 32'sd1165772, -32'sd316679, -32'sd48424, -32'sd740154, -32'sd347115, 32'sd530571, 32'sd511548, 32'sd0, 32'sd0, 32'sd0, -32'sd628361, 32'sd1219113, -32'sd590336, -32'sd738671, -32'sd2276601, -32'sd2961477, -32'sd2150945, -32'sd2207282, -32'sd950428, -32'sd445310, 32'sd526392, 32'sd122308, -32'sd774189, 32'sd509148, 32'sd591389, 32'sd1937275, -32'sd265710, -32'sd685924, 32'sd2335115, 32'sd1131163, -32'sd592699, -32'sd91504, 32'sd387129, -32'sd276462, 32'sd278624, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd824486, -32'sd212843, -32'sd520819, -32'sd996600, 32'sd1028663, 32'sd33700, -32'sd419663, 32'sd604217, 32'sd515982, 32'sd710095, 32'sd1113194, 32'sd239282, 32'sd1170624, 32'sd619500, 32'sd1214103, -32'sd32929, 32'sd37027, 32'sd1182641, -32'sd1126181, -32'sd1111504, 32'sd484771, -32'sd579937, 32'sd690738, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd478138, 32'sd1086924, -32'sd4218, 32'sd641940, -32'sd1148253, 32'sd618098, 32'sd443478, -32'sd797215, -32'sd6955, 32'sd735126, -32'sd898392, 32'sd1185037, 32'sd294465, -32'sd522281, 32'sd1210446, -32'sd149876, -32'sd197928, -32'sd155380, 32'sd1252566, 32'sd388751, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1657394, 32'sd1464868, 32'sd1619951, 32'sd1950900, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd587292, 32'sd1778713, 32'sd1053199, 32'sd554889, 32'sd1155994, -32'sd513740, 32'sd2239809, 32'sd2330877, 32'sd1976824, 32'sd1096781, -32'sd29268, -32'sd815909, 32'sd66621, -32'sd1514137, -32'sd726559, -32'sd144535, -32'sd894330, -32'sd176608, -32'sd60667, 32'sd29552, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd33546, -32'sd219759, -32'sd425115, 32'sd1146861, 32'sd1296818, 32'sd2099545, 32'sd991347, 32'sd980574, -32'sd249615, 32'sd54297, 32'sd221703, -32'sd271968, -32'sd23067, 32'sd195657, -32'sd576705, -32'sd1033620, 32'sd481990, 32'sd788650, -32'sd314483, 32'sd1616404, 32'sd2616265, 32'sd780196, 32'sd446301, -32'sd303445, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd681138, -32'sd318165, 32'sd504950, 32'sd1124915, 32'sd1168813, 32'sd114879, 32'sd1453791, 32'sd35215, -32'sd1724583, 32'sd5470, -32'sd485996, -32'sd1365693, -32'sd459024, 32'sd104481, -32'sd1398322, 32'sd663482, 32'sd710441, 32'sd184777, 32'sd28220, 32'sd1757928, -32'sd491719, 32'sd2316279, -32'sd335981, -32'sd95592, -32'sd2337227, 32'sd0, 32'sd0, 32'sd1212435, 32'sd917008, -32'sd460535, -32'sd1536755, -32'sd1857639, 32'sd1188771, 32'sd104242, -32'sd1649947, 32'sd426002, -32'sd414060, -32'sd122933, -32'sd35403, 32'sd2154824, 32'sd1311271, 32'sd1082363, -32'sd684017, 32'sd1250136, 32'sd1561677, 32'sd1724938, 32'sd1479559, 32'sd2829106, 32'sd1241357, 32'sd164875, -32'sd1405600, -32'sd438091, -32'sd1420251, 32'sd1202965, 32'sd0, 32'sd636584, -32'sd637273, 32'sd1110457, -32'sd269974, -32'sd301433, 32'sd435598, -32'sd1137199, 32'sd984980, 32'sd1232020, 32'sd2015490, -32'sd260842, -32'sd1830905, -32'sd2513322, -32'sd1277107, -32'sd1367432, -32'sd577627, -32'sd188894, -32'sd989249, 32'sd646244, 32'sd1286305, 32'sd1235258, 32'sd3406136, 32'sd1092655, 32'sd406929, 32'sd982817, -32'sd2507664, 32'sd327369, 32'sd0, 32'sd12143, -32'sd949850, -32'sd115692, -32'sd239580, -32'sd902909, -32'sd749263, -32'sd403880, 32'sd604864, 32'sd1147503, 32'sd5631, -32'sd835630, -32'sd1630610, -32'sd203134, -32'sd1880457, -32'sd1161510, -32'sd2558418, 32'sd808514, -32'sd364807, -32'sd510805, 32'sd1260823, -32'sd423426, 32'sd770522, 32'sd541905, 32'sd2361154, -32'sd735560, -32'sd479575, -32'sd961616, 32'sd480952, 32'sd257938, -32'sd395369, -32'sd3, -32'sd84462, -32'sd2312013, -32'sd2280793, -32'sd2444904, 32'sd650911, 32'sd1296664, -32'sd1476302, -32'sd3082998, -32'sd3008096, -32'sd1225129, 32'sd913853, 32'sd915891, -32'sd698115, 32'sd509721, -32'sd1401723, 32'sd906426, 32'sd537965, -32'sd206015, 32'sd156953, 32'sd816157, 32'sd326663, 32'sd392184, 32'sd726529, -32'sd564808, 32'sd968579, 32'sd44337, -32'sd1049775, 32'sd935914, -32'sd1188569, -32'sd209448, -32'sd723762, -32'sd388890, -32'sd925693, -32'sd407742, -32'sd1103106, 32'sd173822, -32'sd2986390, -32'sd669766, 32'sd2574785, -32'sd421906, -32'sd2286751, -32'sd1779519, 32'sd14214, 32'sd10360, -32'sd21142, 32'sd394925, 32'sd564163, 32'sd1858047, 32'sd573178, -32'sd906897, -32'sd235941, -32'sd971467, 32'sd1806464, -32'sd634302, 32'sd300923, 32'sd1779589, -32'sd934162, -32'sd285440, 32'sd591320, 32'sd1126570, -32'sd211232, 32'sd1550798, 32'sd801805, -32'sd118334, -32'sd2133359, -32'sd1576859, -32'sd1051873, 32'sd644413, 32'sd330154, -32'sd974452, -32'sd1390528, 32'sd1827173, 32'sd336552, 32'sd974073, 32'sd1330476, 32'sd2178732, -32'sd688571, 32'sd309207, -32'sd1019612, -32'sd940459, -32'sd108692, 32'sd1041060, -32'sd422995, -32'sd1061396, 32'sd284240, 32'sd1074980, -32'sd684598, 32'sd2493886, 32'sd1693562, 32'sd1965893, 32'sd1067759, 32'sd1108516, -32'sd2161653, -32'sd439814, -32'sd1559325, 32'sd522807, -32'sd1807114, -32'sd1864025, -32'sd58285, -32'sd1505497, -32'sd214880, -32'sd1282092, -32'sd458374, -32'sd385342, 32'sd404885, -32'sd1586104, -32'sd82198, -32'sd268763, 32'sd1126724, 32'sd176774, -32'sd967854, -32'sd307920, 32'sd611276, 32'sd1465918, 32'sd1223429, 32'sd1228836, 32'sd2636880, 32'sd3192766, 32'sd2622261, 32'sd1449428, 32'sd859321, -32'sd1433101, 32'sd167862, 32'sd588053, -32'sd1980307, -32'sd1769987, -32'sd1286176, -32'sd1782386, -32'sd619154, 32'sd800578, -32'sd538632, -32'sd835434, -32'sd172637, -32'sd548737, 32'sd1770226, 32'sd491820, 32'sd703540, 32'sd535566, 32'sd335536, 32'sd1465391, 32'sd653608, 32'sd1223871, -32'sd1136916, 32'sd1663773, 32'sd1296043, 32'sd2678006, 32'sd2755614, 32'sd1237963, 32'sd1325832, -32'sd2179464, -32'sd174073, 32'sd169846, 32'sd466542, -32'sd677113, -32'sd2614920, -32'sd276803, 32'sd205404, -32'sd481339, -32'sd2287576, -32'sd1119280, 32'sd1025678, -32'sd240363, -32'sd211769, 32'sd1339214, 32'sd994804, 32'sd263005, 32'sd702340, 32'sd1185639, 32'sd483166, 32'sd817794, -32'sd1105726, 32'sd490650, 32'sd1705757, 32'sd2173360, 32'sd895342, 32'sd1808, 32'sd783630, -32'sd2051687, 32'sd551863, 32'sd2006247, -32'sd1119627, -32'sd1160730, 32'sd797301, -32'sd1946917, -32'sd350281, -32'sd2314971, -32'sd86781, 32'sd805669, -32'sd2179942, 32'sd1316560, 32'sd823642, -32'sd815877, -32'sd552005, 32'sd1754199, -32'sd797622, -32'sd311817, -32'sd1291141, 32'sd899458, 32'sd65434, 32'sd867858, -32'sd435474, 32'sd954376, 32'sd8449, 32'sd2418434, 32'sd89013, -32'sd389645, 32'sd596658, -32'sd1857234, -32'sd780318, -32'sd1661007, -32'sd648627, -32'sd1770234, -32'sd486491, 32'sd196417, -32'sd477703, -32'sd959230, -32'sd798115, -32'sd385493, 32'sd1052549, -32'sd1044460, 32'sd632921, 32'sd396015, 32'sd931035, -32'sd2429993, -32'sd116163, 32'sd158581, 32'sd1359640, 32'sd1994211, 32'sd1195273, 32'sd168502, -32'sd83361, 32'sd1696817, 32'sd1077739, -32'sd741531, 32'sd960406, -32'sd1665001, -32'sd634756, -32'sd2411603, -32'sd580863, 32'sd27917, 32'sd135763, -32'sd1267015, -32'sd1670869, -32'sd1525367, -32'sd437737, 32'sd104530, -32'sd1115729, -32'sd370749, 32'sd178442, 32'sd109109, 32'sd25692, -32'sd1516990, -32'sd1365811, -32'sd1017781, -32'sd784401, -32'sd278792, 32'sd1336219, 32'sd1332832, 32'sd435097, 32'sd1568713, -32'sd468779, -32'sd804666, 32'sd292599, 32'sd4380, 32'sd562159, 32'sd1286858, -32'sd439565, 32'sd621873, 32'sd220962, 32'sd218039, -32'sd65906, 32'sd883116, 32'sd957399, 32'sd1104468, -32'sd445663, -32'sd143843, 32'sd0, 32'sd913900, -32'sd1384766, 32'sd245184, -32'sd655063, -32'sd1839512, 32'sd1188705, 32'sd932991, 32'sd1334147, -32'sd1097863, 32'sd595693, -32'sd790821, -32'sd40474, 32'sd53839, 32'sd1346150, -32'sd170899, 32'sd705888, 32'sd1174370, 32'sd1510089, -32'sd68107, 32'sd1361519, -32'sd347887, -32'sd268926, -32'sd896804, -32'sd324664, -32'sd531948, -32'sd854729, 32'sd1745323, -32'sd380521, -32'sd513337, -32'sd99482, -32'sd1380694, -32'sd423963, -32'sd922262, -32'sd297794, 32'sd2311299, 32'sd1639534, 32'sd1722876, 32'sd861754, -32'sd1898468, 32'sd1385382, 32'sd184242, 32'sd2110591, 32'sd3183979, 32'sd599873, -32'sd1125975, 32'sd691157, 32'sd1274859, -32'sd71391, -32'sd1401332, 32'sd260458, -32'sd660606, -32'sd316900, 32'sd666675, 32'sd324090, -32'sd388836, -32'sd65118, 32'sd245195, -32'sd1010592, 32'sd666963, -32'sd1819487, -32'sd2171685, 32'sd601977, 32'sd531737, 32'sd1025306, 32'sd437566, 32'sd840882, -32'sd1332778, -32'sd371441, 32'sd2762743, 32'sd1285195, 32'sd1350740, 32'sd57003, -32'sd19577, -32'sd1193307, -32'sd1003264, -32'sd173109, 32'sd432254, 32'sd930457, 32'sd299843, -32'sd1199988, -32'sd370199, 32'sd159522, -32'sd455571, 32'sd0, 32'sd104518, -32'sd1372975, -32'sd394998, -32'sd1593714, -32'sd1596907, -32'sd837437, -32'sd121393, -32'sd470957, 32'sd28073, -32'sd1275995, -32'sd867121, 32'sd1183467, -32'sd92259, 32'sd1791069, 32'sd2052305, -32'sd1137063, -32'sd702204, -32'sd649281, -32'sd403987, -32'sd564836, 32'sd796757, 32'sd1083621, -32'sd1238389, 32'sd198495, 32'sd193445, 32'sd2263040, 32'sd2443182, -32'sd518360, -32'sd585669, 32'sd629206, -32'sd1416923, -32'sd763236, -32'sd1985294, -32'sd544789, -32'sd1255965, -32'sd781927, -32'sd453537, -32'sd824010, 32'sd595584, 32'sd1741918, 32'sd1279486, 32'sd423465, 32'sd428947, 32'sd1015097, 32'sd1047971, -32'sd1254742, 32'sd269995, 32'sd1551074, 32'sd1025826, -32'sd545339, 32'sd1083204, -32'sd1503546, 32'sd1093155, -32'sd204642, -32'sd314901, 32'sd573149, 32'sd6117, -32'sd1174066, -32'sd1007773, -32'sd642014, -32'sd1176397, -32'sd121821, -32'sd1886438, -32'sd1187764, -32'sd1359601, -32'sd1221771, -32'sd448006, 32'sd1693433, 32'sd2843775, 32'sd64806, 32'sd1972389, 32'sd2598411, 32'sd1727548, 32'sd1817595, 32'sd2131115, 32'sd89959, 32'sd1204363, 32'sd482698, -32'sd2095834, -32'sd2181273, -32'sd1765213, 32'sd1334732, 32'sd119763, 32'sd0, -32'sd290859, -32'sd864124, 32'sd383712, 32'sd912953, 32'sd209369, 32'sd139394, 32'sd932580, -32'sd328795, -32'sd1815807, 32'sd247226, -32'sd815418, 32'sd695850, -32'sd537676, 32'sd1787719, -32'sd1263060, 32'sd653288, 32'sd1027434, 32'sd2230068, 32'sd1327248, -32'sd376288, 32'sd113349, -32'sd1120900, -32'sd1151497, -32'sd39480, 32'sd681728, -32'sd1027675, 32'sd0, 32'sd0, 32'sd0, -32'sd579350, -32'sd414009, 32'sd1382507, 32'sd768616, 32'sd576552, 32'sd668690, 32'sd968636, 32'sd237703, -32'sd186883, -32'sd2079211, -32'sd2491559, -32'sd2564717, -32'sd1002202, -32'sd128530, 32'sd443206, 32'sd440629, -32'sd78152, 32'sd34655, -32'sd1239156, -32'sd1704139, -32'sd1930731, -32'sd1368028, -32'sd308959, 32'sd646203, -32'sd357604, 32'sd0, 32'sd0, 32'sd0, 32'sd1243927, 32'sd573399, -32'sd704621, -32'sd809586, 32'sd716413, 32'sd610925, -32'sd1513621, -32'sd316848, -32'sd1355816, -32'sd1295374, -32'sd2041199, -32'sd1770794, -32'sd774644, -32'sd612726, -32'sd569461, 32'sd1461267, 32'sd1395379, -32'sd1505702, -32'sd1026540, -32'sd968066, -32'sd354831, -32'sd89711, 32'sd95213, 32'sd665494, 32'sd585064, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd322090, 32'sd250265, -32'sd742002, 32'sd105209, -32'sd1482239, -32'sd2464698, -32'sd1158595, -32'sd469072, 32'sd1592136, 32'sd641325, 32'sd1734516, 32'sd600183, 32'sd840250, -32'sd1838511, -32'sd408639, -32'sd1397777, -32'sd1752029, -32'sd1556832, -32'sd736122, 32'sd705846, 32'sd790908, -32'sd215071, 32'sd466126, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd763493, -32'sd542721, 32'sd306113, 32'sd352806, -32'sd716956, 32'sd316665, 32'sd291996, -32'sd14886, -32'sd399170, -32'sd143423, 32'sd539471, 32'sd570468, 32'sd447663, -32'sd447811, 32'sd878283, -32'sd399215, -32'sd399056, 32'sd1899052, 32'sd608540, 32'sd877748, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd890822, -32'sd927951, -32'sd452654, 32'sd221376, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1586395, -32'sd765044, -32'sd652386, -32'sd21007, 32'sd28870, -32'sd987787, 32'sd661042, 32'sd628120, 32'sd2102571, -32'sd532794, 32'sd1003175, -32'sd2236068, -32'sd398090, -32'sd72161, 32'sd93531, -32'sd286312, 32'sd1325532, 32'sd589809, -32'sd321524, -32'sd359325, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd308604, -32'sd333906, -32'sd150743, -32'sd519575, 32'sd243532, -32'sd42184, -32'sd1778219, -32'sd2254211, -32'sd69619, 32'sd1392736, -32'sd323897, -32'sd424607, -32'sd239691, -32'sd682954, 32'sd618314, 32'sd844928, 32'sd1352579, 32'sd156690, 32'sd1102559, 32'sd1745188, 32'sd1781383, 32'sd812699, -32'sd842052, 32'sd118630, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd74835, -32'sd604482, -32'sd1647210, -32'sd226811, 32'sd183332, -32'sd1728453, -32'sd1965315, -32'sd206161, -32'sd439655, -32'sd32891, -32'sd3060721, -32'sd2706361, 32'sd107387, -32'sd1584853, -32'sd2720189, 32'sd1612144, -32'sd479600, -32'sd362404, -32'sd1657021, -32'sd1144481, 32'sd1227161, -32'sd1282666, 32'sd515742, 32'sd606446, -32'sd87971, 32'sd0, 32'sd0, -32'sd285862, -32'sd555976, 32'sd1219042, -32'sd1648502, -32'sd1330468, -32'sd982683, -32'sd1228731, -32'sd1758051, 32'sd287586, 32'sd391762, -32'sd923808, -32'sd907769, -32'sd195038, -32'sd1001849, -32'sd1120128, -32'sd845249, 32'sd368285, 32'sd1950925, 32'sd908013, 32'sd521340, 32'sd395827, -32'sd287619, -32'sd977986, 32'sd5261, 32'sd791018, 32'sd85476, 32'sd480266, 32'sd0, 32'sd562727, -32'sd293029, 32'sd684604, -32'sd447473, -32'sd1111181, -32'sd3651435, -32'sd1807799, -32'sd838444, 32'sd985009, 32'sd2237934, -32'sd106660, -32'sd513632, 32'sd141172, -32'sd888223, -32'sd1928481, -32'sd1000338, 32'sd1768869, 32'sd778408, 32'sd73653, 32'sd856419, 32'sd1225495, -32'sd1926303, -32'sd1906387, -32'sd1529077, 32'sd77392, 32'sd727191, -32'sd1002623, 32'sd0, -32'sd243079, -32'sd468785, -32'sd577967, 32'sd1486392, 32'sd537604, -32'sd4977648, -32'sd1877980, -32'sd827763, 32'sd1779046, 32'sd55221, 32'sd168819, 32'sd747174, -32'sd165251, -32'sd997188, -32'sd1906438, -32'sd247866, 32'sd26700, 32'sd288812, 32'sd425659, 32'sd1950940, -32'sd816914, 32'sd363144, -32'sd1058337, -32'sd1468974, -32'sd558929, -32'sd1477424, 32'sd1491698, -32'sd831811, -32'sd507907, -32'sd2224880, -32'sd1200491, -32'sd1599871, -32'sd3102886, -32'sd3807419, -32'sd2394103, 32'sd1414977, 32'sd958426, 32'sd1512768, 32'sd1886209, 32'sd542279, -32'sd776167, -32'sd307401, 32'sd1242919, 32'sd1541880, 32'sd1502208, 32'sd1229631, -32'sd147361, 32'sd1262831, -32'sd851816, -32'sd1210687, -32'sd1408180, 32'sd710909, -32'sd1398779, 32'sd548500, -32'sd1073116, -32'sd151899, -32'sd187974, 32'sd499461, 32'sd472055, -32'sd748143, -32'sd3633444, -32'sd4603698, -32'sd1856021, 32'sd1027732, 32'sd577140, -32'sd1128187, 32'sd2555914, -32'sd330661, 32'sd164356, -32'sd833623, -32'sd856916, 32'sd512264, 32'sd720869, -32'sd453578, -32'sd3722824, -32'sd2051139, -32'sd2522371, -32'sd2329067, -32'sd1420639, 32'sd1432743, -32'sd2292368, -32'sd470241, 32'sd74687, -32'sd596722, -32'sd1592355, 32'sd482735, -32'sd128625, -32'sd1159890, -32'sd3579684, -32'sd3058313, -32'sd548541, 32'sd167466, -32'sd297725, -32'sd567314, 32'sd1916727, 32'sd472424, 32'sd154968, -32'sd2962916, -32'sd1254123, 32'sd1979013, -32'sd1941221, -32'sd3741426, -32'sd3221512, -32'sd1963472, -32'sd1826142, -32'sd2647804, -32'sd937722, -32'sd973029, 32'sd638307, 32'sd737987, 32'sd324968, -32'sd1075722, 32'sd144303, -32'sd1085895, -32'sd646896, -32'sd939535, -32'sd2365072, -32'sd5589960, -32'sd1813128, 32'sd745070, 32'sd1812617, -32'sd311577, 32'sd1488727, 32'sd462877, -32'sd475198, -32'sd3341138, 32'sd771587, -32'sd934132, -32'sd2565335, -32'sd2388874, -32'sd3401153, -32'sd806775, -32'sd1104653, -32'sd1183347, -32'sd1011814, 32'sd990770, -32'sd298158, 32'sd976484, -32'sd1174324, -32'sd713379, -32'sd478611, 32'sd124260, -32'sd1139032, -32'sd1286681, -32'sd982624, -32'sd3030556, -32'sd1543470, 32'sd1464678, 32'sd2232028, 32'sd778564, 32'sd484235, 32'sd2118844, 32'sd326488, -32'sd2691152, -32'sd2497963, 32'sd1158000, 32'sd379577, 32'sd139111, 32'sd703753, -32'sd1055014, -32'sd831174, -32'sd1928516, 32'sd574628, -32'sd771738, -32'sd1264989, 32'sd936699, -32'sd1811734, -32'sd632002, 32'sd338051, -32'sd1517758, -32'sd96911, -32'sd368977, -32'sd1425721, -32'sd2439339, -32'sd604745, -32'sd597312, -32'sd27286, 32'sd1458109, 32'sd2915674, 32'sd3521323, -32'sd1185371, -32'sd2484658, -32'sd124372, -32'sd2552549, -32'sd262788, -32'sd923162, -32'sd1706800, -32'sd259756, -32'sd43162, 32'sd333916, -32'sd427643, -32'sd380549, -32'sd2659, 32'sd413553, -32'sd694085, -32'sd747436, 32'sd13121, -32'sd245144, -32'sd1113651, 32'sd1353125, -32'sd862276, -32'sd3164856, -32'sd1467244, -32'sd1495199, -32'sd728953, 32'sd1863293, 32'sd216685, 32'sd1756463, -32'sd969612, -32'sd2771469, -32'sd1910047, -32'sd2440121, -32'sd1294381, -32'sd1183081, 32'sd43778, 32'sd1182419, 32'sd731986, 32'sd373849, -32'sd2757565, -32'sd2203432, -32'sd4130626, -32'sd1031112, -32'sd780305, 32'sd739019, -32'sd443504, 32'sd202760, -32'sd1339980, 32'sd6731, 32'sd495094, -32'sd2374707, -32'sd1256255, -32'sd1318875, 32'sd899952, 32'sd1234170, -32'sd184234, 32'sd1435629, 32'sd940654, -32'sd647978, -32'sd1937074, -32'sd441503, -32'sd1190078, 32'sd15040, 32'sd98943, 32'sd1034360, 32'sd695294, -32'sd663278, -32'sd964529, 32'sd327492, -32'sd2167567, -32'sd643852, 32'sd173501, 32'sd701768, 32'sd53365, -32'sd2170151, -32'sd895359, -32'sd460935, 32'sd646549, -32'sd2429704, -32'sd1416895, -32'sd1740443, 32'sd1445373, 32'sd1434800, 32'sd2558245, 32'sd1082595, -32'sd868741, -32'sd1920885, -32'sd1117549, -32'sd2176587, -32'sd672660, -32'sd301949, -32'sd484545, 32'sd956863, 32'sd950044, -32'sd1710727, 32'sd101302, -32'sd1509337, -32'sd1866937, -32'sd1494915, 32'sd284818, 32'sd722444, -32'sd197126, -32'sd1429777, 32'sd706190, -32'sd483420, 32'sd1413155, -32'sd730603, -32'sd526569, -32'sd158638, 32'sd513048, 32'sd1365686, 32'sd1992901, -32'sd437074, 32'sd120158, -32'sd1293502, -32'sd1990067, -32'sd1862866, -32'sd641433, 32'sd2365711, 32'sd1088346, 32'sd544856, 32'sd2143991, -32'sd1998402, 32'sd118515, -32'sd1143536, -32'sd1727703, -32'sd1992872, -32'sd1258992, 32'sd0, -32'sd884182, 32'sd697215, -32'sd2142268, 32'sd529934, 32'sd672779, 32'sd1074497, 32'sd1114284, 32'sd1074335, -32'sd722257, 32'sd1062357, 32'sd1507715, 32'sd560154, -32'sd111689, 32'sd45315, -32'sd2419084, -32'sd61851, 32'sd2797579, 32'sd2459367, 32'sd1266903, 32'sd1679490, 32'sd1576467, -32'sd571407, -32'sd2305416, -32'sd545950, -32'sd1699210, -32'sd615642, -32'sd1269972, -32'sd104229, -32'sd304127, -32'sd664861, 32'sd264587, 32'sd620676, 32'sd1350047, 32'sd745108, 32'sd427618, 32'sd2054392, -32'sd124524, 32'sd268482, 32'sd182966, -32'sd712368, 32'sd710, 32'sd159607, 32'sd1711299, 32'sd169641, 32'sd2047316, 32'sd848037, 32'sd955046, 32'sd1203548, -32'sd506567, -32'sd2161662, -32'sd2842453, -32'sd1356380, -32'sd2386131, 32'sd1170562, -32'sd381689, -32'sd3193, -32'sd559051, 32'sd1018369, 32'sd1577759, 32'sd247981, 32'sd367093, 32'sd2216273, 32'sd1140105, 32'sd1593804, 32'sd61283, -32'sd439989, 32'sd176262, -32'sd826623, -32'sd303980, -32'sd639716, 32'sd2319214, 32'sd2240618, 32'sd285570, 32'sd238588, 32'sd1781329, 32'sd1954323, -32'sd549263, -32'sd1882328, -32'sd1486439, -32'sd41743, -32'sd2487481, -32'sd983363, -32'sd428989, 32'sd0, 32'sd87530, 32'sd1240975, -32'sd495091, 32'sd174758, -32'sd1528968, 32'sd1059085, -32'sd759938, 32'sd76431, 32'sd269796, -32'sd502390, -32'sd1081147, -32'sd3884138, -32'sd2317476, -32'sd976195, 32'sd1987020, 32'sd1380939, 32'sd2843108, 32'sd2247379, 32'sd2231759, -32'sd131519, -32'sd384554, 32'sd1379862, -32'sd2513515, -32'sd1328722, -32'sd792639, 32'sd121899, 32'sd420565, 32'sd319208, -32'sd1488549, -32'sd610043, 32'sd292478, -32'sd212114, -32'sd575845, -32'sd836189, -32'sd2408134, -32'sd786472, -32'sd1155951, -32'sd1317004, -32'sd1097275, -32'sd1785822, -32'sd3106232, 32'sd1218685, 32'sd549352, 32'sd1259514, 32'sd1472701, 32'sd1433528, 32'sd720676, 32'sd2411582, -32'sd34306, 32'sd1181344, -32'sd2825286, -32'sd874659, -32'sd435994, 32'sd82449, -32'sd729078, -32'sd346448, -32'sd256696, 32'sd348052, -32'sd628475, 32'sd898197, 32'sd521519, -32'sd184614, -32'sd2169367, -32'sd444071, -32'sd1360328, 32'sd462068, -32'sd1362975, -32'sd2284592, -32'sd2646131, 32'sd1118040, -32'sd1062855, 32'sd2261528, 32'sd2459298, 32'sd2003027, 32'sd162582, 32'sd1003673, -32'sd400919, 32'sd209247, -32'sd807332, 32'sd239458, -32'sd1040402, 32'sd856031, -32'sd667195, 32'sd0, 32'sd175317, 32'sd129327, 32'sd453778, 32'sd251220, 32'sd1178292, 32'sd202182, -32'sd1244799, 32'sd45763, -32'sd2030847, -32'sd1904630, -32'sd522524, -32'sd395224, -32'sd803054, 32'sd9520, 32'sd540939, 32'sd1967576, 32'sd2342150, 32'sd1166052, 32'sd1024509, 32'sd470397, -32'sd1077135, -32'sd1696415, -32'sd431042, -32'sd652241, -32'sd56654, 32'sd99445, 32'sd0, 32'sd0, 32'sd0, -32'sd1230234, 32'sd239621, 32'sd892055, -32'sd1427768, -32'sd2117106, -32'sd1388370, -32'sd1511592, -32'sd1304686, -32'sd385721, -32'sd1141883, -32'sd1801555, 32'sd1180639, 32'sd173805, 32'sd879434, 32'sd1994715, 32'sd2093580, 32'sd589337, 32'sd1259803, -32'sd884268, -32'sd2578218, -32'sd230676, -32'sd276669, 32'sd416439, -32'sd209527, 32'sd221411, 32'sd0, 32'sd0, 32'sd0, -32'sd857115, 32'sd703298, -32'sd348681, 32'sd340188, 32'sd884305, -32'sd1107357, -32'sd1064167, 32'sd1987975, 32'sd137102, 32'sd58305, -32'sd583080, 32'sd47545, 32'sd377175, 32'sd2058361, 32'sd3555883, 32'sd1278274, 32'sd520206, -32'sd1813671, -32'sd267075, 32'sd629541, 32'sd720573, -32'sd162413, -32'sd10117, 32'sd284043, -32'sd500657, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd148204, -32'sd876439, 32'sd937470, -32'sd674411, -32'sd566880, -32'sd157874, 32'sd240595, -32'sd2804796, 32'sd610714, -32'sd299917, 32'sd138011, -32'sd664314, 32'sd673437, 32'sd728730, -32'sd2022591, -32'sd1781269, 32'sd940047, 32'sd460091, 32'sd258845, -32'sd399753, 32'sd925158, 32'sd1332856, -32'sd546317, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd309721, 32'sd1009577, 32'sd984539, 32'sd815237, -32'sd8271, 32'sd57181, 32'sd603314, -32'sd1207641, 32'sd107129, -32'sd580044, -32'sd334547, 32'sd1850843, -32'sd1274753, 32'sd631243, 32'sd598191, 32'sd379787, -32'sd1564972, -32'sd32838, -32'sd302725, -32'sd148001, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd540057, 32'sd2286985, 32'sd1125399, 32'sd1692024, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd455485, 32'sd1953993, 32'sd1335290, 32'sd1737764, 32'sd992644, 32'sd1803740, 32'sd2106131, 32'sd988712, 32'sd351915, -32'sd436650, -32'sd1562545, 32'sd910684, 32'sd2259350, 32'sd2209424, 32'sd1492276, 32'sd604845, -32'sd193167, -32'sd207726, 32'sd1441062, 32'sd672101, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1147843, -32'sd406068, -32'sd23792, 32'sd1473202, 32'sd446532, -32'sd423440, 32'sd1015456, 32'sd1397272, 32'sd581523, -32'sd548515, -32'sd1139499, -32'sd719725, 32'sd357644, 32'sd754438, 32'sd837930, 32'sd986364, 32'sd340164, 32'sd3798424, 32'sd3019456, 32'sd1220979, -32'sd90338, 32'sd2458057, 32'sd102608, 32'sd1418857, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd351410, 32'sd559737, -32'sd136121, -32'sd84000, -32'sd668000, -32'sd2097876, -32'sd764385, 32'sd1238980, 32'sd98404, 32'sd1155075, -32'sd269158, 32'sd1322588, 32'sd8534, -32'sd1001127, -32'sd768149, 32'sd255174, 32'sd1114595, 32'sd1011938, 32'sd696819, 32'sd90658, -32'sd686499, -32'sd2720968, -32'sd1104474, -32'sd1171869, 32'sd858860, 32'sd0, 32'sd0, 32'sd871710, 32'sd521715, -32'sd5991, -32'sd376670, -32'sd628151, -32'sd2369577, -32'sd1926569, -32'sd1622483, -32'sd1130998, -32'sd903048, 32'sd1055989, 32'sd569248, -32'sd293427, -32'sd1189992, -32'sd1116309, -32'sd1321925, -32'sd1159002, -32'sd730960, -32'sd186935, -32'sd1892664, -32'sd494914, -32'sd1158804, 32'sd473500, 32'sd179831, 32'sd1018751, 32'sd1373823, 32'sd797067, 32'sd0, 32'sd869355, -32'sd746857, -32'sd111726, -32'sd1617610, -32'sd1464724, -32'sd486203, -32'sd2491052, -32'sd1723157, -32'sd1874432, 32'sd267667, 32'sd458790, -32'sd204155, 32'sd304914, 32'sd483493, 32'sd78685, -32'sd306920, 32'sd627611, -32'sd42004, 32'sd1229352, 32'sd1849492, 32'sd2090967, 32'sd664312, -32'sd291711, 32'sd2088690, 32'sd2092726, 32'sd2214984, -32'sd1091933, 32'sd0, 32'sd548015, -32'sd864572, -32'sd457468, -32'sd2192046, -32'sd998073, -32'sd1270277, 32'sd115355, -32'sd2131949, -32'sd2926684, -32'sd151159, 32'sd1729899, 32'sd123393, -32'sd281447, 32'sd669002, -32'sd296682, 32'sd1240273, 32'sd1684274, 32'sd1827112, 32'sd1393406, 32'sd1729337, 32'sd384132, 32'sd8815, -32'sd176731, -32'sd132785, -32'sd656022, 32'sd801277, -32'sd246238, 32'sd1700487, -32'sd1102157, -32'sd226736, 32'sd379527, -32'sd1616783, -32'sd737034, 32'sd1490623, -32'sd1439599, -32'sd717816, -32'sd306802, 32'sd903576, 32'sd1243042, -32'sd2267910, -32'sd1897244, -32'sd215786, -32'sd1598308, -32'sd1742922, 32'sd195878, -32'sd878245, 32'sd2395336, 32'sd1047288, 32'sd922631, 32'sd2896079, -32'sd463666, -32'sd409679, 32'sd232195, -32'sd1188843, -32'sd282023, -32'sd20067, 32'sd393484, 32'sd1351528, -32'sd1069388, -32'sd1885979, 32'sd282950, -32'sd399991, -32'sd578321, -32'sd1464861, -32'sd1013434, 32'sd1321264, 32'sd1858974, -32'sd1304697, -32'sd1902579, -32'sd997994, -32'sd2102424, -32'sd185517, -32'sd87271, -32'sd712745, 32'sd1084197, 32'sd3136499, 32'sd860984, 32'sd1369419, 32'sd1142332, -32'sd685857, 32'sd603387, -32'sd755702, -32'sd207962, 32'sd749777, -32'sd336113, -32'sd602095, 32'sd2809360, 32'sd3534748, 32'sd2356619, 32'sd1634898, 32'sd43050, -32'sd90267, 32'sd65310, -32'sd264690, 32'sd1020232, -32'sd1785577, -32'sd1619130, -32'sd421871, -32'sd3609192, -32'sd4092696, -32'sd3138433, 32'sd815800, 32'sd1116757, 32'sd2011547, 32'sd1366732, 32'sd1834362, 32'sd1001423, -32'sd253296, 32'sd1552827, 32'sd562065, -32'sd842382, -32'sd208421, 32'sd73062, 32'sd1089928, 32'sd44615, 32'sd1098152, 32'sd2088134, -32'sd166517, -32'sd363648, 32'sd509517, 32'sd1874108, 32'sd2258011, 32'sd2921319, 32'sd1180894, 32'sd472298, -32'sd1062968, -32'sd1037599, -32'sd1414888, -32'sd2073859, -32'sd190914, -32'sd94642, 32'sd1359676, 32'sd169460, 32'sd2272569, 32'sd1504946, -32'sd1108680, -32'sd647388, -32'sd1258506, 32'sd28034, 32'sd507199, 32'sd1732597, 32'sd1583787, 32'sd651913, 32'sd1232988, 32'sd44295, -32'sd1319155, 32'sd1648454, -32'sd516227, 32'sd1914633, 32'sd1592396, 32'sd75773, 32'sd517523, 32'sd1890402, 32'sd1054057, -32'sd1208067, -32'sd2082481, -32'sd2530160, -32'sd1304200, 32'sd180813, 32'sd703968, 32'sd632035, 32'sd2695981, 32'sd1302764, 32'sd730303, 32'sd1494384, 32'sd1102097, 32'sd1018850, 32'sd1164431, 32'sd821232, -32'sd288909, -32'sd132948, 32'sd348721, -32'sd1352400, 32'sd974590, 32'sd2353024, 32'sd1009911, 32'sd2073267, 32'sd1063347, 32'sd914650, -32'sd153508, -32'sd1660829, -32'sd2836426, -32'sd1192919, -32'sd2554878, -32'sd2992485, -32'sd1919918, -32'sd1694991, 32'sd348979, -32'sd889335, 32'sd373877, 32'sd1319379, 32'sd120747, -32'sd384709, 32'sd238054, 32'sd2227244, 32'sd1005974, -32'sd79068, -32'sd1391402, -32'sd2251166, 32'sd412034, 32'sd295437, 32'sd1328204, 32'sd806641, -32'sd253517, -32'sd717867, -32'sd678017, -32'sd1118637, -32'sd2231658, -32'sd511808, -32'sd1739776, -32'sd2795545, -32'sd221681, -32'sd1443158, -32'sd2231253, -32'sd1013462, 32'sd287665, -32'sd58965, -32'sd855182, -32'sd437595, 32'sd2179112, 32'sd843706, 32'sd1988346, 32'sd2886879, 32'sd1188734, -32'sd907214, -32'sd214922, -32'sd2488677, -32'sd476170, 32'sd804812, -32'sd1204271, -32'sd277628, 32'sd64252, -32'sd2103390, -32'sd1432469, -32'sd2618954, -32'sd1832938, -32'sd2148582, -32'sd797373, -32'sd2873493, -32'sd2540728, 32'sd1706552, 32'sd906031, -32'sd385785, 32'sd1724476, -32'sd387317, -32'sd83915, 32'sd740615, -32'sd194894, 32'sd770868, -32'sd1094197, 32'sd2904623, 32'sd1049575, 32'sd534406, -32'sd344044, -32'sd393500, 32'sd760145, -32'sd380860, -32'sd119212, -32'sd737262, -32'sd186422, 32'sd323666, -32'sd1681809, -32'sd278085, -32'sd2056327, -32'sd633717, -32'sd903354, -32'sd1193357, -32'sd914178, 32'sd1594726, 32'sd1152508, 32'sd2061651, 32'sd89265, -32'sd149130, -32'sd899812, -32'sd141036, -32'sd56183, -32'sd1438634, 32'sd463186, 32'sd792383, 32'sd1009871, -32'sd1185847, -32'sd228257, 32'sd759228, -32'sd630901, 32'sd1723656, 32'sd1361371, 32'sd1939899, -32'sd27019, 32'sd240872, 32'sd466699, 32'sd342682, -32'sd1691656, 32'sd51581, -32'sd1005152, -32'sd547925, -32'sd863000, 32'sd2685164, 32'sd158415, 32'sd903544, 32'sd1646396, 32'sd201196, -32'sd729567, -32'sd472652, -32'sd621542, 32'sd1212559, 32'sd1268807, 32'sd1751034, 32'sd0, 32'sd886912, -32'sd1244213, -32'sd522894, 32'sd2113654, 32'sd2121119, -32'sd10004, 32'sd2079753, 32'sd192863, 32'sd1842494, -32'sd1005788, -32'sd1385742, -32'sd1410959, -32'sd86286, 32'sd838273, -32'sd353356, -32'sd169845, 32'sd1302413, 32'sd1407782, -32'sd1589054, 32'sd1085625, -32'sd989467, -32'sd612059, 32'sd539928, 32'sd1150845, 32'sd1329202, -32'sd651155, 32'sd87509, -32'sd329984, 32'sd902029, 32'sd701724, -32'sd1571574, 32'sd1543385, 32'sd1841575, -32'sd376641, 32'sd1418445, 32'sd1111534, 32'sd242200, -32'sd2982105, -32'sd2174805, -32'sd3087533, -32'sd1039945, 32'sd231402, -32'sd906025, -32'sd1976064, -32'sd145637, 32'sd807176, -32'sd2424676, 32'sd596969, 32'sd330532, -32'sd1091940, 32'sd968968, 32'sd152997, -32'sd313743, -32'sd323048, 32'sd1852010, 32'sd879374, -32'sd1135536, 32'sd435227, -32'sd1206314, 32'sd2020277, 32'sd1820361, 32'sd43207, 32'sd534635, 32'sd1995022, 32'sd1928910, -32'sd1609210, -32'sd2106139, -32'sd149669, -32'sd986166, -32'sd1477004, -32'sd853119, -32'sd253762, -32'sd298274, -32'sd1365597, -32'sd634085, -32'sd1401031, -32'sd149779, -32'sd1202929, -32'sd81678, -32'sd757423, -32'sd196472, -32'sd1433428, -32'sd594466, 32'sd0, -32'sd288306, 32'sd323717, 32'sd508046, 32'sd1843540, 32'sd2360240, 32'sd1785373, 32'sd2727020, 32'sd1001070, -32'sd739917, -32'sd576120, 32'sd413895, -32'sd1575494, -32'sd1320775, -32'sd1953777, -32'sd2854761, -32'sd2631438, -32'sd2417281, -32'sd1682846, 32'sd135677, -32'sd513884, -32'sd1084442, -32'sd773899, -32'sd1017619, -32'sd781882, -32'sd1404271, -32'sd1466685, 32'sd961653, 32'sd1053663, 32'sd376244, -32'sd80847, 32'sd344074, 32'sd539139, 32'sd1590389, 32'sd2142729, 32'sd2154048, 32'sd1726772, 32'sd58195, -32'sd587559, 32'sd460819, -32'sd1025400, -32'sd1118845, -32'sd1130621, 32'sd22672, -32'sd1030506, 32'sd595275, -32'sd1162308, -32'sd1053124, -32'sd536874, 32'sd227192, 32'sd701703, -32'sd533180, 32'sd3121, -32'sd659425, 32'sd847717, 32'sd1173297, 32'sd1306810, 32'sd311023, -32'sd180917, 32'sd1754602, -32'sd170731, 32'sd346124, 32'sd3389368, 32'sd1942977, 32'sd268031, -32'sd988612, -32'sd255288, 32'sd538357, 32'sd924974, -32'sd1601798, -32'sd1077981, -32'sd147198, 32'sd552942, -32'sd546010, -32'sd1478565, -32'sd344527, -32'sd488817, 32'sd419340, -32'sd1030189, -32'sd2387269, -32'sd614463, -32'sd173639, 32'sd656156, 32'sd2030714, 32'sd0, 32'sd893456, 32'sd1800107, 32'sd1840265, 32'sd250858, -32'sd589943, 32'sd1610876, 32'sd1970465, 32'sd2392641, -32'sd515284, 32'sd915023, -32'sd716399, -32'sd1457713, -32'sd685085, -32'sd991972, 32'sd53052, 32'sd90135, 32'sd1058975, 32'sd232701, 32'sd140138, 32'sd524239, -32'sd1576750, -32'sd56009, -32'sd682914, 32'sd594062, -32'sd251871, -32'sd116567, 32'sd0, 32'sd0, 32'sd0, 32'sd381563, 32'sd1233971, 32'sd2336767, 32'sd232782, 32'sd418270, 32'sd1896962, 32'sd2435171, 32'sd538939, 32'sd1211679, 32'sd82065, 32'sd651530, 32'sd358764, -32'sd2151509, -32'sd1252551, -32'sd1642438, -32'sd668556, 32'sd615919, 32'sd588849, 32'sd529113, 32'sd582369, -32'sd236558, 32'sd549813, -32'sd1034390, 32'sd1070140, 32'sd738725, 32'sd0, 32'sd0, 32'sd0, -32'sd1182245, -32'sd193380, -32'sd458219, -32'sd1790308, -32'sd1787036, -32'sd579614, 32'sd848259, 32'sd1408394, 32'sd1363258, -32'sd687130, 32'sd440913, 32'sd825149, 32'sd1368721, -32'sd429169, 32'sd1101113, -32'sd1237844, -32'sd716593, 32'sd2102206, 32'sd734331, 32'sd1457383, -32'sd1226803, 32'sd872164, -32'sd274242, 32'sd958569, 32'sd1743935, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1564392, 32'sd365072, -32'sd1763911, -32'sd704755, -32'sd988591, -32'sd344660, 32'sd588170, 32'sd1059761, 32'sd41381, 32'sd1208059, -32'sd1252337, -32'sd331385, -32'sd755308, 32'sd2041021, 32'sd288128, 32'sd1321626, 32'sd1499142, 32'sd5889, -32'sd554428, 32'sd2418818, 32'sd1438863, -32'sd393462, 32'sd1760083, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1709196, 32'sd993463, 32'sd469403, 32'sd1313508, 32'sd39221, -32'sd148601, 32'sd1661594, -32'sd243917, 32'sd1383955, 32'sd784847, 32'sd1950962, 32'sd1409673, 32'sd243677, 32'sd661043, 32'sd833402, -32'sd1058307, 32'sd185459, 32'sd214897, 32'sd993306, 32'sd1529708, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd98403, -32'sd260283, -32'sd296132, -32'sd5841, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd725330, -32'sd907728, -32'sd198640, 32'sd516755, 32'sd83373, 32'sd59713, 32'sd1797483, -32'sd1074514, 32'sd75591, -32'sd1102146, 32'sd128342, 32'sd133196, 32'sd906590, 32'sd1172352, 32'sd1153552, -32'sd734669, 32'sd1463765, 32'sd703823, 32'sd1739129, 32'sd159505, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1158096, 32'sd1608416, 32'sd452371, -32'sd584794, 32'sd289929, -32'sd720072, -32'sd251067, -32'sd703508, 32'sd1001977, 32'sd111118, -32'sd1082686, -32'sd344175, -32'sd222642, 32'sd1512805, 32'sd1857204, -32'sd243717, 32'sd2072811, 32'sd3643714, 32'sd1301300, -32'sd287349, 32'sd410462, 32'sd1563250, -32'sd1569, 32'sd819845, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd558465, 32'sd485197, 32'sd409962, -32'sd1539693, -32'sd1455589, -32'sd338291, -32'sd1002928, 32'sd1235750, 32'sd585775, -32'sd976551, 32'sd805446, 32'sd2389956, 32'sd1952164, 32'sd1466575, 32'sd209804, -32'sd1148987, -32'sd129479, -32'sd444394, -32'sd1492872, -32'sd522833, 32'sd1093944, 32'sd204908, 32'sd996565, 32'sd1144009, 32'sd236559, 32'sd0, 32'sd0, 32'sd169061, 32'sd683956, -32'sd1335112, 32'sd391921, -32'sd1717, 32'sd928895, -32'sd1240305, -32'sd499003, -32'sd851602, -32'sd955752, 32'sd1190397, 32'sd442523, -32'sd1062337, 32'sd2066838, 32'sd2893906, -32'sd800914, -32'sd382993, -32'sd1092646, -32'sd698916, -32'sd809479, 32'sd2184483, 32'sd287478, 32'sd1932473, -32'sd685102, 32'sd1644938, 32'sd197400, 32'sd718485, 32'sd0, 32'sd313187, -32'sd674191, 32'sd198694, -32'sd390238, 32'sd270284, -32'sd55611, -32'sd801826, 32'sd1494525, -32'sd1393206, 32'sd588863, 32'sd1084465, 32'sd896643, 32'sd1529776, -32'sd191273, 32'sd2357762, 32'sd668109, 32'sd940444, 32'sd1778305, -32'sd177367, 32'sd1877997, 32'sd685384, 32'sd564954, 32'sd1868578, 32'sd1597270, 32'sd659231, 32'sd308827, 32'sd807281, 32'sd0, -32'sd423803, -32'sd112685, 32'sd1018417, 32'sd847828, 32'sd281339, -32'sd870579, -32'sd562741, 32'sd2255275, 32'sd568162, -32'sd762194, 32'sd1960880, 32'sd2118695, 32'sd3404405, 32'sd1434263, 32'sd3167035, 32'sd2808154, 32'sd2218021, 32'sd1274337, 32'sd52594, -32'sd833694, 32'sd60209, -32'sd29457, -32'sd1908731, -32'sd1407795, -32'sd1225268, -32'sd690242, 32'sd1066154, 32'sd1496666, 32'sd998418, 32'sd1517057, 32'sd926472, -32'sd81689, -32'sd552515, 32'sd250076, -32'sd120908, 32'sd2007882, 32'sd993316, 32'sd1165228, 32'sd1545097, 32'sd3148187, 32'sd2641985, 32'sd2312724, -32'sd100840, 32'sd221165, -32'sd2461310, -32'sd1195728, -32'sd705098, -32'sd1369348, -32'sd716132, -32'sd434988, -32'sd2450472, -32'sd1332586, 32'sd1304849, -32'sd1274173, 32'sd30508, 32'sd1267290, 32'sd1326591, 32'sd280576, -32'sd1105267, -32'sd2596996, 32'sd729345, -32'sd868042, 32'sd1136992, 32'sd1804520, 32'sd88272, 32'sd1996493, 32'sd3037581, 32'sd1888664, -32'sd524125, 32'sd359516, -32'sd3408657, -32'sd5123206, -32'sd4029413, -32'sd3499283, -32'sd3669808, -32'sd2745932, -32'sd1335096, -32'sd1248105, -32'sd2613443, -32'sd1571481, -32'sd1496974, -32'sd246988, -32'sd617505, -32'sd386353, 32'sd1960384, 32'sd1401198, -32'sd1423604, 32'sd151572, -32'sd196383, 32'sd1928912, -32'sd186847, 32'sd1798026, 32'sd218108, 32'sd1394608, 32'sd1851934, -32'sd2061260, -32'sd3103116, -32'sd1396861, -32'sd2335239, -32'sd3244309, -32'sd1908236, -32'sd3973834, -32'sd4876414, -32'sd4422285, -32'sd3864130, -32'sd2996321, -32'sd3192412, -32'sd1910590, -32'sd345197, -32'sd279130, 32'sd94269, 32'sd87805, -32'sd275360, 32'sd1383086, -32'sd1257849, -32'sd1356311, 32'sd1193377, 32'sd1351100, 32'sd143767, -32'sd943141, 32'sd78609, -32'sd240963, -32'sd425110, -32'sd3415033, 32'sd39328, 32'sd1064632, 32'sd327841, 32'sd1379230, 32'sd577868, 32'sd1199555, -32'sd944478, -32'sd1724359, -32'sd2043768, -32'sd200984, -32'sd1235071, -32'sd799545, -32'sd582029, -32'sd451357, 32'sd358142, 32'sd846438, -32'sd307823, -32'sd1410667, -32'sd620134, -32'sd1561411, -32'sd438560, 32'sd1265842, 32'sd1009993, -32'sd54008, -32'sd1039969, 32'sd1144131, 32'sd509417, -32'sd391377, 32'sd3993861, 32'sd2445489, 32'sd4339082, 32'sd5514425, 32'sd5128042, 32'sd2110810, 32'sd221055, 32'sd632316, 32'sd1287224, -32'sd754833, 32'sd112297, -32'sd282181, -32'sd3166953, -32'sd104579, -32'sd338378, 32'sd394542, 32'sd348707, 32'sd683192, -32'sd207743, 32'sd970634, 32'sd32797, 32'sd58360, 32'sd1389474, 32'sd1918568, 32'sd1201136, -32'sd169592, 32'sd704190, -32'sd229437, 32'sd1868980, 32'sd899677, 32'sd3033372, 32'sd1699091, 32'sd1141342, 32'sd1999417, 32'sd2322999, 32'sd2924997, 32'sd1255240, 32'sd865749, 32'sd2095085, -32'sd937373, -32'sd4854880, -32'sd2070216, -32'sd470498, 32'sd691276, 32'sd938241, 32'sd934108, 32'sd210461, -32'sd227072, 32'sd1138374, 32'sd813594, 32'sd1021963, 32'sd14418, 32'sd719899, 32'sd466975, -32'sd1663470, -32'sd621341, -32'sd2351685, -32'sd2404023, -32'sd138160, 32'sd1435926, -32'sd895808, -32'sd133060, 32'sd836590, 32'sd2264230, 32'sd990969, 32'sd990994, 32'sd2420693, -32'sd232313, -32'sd1502613, 32'sd112363, -32'sd525170, 32'sd911339, 32'sd450925, 32'sd655011, -32'sd1710707, -32'sd894374, -32'sd1459801, 32'sd1162734, 32'sd247889, 32'sd461442, -32'sd1048619, 32'sd1017970, 32'sd1166106, 32'sd874147, -32'sd151010, -32'sd1853998, -32'sd2949127, -32'sd748613, -32'sd1081709, 32'sd1831903, 32'sd1193269, 32'sd52134, 32'sd746011, 32'sd611680, 32'sd2857170, 32'sd1348522, -32'sd57013, 32'sd814007, 32'sd344872, 32'sd1567154, -32'sd1258467, -32'sd370719, -32'sd2380552, -32'sd2354222, -32'sd1806435, 32'sd109429, -32'sd1032309, -32'sd478227, -32'sd1098881, -32'sd114530, -32'sd1218099, -32'sd929447, -32'sd2341675, -32'sd3547961, -32'sd1897351, -32'sd587256, -32'sd215668, 32'sd197146, -32'sd180900, 32'sd1016807, 32'sd97933, -32'sd45769, 32'sd153616, -32'sd429492, -32'sd1353872, 32'sd59801, -32'sd221918, 32'sd163547, -32'sd717510, -32'sd1847966, -32'sd213529, -32'sd342342, -32'sd556182, -32'sd419139, -32'sd2510223, -32'sd2574378, -32'sd2355160, -32'sd1415324, -32'sd2449336, -32'sd2583493, -32'sd1688597, -32'sd2298574, -32'sd372543, -32'sd1082732, 32'sd64469, -32'sd1040990, 32'sd1495259, 32'sd1239163, 32'sd2645226, -32'sd797656, 32'sd389583, 32'sd763543, -32'sd1350201, -32'sd827001, -32'sd1057315, 32'sd0, 32'sd838323, 32'sd250732, 32'sd1119937, -32'sd1886039, -32'sd292078, 32'sd1412398, -32'sd798282, 32'sd341086, -32'sd1035530, -32'sd2245496, -32'sd1294767, -32'sd2691120, -32'sd3321512, 32'sd161046, -32'sd753552, 32'sd417944, -32'sd580230, 32'sd1115670, 32'sd98150, -32'sd541557, -32'sd167946, 32'sd552439, -32'sd783836, 32'sd1174408, 32'sd875329, 32'sd768137, 32'sd342896, -32'sd506907, 32'sd346068, -32'sd548549, 32'sd1043561, 32'sd1290087, 32'sd1697953, -32'sd1110564, -32'sd1546585, -32'sd464889, -32'sd1652285, -32'sd214935, -32'sd1042293, 32'sd178617, -32'sd1229796, 32'sd86144, 32'sd1411976, 32'sd929920, 32'sd1318595, 32'sd467735, 32'sd71043, 32'sd50996, -32'sd1255060, -32'sd1733996, -32'sd105715, 32'sd298700, -32'sd465837, -32'sd385580, -32'sd851232, 32'sd931426, -32'sd74785, -32'sd526751, -32'sd13647, 32'sd113325, 32'sd828378, -32'sd682181, -32'sd686727, -32'sd1860225, -32'sd539810, -32'sd2392099, -32'sd676664, -32'sd96325, -32'sd703189, 32'sd858620, 32'sd304178, -32'sd338527, -32'sd521160, -32'sd1725747, 32'sd52682, -32'sd2055103, -32'sd639302, -32'sd1206552, 32'sd619360, 32'sd1153440, 32'sd82589, -32'sd217384, -32'sd248693, 32'sd0, 32'sd330830, -32'sd1429691, 32'sd1412732, 32'sd1390527, 32'sd555128, 32'sd55183, 32'sd268374, 32'sd403846, 32'sd505977, 32'sd1010334, 32'sd817206, 32'sd480459, -32'sd788949, 32'sd86110, -32'sd335041, -32'sd203627, 32'sd583199, -32'sd1466183, -32'sd154942, -32'sd1085190, 32'sd49078, -32'sd892434, 32'sd553362, 32'sd1606456, 32'sd174398, -32'sd324004, 32'sd693458, 32'sd1132182, -32'sd9658, 32'sd1338569, -32'sd1253408, -32'sd627904, -32'sd235018, 32'sd1561488, 32'sd383050, 32'sd1191911, 32'sd351925, 32'sd1166933, 32'sd551540, 32'sd588366, -32'sd925494, 32'sd904407, 32'sd879139, -32'sd1635429, 32'sd173118, -32'sd362010, -32'sd1385304, 32'sd1036829, 32'sd1583714, -32'sd905527, 32'sd137092, 32'sd1658128, 32'sd651795, 32'sd261433, 32'sd582391, 32'sd1933413, 32'sd1396019, 32'sd402342, 32'sd373441, 32'sd395842, -32'sd1898033, -32'sd1114297, -32'sd171966, 32'sd1025831, 32'sd1206559, 32'sd2109512, 32'sd604466, 32'sd1035254, 32'sd230878, 32'sd1019166, 32'sd365001, -32'sd139998, -32'sd453690, -32'sd586445, -32'sd2346319, -32'sd745284, -32'sd500248, 32'sd502384, 32'sd1863337, 32'sd745025, 32'sd246292, 32'sd319676, 32'sd506910, 32'sd0, -32'sd70418, -32'sd328619, -32'sd413403, 32'sd467160, 32'sd1199359, -32'sd1473977, 32'sd99760, 32'sd2207129, 32'sd1780006, 32'sd236729, 32'sd270350, 32'sd332710, 32'sd1088999, 32'sd13826, 32'sd257909, -32'sd118841, 32'sd438118, 32'sd31164, -32'sd893228, 32'sd1393653, -32'sd426237, 32'sd483355, 32'sd122509, 32'sd946713, -32'sd154871, 32'sd112638, 32'sd0, 32'sd0, 32'sd0, -32'sd978486, 32'sd540143, -32'sd970347, 32'sd684799, 32'sd485525, 32'sd1573983, 32'sd3027241, 32'sd1071900, 32'sd2098242, 32'sd235571, -32'sd1322749, -32'sd2618104, -32'sd1704983, 32'sd385031, 32'sd1688497, -32'sd31646, -32'sd845540, 32'sd1035458, -32'sd130845, 32'sd122571, -32'sd888478, 32'sd741927, 32'sd1215995, -32'sd926586, -32'sd1333340, 32'sd0, 32'sd0, 32'sd0, 32'sd636377, 32'sd973471, -32'sd1465313, -32'sd484418, 32'sd2699981, 32'sd1443085, 32'sd1288750, 32'sd1983766, 32'sd57114, 32'sd424540, 32'sd1509269, -32'sd500924, 32'sd594223, 32'sd2727120, 32'sd2911490, -32'sd538623, -32'sd1570431, 32'sd1823204, -32'sd871700, -32'sd1111773, -32'sd2495077, -32'sd854709, -32'sd2025146, 32'sd812394, 32'sd301012, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1547645, -32'sd338557, 32'sd939932, 32'sd39301, 32'sd651213, -32'sd707118, -32'sd1425766, 32'sd175486, 32'sd1340626, 32'sd515937, 32'sd925394, 32'sd1780874, 32'sd1004228, 32'sd239350, 32'sd949325, -32'sd360756, -32'sd249733, 32'sd149938, -32'sd1432929, -32'sd56229, -32'sd227169, 32'sd332943, -32'sd73848, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd264790, -32'sd887383, 32'sd1524545, 32'sd1381595, 32'sd1029349, 32'sd962459, -32'sd244312, -32'sd631606, -32'sd50654, -32'sd272291, 32'sd1293356, 32'sd343792, -32'sd1065558, 32'sd1335042, -32'sd1387917, -32'sd1216209, 32'sd704880, -32'sd319440, 32'sd147293, 32'sd521937, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd197037, -32'sd1180780, 32'sd530883, 32'sd95340, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd342268, -32'sd870943, -32'sd515046, -32'sd922477, -32'sd580079, -32'sd1305913, -32'sd1084190, -32'sd778492, -32'sd974296, 32'sd586145, -32'sd991862, -32'sd1431954, -32'sd1089820, -32'sd1479320, -32'sd105748, -32'sd595282, 32'sd1103484, 32'sd66567, -32'sd1006979, 32'sd382085, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd839199, -32'sd94405, -32'sd766084, -32'sd1064686, 32'sd372809, -32'sd291870, -32'sd985659, 32'sd652251, -32'sd565516, -32'sd2938554, 32'sd2166700, 32'sd558553, -32'sd606768, -32'sd1364899, -32'sd196454, -32'sd224901, 32'sd486662, -32'sd1483650, -32'sd156669, -32'sd1176597, -32'sd1455909, -32'sd753887, -32'sd214601, -32'sd870591, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd172772, -32'sd458470, -32'sd854654, -32'sd646280, 32'sd991860, -32'sd911794, -32'sd1422602, -32'sd928282, -32'sd578602, -32'sd2355531, -32'sd2028350, -32'sd2067192, -32'sd1164626, -32'sd362750, -32'sd394526, -32'sd1627407, 32'sd403581, -32'sd616772, 32'sd817209, 32'sd699852, -32'sd925909, -32'sd145812, -32'sd355545, 32'sd189507, -32'sd399584, 32'sd0, 32'sd0, -32'sd381519, -32'sd554114, -32'sd920616, -32'sd795701, 32'sd468264, -32'sd22184, 32'sd280532, -32'sd1729644, -32'sd2106899, -32'sd1835918, -32'sd2240714, -32'sd367936, -32'sd2642897, -32'sd1866226, -32'sd3835921, -32'sd3586905, -32'sd1309019, -32'sd758932, -32'sd382193, 32'sd1045400, 32'sd1963501, 32'sd1140555, -32'sd562047, -32'sd239627, -32'sd1064843, -32'sd1377412, 32'sd1395421, 32'sd0, 32'sd161076, -32'sd1027186, -32'sd1211808, -32'sd2232975, 32'sd168841, 32'sd377222, 32'sd1367558, 32'sd2235126, -32'sd318475, 32'sd1548509, 32'sd350241, 32'sd2255052, -32'sd80155, -32'sd511461, 32'sd140934, -32'sd827921, 32'sd1368673, -32'sd2394942, -32'sd3794979, -32'sd1039881, 32'sd2103363, 32'sd2521603, -32'sd481896, -32'sd1284463, -32'sd1522585, 32'sd692633, 32'sd499764, 32'sd0, -32'sd835204, 32'sd283319, 32'sd869820, 32'sd487182, -32'sd138483, -32'sd1032920, 32'sd1313727, 32'sd294033, 32'sd1215079, 32'sd2564605, 32'sd1281618, 32'sd1114665, 32'sd1633873, -32'sd253122, -32'sd473318, 32'sd2111956, 32'sd2587530, 32'sd545840, -32'sd1599567, -32'sd498052, 32'sd1621556, 32'sd2743405, 32'sd2363315, 32'sd765771, 32'sd1061496, 32'sd1155323, -32'sd2421723, 32'sd203591, -32'sd574015, 32'sd1642977, -32'sd179225, -32'sd1323247, -32'sd3130218, -32'sd1750157, 32'sd477442, -32'sd678168, 32'sd37468, 32'sd440991, 32'sd2542198, 32'sd1733929, 32'sd1344274, -32'sd1346779, -32'sd2891026, -32'sd23719, 32'sd382737, 32'sd47849, -32'sd1383615, -32'sd442864, 32'sd1700292, 32'sd1724805, 32'sd1982086, 32'sd981411, -32'sd1837608, 32'sd579700, -32'sd1003952, -32'sd881415, -32'sd677531, 32'sd1452128, 32'sd150969, 32'sd94650, -32'sd296152, 32'sd479819, -32'sd367784, 32'sd1434672, 32'sd59303, 32'sd1069004, 32'sd2449538, 32'sd2442134, -32'sd1749036, -32'sd1460029, -32'sd786637, -32'sd281029, -32'sd854497, -32'sd23304, -32'sd97318, 32'sd1027774, 32'sd521256, 32'sd1283349, 32'sd2489637, -32'sd489945, -32'sd1331156, -32'sd2262604, 32'sd210090, 32'sd1119981, 32'sd1558960, -32'sd763371, 32'sd844132, 32'sd1905578, -32'sd582778, 32'sd601760, 32'sd855616, -32'sd254991, 32'sd804005, 32'sd882218, 32'sd1093864, 32'sd2345340, -32'sd928507, -32'sd866566, -32'sd2028590, -32'sd1433124, 32'sd769027, 32'sd1215146, 32'sd972973, 32'sd2247468, 32'sd635019, -32'sd485248, 32'sd83899, -32'sd668571, 32'sd422253, 32'sd227161, 32'sd439101, -32'sd582251, 32'sd448903, 32'sd321214, -32'sd61023, 32'sd2609349, 32'sd245247, 32'sd25155, -32'sd1110054, 32'sd1123005, 32'sd1430954, 32'sd1183133, 32'sd2782469, -32'sd273967, 32'sd893835, -32'sd544526, 32'sd224162, 32'sd293246, -32'sd801415, 32'sd1613178, 32'sd1312128, 32'sd819670, 32'sd616706, 32'sd1157356, 32'sd504407, 32'sd267513, 32'sd1643599, 32'sd731755, 32'sd452091, -32'sd653351, -32'sd193498, 32'sd1319326, 32'sd931640, 32'sd923938, 32'sd762419, -32'sd218646, 32'sd2795266, 32'sd3578827, 32'sd1619157, 32'sd593936, 32'sd2698834, 32'sd3414479, 32'sd976010, 32'sd11248, 32'sd2941112, 32'sd370771, -32'sd206390, -32'sd516229, 32'sd1592689, 32'sd2475835, 32'sd1318359, -32'sd412369, -32'sd166873, 32'sd210426, 32'sd37353, 32'sd931866, 32'sd768847, 32'sd40095, 32'sd415105, -32'sd162525, -32'sd751636, -32'sd602888, -32'sd945634, -32'sd1293702, 32'sd2621188, 32'sd2291177, 32'sd581026, 32'sd2825155, 32'sd2690114, 32'sd1951164, 32'sd1459498, -32'sd2081307, 32'sd1303052, -32'sd1007623, -32'sd552674, 32'sd165138, -32'sd220840, -32'sd839962, 32'sd142491, -32'sd216635, -32'sd1058366, -32'sd135644, 32'sd21711, -32'sd1217081, -32'sd1392804, -32'sd637673, -32'sd1049556, -32'sd671876, 32'sd104176, -32'sd302880, -32'sd53590, 32'sd2081521, 32'sd2423155, 32'sd529867, -32'sd573637, -32'sd1576090, -32'sd975602, -32'sd488761, -32'sd225159, -32'sd2071716, 32'sd967959, -32'sd770606, -32'sd1091081, 32'sd702063, -32'sd610269, -32'sd2112382, -32'sd504072, -32'sd1236491, 32'sd8898, 32'sd2650278, 32'sd1813426, 32'sd765609, -32'sd682465, -32'sd912459, 32'sd266672, -32'sd782512, 32'sd200335, 32'sd1629332, 32'sd285899, 32'sd2007970, 32'sd1273452, 32'sd1378319, 32'sd275307, -32'sd1397773, -32'sd1867375, 32'sd1163638, -32'sd848802, -32'sd1970108, -32'sd902795, -32'sd2656140, 32'sd606264, -32'sd267093, 32'sd47231, -32'sd2230698, -32'sd1962122, -32'sd1181514, -32'sd1470548, 32'sd8506, 32'sd283054, -32'sd2037344, 32'sd310085, 32'sd940110, 32'sd67342, -32'sd1742104, -32'sd788744, -32'sd115997, -32'sd411888, 32'sd1677117, 32'sd918135, -32'sd1099198, -32'sd1657882, 32'sd252262, -32'sd1896349, -32'sd2173345, -32'sd1992055, -32'sd1336406, 32'sd1234894, -32'sd1600422, -32'sd1237109, -32'sd433473, 32'sd222025, -32'sd1587489, -32'sd227388, -32'sd250648, -32'sd759911, -32'sd763182, -32'sd819466, 32'sd90858, 32'sd878548, 32'sd196975, -32'sd629005, -32'sd1161470, -32'sd1591273, -32'sd765175, 32'sd25177, -32'sd1605029, -32'sd805758, 32'sd747879, -32'sd2280182, -32'sd179476, -32'sd2764489, -32'sd2370034, -32'sd1371355, 32'sd166766, 32'sd1460451, -32'sd257591, 32'sd974818, -32'sd5114, -32'sd288664, -32'sd1015921, 32'sd446170, 32'sd1559695, 32'sd1209359, -32'sd328740, 32'sd1163418, -32'sd117234, -32'sd619220, 32'sd0, -32'sd76304, 32'sd48185, -32'sd2243945, -32'sd1642170, -32'sd1781182, -32'sd2337527, -32'sd1355228, -32'sd214999, -32'sd1833462, -32'sd88265, -32'sd820391, -32'sd2543593, -32'sd1200603, -32'sd2155217, 32'sd686511, -32'sd508611, -32'sd549121, -32'sd567360, -32'sd1412745, 32'sd363902, 32'sd1599863, 32'sd937670, -32'sd791873, 32'sd419005, 32'sd956512, 32'sd1695610, -32'sd52281, -32'sd736860, -32'sd153290, 32'sd146569, 32'sd605913, 32'sd154013, -32'sd3486322, -32'sd2157921, -32'sd2615188, -32'sd1103576, -32'sd2544721, -32'sd112031, -32'sd2694763, -32'sd1118977, 32'sd1130913, 32'sd47454, 32'sd361860, -32'sd17922, -32'sd1056990, -32'sd2253348, -32'sd2666516, -32'sd774485, 32'sd1274276, 32'sd626105, -32'sd439237, -32'sd2379411, -32'sd2166511, -32'sd368874, -32'sd766872, -32'sd807015, 32'sd132811, 32'sd649627, -32'sd1229477, 32'sd478037, -32'sd1970554, -32'sd2358562, -32'sd3297065, -32'sd1872370, -32'sd1671591, -32'sd2836067, -32'sd2913803, 32'sd1925265, 32'sd1054383, 32'sd1531016, -32'sd966321, -32'sd1810990, -32'sd1992784, -32'sd2323945, -32'sd3431400, -32'sd1982246, -32'sd26217, 32'sd16832, 32'sd1310400, -32'sd1331204, -32'sd1059162, 32'sd999754, -32'sd1462703, 32'sd0, 32'sd412429, 32'sd477042, -32'sd1133483, -32'sd2471383, -32'sd2940274, -32'sd2923462, -32'sd1788691, 32'sd24883, 32'sd865663, -32'sd1783567, 32'sd127567, 32'sd2346740, 32'sd963659, -32'sd1475306, -32'sd2415997, -32'sd2900989, -32'sd2718016, -32'sd2460156, -32'sd1892889, -32'sd755005, -32'sd441637, -32'sd1127137, 32'sd1232589, -32'sd658649, -32'sd158109, 32'sd13213, -32'sd131380, 32'sd1213, -32'sd245498, -32'sd1155348, -32'sd2017748, -32'sd511437, -32'sd2211418, -32'sd1335290, -32'sd2133186, -32'sd615657, -32'sd1061067, -32'sd1815137, 32'sd260216, 32'sd1112058, -32'sd610927, -32'sd604567, -32'sd1233964, -32'sd741617, -32'sd1238809, -32'sd2758078, -32'sd2013893, 32'sd401979, 32'sd1901479, 32'sd1468824, 32'sd56998, 32'sd66014, -32'sd155146, -32'sd766935, -32'sd284321, -32'sd127839, -32'sd2262371, 32'sd1117299, -32'sd923869, -32'sd435226, -32'sd2475244, 32'sd237866, 32'sd1325720, -32'sd1211305, 32'sd38995, 32'sd1134868, -32'sd168258, -32'sd147053, -32'sd396385, -32'sd827015, -32'sd90313, -32'sd1930765, -32'sd1587777, -32'sd1629494, -32'sd2088703, 32'sd55453, 32'sd86193, -32'sd1704287, -32'sd699695, -32'sd686832, 32'sd122856, -32'sd889394, -32'sd153162, 32'sd0, -32'sd334109, 32'sd950044, 32'sd1764418, 32'sd1605632, -32'sd1807835, 32'sd1409723, 32'sd1530675, 32'sd1214307, 32'sd1213638, -32'sd1301932, 32'sd1297471, -32'sd221592, -32'sd432670, 32'sd725633, -32'sd1543756, 32'sd109113, -32'sd933970, -32'sd3120000, -32'sd3684033, -32'sd220288, 32'sd1161064, -32'sd696287, -32'sd1226920, -32'sd1454884, 32'sd662426, -32'sd323612, 32'sd0, 32'sd0, 32'sd0, -32'sd1385998, -32'sd539540, -32'sd1162632, -32'sd1122713, 32'sd214888, -32'sd196390, 32'sd1493282, -32'sd691990, 32'sd1381561, 32'sd2302753, -32'sd664448, 32'sd1193630, 32'sd688276, 32'sd1624244, -32'sd431851, 32'sd277804, -32'sd1489771, -32'sd3855554, -32'sd1184054, -32'sd1468836, 32'sd2192203, -32'sd50615, 32'sd482446, -32'sd475953, -32'sd360274, 32'sd0, 32'sd0, 32'sd0, -32'sd753463, 32'sd682788, 32'sd278242, 32'sd102688, -32'sd1091491, 32'sd1278608, -32'sd358485, 32'sd180313, -32'sd90112, -32'sd514430, -32'sd1435901, -32'sd750749, 32'sd636348, 32'sd313586, 32'sd934255, 32'sd721406, -32'sd943642, -32'sd3137558, -32'sd2453315, -32'sd1585414, 32'sd985085, -32'sd21232, -32'sd387240, -32'sd775206, -32'sd664517, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd62187, -32'sd910506, -32'sd1063903, 32'sd89746, -32'sd1466651, 32'sd1276296, -32'sd155456, 32'sd1322190, -32'sd474591, 32'sd611498, 32'sd1048024, 32'sd363812, -32'sd2041999, -32'sd601906, 32'sd2013054, 32'sd997213, -32'sd1182503, 32'sd1012434, 32'sd244409, 32'sd503674, 32'sd643578, -32'sd2100975, 32'sd843894, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd696704, -32'sd511917, 32'sd166593, 32'sd252763, -32'sd859294, 32'sd800108, -32'sd459853, -32'sd985607, 32'sd172195, -32'sd1340265, 32'sd1186085, -32'sd22917, 32'sd144848, 32'sd1795524, 32'sd264039, -32'sd598780, -32'sd722082, 32'sd215286, 32'sd1279448, 32'sd1601429, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1359111, 32'sd1557097, -32'sd331106, -32'sd29936, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd336456, 32'sd9192, -32'sd168555, 32'sd455810, 32'sd242631, -32'sd86324, -32'sd448342, 32'sd1829869, -32'sd351174, -32'sd604886, 32'sd723389, -32'sd1244139, -32'sd1885789, 32'sd26373, -32'sd674161, 32'sd496761, 32'sd14240, -32'sd55122, -32'sd292723, -32'sd38628, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd314127, 32'sd379700, 32'sd1161636, 32'sd170949, 32'sd198309, -32'sd624672, 32'sd138893, -32'sd497446, -32'sd850044, -32'sd226120, 32'sd132067, -32'sd425035, -32'sd108042, -32'sd1148716, -32'sd1811, -32'sd1603993, -32'sd3018307, 32'sd306014, 32'sd1665500, -32'sd190842, 32'sd1691796, -32'sd524770, -32'sd222426, -32'sd82124, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd519962, -32'sd1505098, 32'sd372118, -32'sd1985564, -32'sd563636, -32'sd1558738, 32'sd687193, 32'sd581062, 32'sd73415, -32'sd44314, -32'sd202, 32'sd973641, 32'sd3336549, 32'sd1903517, 32'sd500609, -32'sd366658, 32'sd616895, -32'sd2206694, -32'sd2763594, -32'sd477805, -32'sd982277, -32'sd1947295, 32'sd34865, 32'sd735439, 32'sd258965, 32'sd0, 32'sd0, 32'sd1165350, 32'sd607558, 32'sd1303995, 32'sd502506, 32'sd626253, 32'sd174933, 32'sd606365, -32'sd2294386, -32'sd443371, -32'sd1378880, 32'sd450896, -32'sd433041, 32'sd74169, 32'sd639276, -32'sd1175470, 32'sd1959059, 32'sd388067, -32'sd123781, 32'sd455600, -32'sd1242818, -32'sd228719, -32'sd2066342, -32'sd1772172, -32'sd1776738, 32'sd837850, -32'sd1384911, 32'sd497457, 32'sd0, -32'sd700085, -32'sd632438, 32'sd1170210, -32'sd356040, -32'sd212801, -32'sd1286472, 32'sd992206, -32'sd2038580, 32'sd610618, 32'sd182148, 32'sd493078, 32'sd870144, 32'sd1708972, -32'sd509629, 32'sd800716, 32'sd525507, 32'sd1660409, -32'sd1711698, 32'sd962278, -32'sd201564, -32'sd2974427, -32'sd683815, 32'sd100985, -32'sd1466606, -32'sd1147232, 32'sd1102054, -32'sd540148, 32'sd0, 32'sd377854, -32'sd2204551, 32'sd93833, 32'sd201676, 32'sd134396, -32'sd446419, 32'sd1848494, 32'sd617111, 32'sd1879531, 32'sd1269362, 32'sd1678887, 32'sd2732131, 32'sd1383009, -32'sd163985, -32'sd1045431, 32'sd53170, 32'sd1416662, -32'sd227956, -32'sd2732926, -32'sd2879856, -32'sd2162933, -32'sd3341884, -32'sd1831178, -32'sd596058, -32'sd2331547, -32'sd1501201, 32'sd392493, -32'sd263665, 32'sd285613, -32'sd181049, -32'sd2567391, -32'sd617455, -32'sd2219925, -32'sd478491, -32'sd1104270, 32'sd127274, 32'sd551045, 32'sd1612285, 32'sd1665739, 32'sd80839, 32'sd1317953, 32'sd399516, -32'sd1063914, -32'sd622589, -32'sd1816272, -32'sd884557, -32'sd238142, -32'sd65691, -32'sd166077, -32'sd1266264, -32'sd549499, -32'sd3165019, -32'sd2737653, -32'sd685468, -32'sd481294, -32'sd297858, -32'sd1240086, 32'sd1695737, -32'sd458216, 32'sd734630, 32'sd424148, -32'sd689066, 32'sd169711, 32'sd3158044, 32'sd305651, -32'sd398785, 32'sd748040, 32'sd1018399, 32'sd316294, -32'sd1632776, -32'sd1085166, -32'sd171489, -32'sd1351106, 32'sd1484395, 32'sd937506, 32'sd209361, -32'sd801492, 32'sd556959, -32'sd1800782, -32'sd2967955, 32'sd244450, -32'sd1559860, 32'sd676186, -32'sd235069, -32'sd209679, 32'sd1871147, -32'sd696887, -32'sd112322, -32'sd359700, -32'sd232114, -32'sd311079, 32'sd744055, 32'sd859863, 32'sd1083511, -32'sd428735, -32'sd1330467, 32'sd110267, -32'sd1624982, 32'sd495940, -32'sd838984, 32'sd2861221, 32'sd821173, 32'sd1095468, 32'sd1667406, 32'sd731048, -32'sd310636, -32'sd1406058, -32'sd1245004, 32'sd446098, -32'sd144841, -32'sd492651, 32'sd1792648, 32'sd577548, -32'sd516175, -32'sd359185, 32'sd68640, -32'sd321631, 32'sd452159, 32'sd1056646, -32'sd141889, 32'sd24628, -32'sd2805212, -32'sd1257189, -32'sd1546584, -32'sd475890, 32'sd1191644, -32'sd1340493, -32'sd401711, 32'sd2777602, 32'sd1452005, 32'sd2518266, 32'sd1931296, 32'sd1031189, 32'sd1871903, -32'sd1541666, -32'sd71166, 32'sd814977, -32'sd1398065, 32'sd663875, 32'sd1111022, 32'sd216150, -32'sd2875316, -32'sd1758878, -32'sd215305, 32'sd488853, 32'sd410492, -32'sd726264, 32'sd2121083, 32'sd442454, -32'sd1913345, -32'sd2616059, 32'sd387160, 32'sd2837371, 32'sd2517717, 32'sd940449, -32'sd1148583, 32'sd2596753, 32'sd1421871, 32'sd2371373, 32'sd1506974, 32'sd27982, -32'sd551221, 32'sd369791, -32'sd1618726, 32'sd1173635, -32'sd990082, -32'sd93462, -32'sd310408, -32'sd309803, -32'sd1143951, -32'sd1846455, 32'sd99888, 32'sd203407, 32'sd771118, -32'sd787215, -32'sd275369, -32'sd2791067, -32'sd1830960, -32'sd275070, -32'sd631975, 32'sd2649015, 32'sd962249, 32'sd2215663, 32'sd465624, 32'sd1441283, 32'sd1219627, -32'sd881423, -32'sd311167, 32'sd586239, -32'sd1350501, 32'sd1442423, -32'sd1150777, -32'sd2129001, -32'sd475425, -32'sd949431, -32'sd312944, 32'sd761247, 32'sd435594, -32'sd1347821, -32'sd1083371, 32'sd235844, 32'sd1914109, 32'sd16974, -32'sd1133987, -32'sd1263908, -32'sd925107, 32'sd459369, 32'sd723271, 32'sd530112, 32'sd63626, -32'sd590925, -32'sd575380, -32'sd610650, -32'sd1008445, -32'sd1106977, -32'sd925329, -32'sd1103971, -32'sd224435, -32'sd2816864, -32'sd1222801, -32'sd824565, -32'sd1178968, 32'sd547853, 32'sd1158585, 32'sd474686, -32'sd1345103, -32'sd758252, 32'sd1022736, -32'sd1308781, -32'sd970456, -32'sd851944, -32'sd1177732, -32'sd55216, -32'sd728861, 32'sd2134754, 32'sd401778, 32'sd2631276, -32'sd1168569, 32'sd1726847, -32'sd595621, 32'sd845996, -32'sd643606, -32'sd1452838, 32'sd556111, -32'sd620477, 32'sd872104, -32'sd1004367, -32'sd3656084, -32'sd1943968, 32'sd567065, -32'sd635284, 32'sd829890, 32'sd340545, 32'sd559484, -32'sd452816, -32'sd1198337, -32'sd369485, -32'sd959867, -32'sd2486811, -32'sd1923456, -32'sd2019038, -32'sd212075, 32'sd36136, 32'sd1760378, 32'sd1280737, 32'sd2223016, 32'sd1224445, 32'sd28612, 32'sd2143017, 32'sd799499, -32'sd1049853, 32'sd219706, -32'sd802206, -32'sd1111488, -32'sd509617, -32'sd2418920, -32'sd592393, -32'sd936583, 32'sd221970, 32'sd890605, -32'sd969254, 32'sd698660, 32'sd491449, 32'sd349767, -32'sd328884, -32'sd2072301, -32'sd3271046, -32'sd3585444, -32'sd2246524, 32'sd2043098, -32'sd31538, -32'sd290762, -32'sd752472, -32'sd680099, -32'sd269585, 32'sd2336550, 32'sd2017946, 32'sd1323645, -32'sd1720704, -32'sd2160877, -32'sd4516920, -32'sd3086790, -32'sd2077876, -32'sd2459280, -32'sd1507148, -32'sd421129, 32'sd453203, 32'sd0, -32'sd60957, -32'sd384800, -32'sd712226, 32'sd837640, -32'sd327148, -32'sd1678907, -32'sd2567498, -32'sd3964123, -32'sd3743340, -32'sd3469425, -32'sd693690, -32'sd78957, 32'sd1704062, -32'sd1294547, -32'sd141200, 32'sd2000788, 32'sd2034290, -32'sd50047, -32'sd327065, -32'sd2288822, -32'sd922393, 32'sd52798, -32'sd512905, -32'sd157214, 32'sd859333, 32'sd926511, 32'sd351052, 32'sd308077, 32'sd762552, -32'sd595787, -32'sd541822, -32'sd221176, -32'sd1649236, 32'sd182275, -32'sd1923259, -32'sd2533068, -32'sd3299913, -32'sd2138693, -32'sd890176, 32'sd42726, -32'sd57778, -32'sd2696310, -32'sd2477951, 32'sd2876294, 32'sd1780229, 32'sd1243745, 32'sd397463, -32'sd3738428, -32'sd2367801, -32'sd1509363, -32'sd1570339, 32'sd411367, -32'sd23884, 32'sd670419, -32'sd642533, 32'sd560436, -32'sd879184, 32'sd535699, 32'sd752619, -32'sd1037466, 32'sd172275, 32'sd1411363, 32'sd847913, 32'sd942867, -32'sd365019, -32'sd2474301, -32'sd515630, -32'sd1100399, -32'sd3348489, -32'sd1648264, -32'sd453666, 32'sd1043987, 32'sd2089612, 32'sd1989657, 32'sd382446, -32'sd3596673, -32'sd2328158, -32'sd1382408, -32'sd1836544, -32'sd1340429, 32'sd1226911, -32'sd425688, 32'sd631932, 32'sd0, -32'sd1340323, -32'sd137269, -32'sd1850839, -32'sd613979, -32'sd249172, 32'sd1207917, 32'sd388475, -32'sd1424659, 32'sd454228, 32'sd305579, -32'sd1938524, -32'sd3176256, -32'sd2171937, -32'sd617634, -32'sd1020951, 32'sd25495, -32'sd313182, -32'sd862891, -32'sd1920989, -32'sd1835131, -32'sd2945510, -32'sd1041404, -32'sd2199693, -32'sd2979767, -32'sd175947, 32'sd1139056, -32'sd698543, 32'sd615626, 32'sd960821, -32'sd266703, -32'sd1164333, -32'sd582687, 32'sd587728, 32'sd1734382, -32'sd361838, -32'sd412890, -32'sd2615986, -32'sd987357, -32'sd2002441, -32'sd1300114, -32'sd3007067, -32'sd347183, -32'sd192810, 32'sd1081315, -32'sd296139, -32'sd499619, -32'sd4146534, -32'sd4574927, -32'sd3749717, -32'sd987493, -32'sd782699, 32'sd727973, -32'sd2239883, 32'sd33057, 32'sd1020248, 32'sd1248150, 32'sd651731, 32'sd346986, -32'sd412168, 32'sd715691, 32'sd799215, 32'sd1698362, 32'sd1613178, -32'sd1094426, -32'sd1716190, -32'sd324537, -32'sd823459, -32'sd815623, -32'sd2344695, 32'sd934106, -32'sd493772, -32'sd30215, -32'sd545994, -32'sd1310178, -32'sd1375087, -32'sd4188897, -32'sd4131596, -32'sd438552, -32'sd1560107, 32'sd1198742, -32'sd1445540, -32'sd1229560, 32'sd288415, 32'sd0, 32'sd995050, 32'sd1297920, 32'sd518467, 32'sd323063, 32'sd839185, -32'sd918366, 32'sd589195, -32'sd535164, -32'sd1191101, -32'sd93096, 32'sd1851901, 32'sd894635, -32'sd656528, 32'sd929899, -32'sd94155, -32'sd338860, -32'sd1155128, -32'sd282079, -32'sd256161, -32'sd3268360, -32'sd2858881, -32'sd1758314, 32'sd584562, -32'sd953546, -32'sd227956, -32'sd652559, 32'sd0, 32'sd0, 32'sd0, 32'sd1005219, 32'sd706526, -32'sd366223, 32'sd1733158, 32'sd1089873, 32'sd361580, 32'sd482898, 32'sd658833, -32'sd531268, -32'sd350606, -32'sd2023399, 32'sd599085, -32'sd239084, -32'sd389019, 32'sd2207553, -32'sd1050941, 32'sd935, -32'sd1571418, -32'sd2316869, -32'sd2836444, -32'sd2014721, -32'sd631676, 32'sd689952, 32'sd1879, 32'sd385036, 32'sd0, 32'sd0, 32'sd0, -32'sd433607, -32'sd526073, -32'sd43817, -32'sd1247671, -32'sd267268, -32'sd588115, -32'sd172457, -32'sd2336466, 32'sd1914916, -32'sd1107465, -32'sd1950412, -32'sd1237281, -32'sd1500022, -32'sd580260, -32'sd1480464, -32'sd748500, 32'sd1395179, 32'sd874505, -32'sd1548697, -32'sd509403, -32'sd3220305, -32'sd593953, 32'sd134544, 32'sd968651, -32'sd1418313, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd358298, -32'sd1728068, 32'sd890112, -32'sd284726, -32'sd1556924, -32'sd1528657, -32'sd1680529, 32'sd617174, -32'sd948650, -32'sd1483749, 32'sd111344, 32'sd787838, -32'sd18121, 32'sd1765831, 32'sd1705531, 32'sd2516774, 32'sd730042, 32'sd1711520, 32'sd2627423, -32'sd1687478, 32'sd281196, 32'sd1168543, 32'sd427202, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd268159, 32'sd893505, -32'sd1114540, 32'sd1159390, -32'sd18663, -32'sd913435, -32'sd2147853, 32'sd558279, -32'sd430604, -32'sd1126292, -32'sd643256, 32'sd1000340, 32'sd1323198, 32'sd734910, -32'sd343131, -32'sd332307, -32'sd1911133, -32'sd648144, 32'sd371411, 32'sd99972, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd330022, 32'sd2098168, 32'sd1252969, 32'sd1009068, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd286893, 32'sd1048490, 32'sd317423, 32'sd1896279, 32'sd1444002, 32'sd1258082, 32'sd1597858, 32'sd1236983, 32'sd839553, 32'sd542982, 32'sd842948, 32'sd510295, 32'sd1198733, 32'sd287426, 32'sd675963, -32'sd281444, 32'sd657401, -32'sd148473, 32'sd516240, 32'sd269666, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1734217, -32'sd39875, -32'sd17136, 32'sd1159977, 32'sd1135365, -32'sd398349, -32'sd209273, 32'sd57485, 32'sd380532, -32'sd205017, 32'sd165047, -32'sd2742309, -32'sd1073644, -32'sd788618, 32'sd19798, 32'sd889727, 32'sd661298, 32'sd385436, 32'sd315375, 32'sd1958688, 32'sd1696723, 32'sd956613, 32'sd1552461, 32'sd1201389, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1297023, -32'sd23792, -32'sd57218, -32'sd625428, -32'sd127801, -32'sd1018075, -32'sd1410432, 32'sd1063379, -32'sd460290, -32'sd342757, 32'sd1449426, -32'sd175605, -32'sd326119, -32'sd1042514, -32'sd771991, -32'sd2421598, -32'sd1625037, 32'sd788421, 32'sd627147, 32'sd2077531, -32'sd286182, -32'sd107356, 32'sd1462102, 32'sd939441, -32'sd362550, 32'sd0, 32'sd0, 32'sd216574, -32'sd1359102, 32'sd430618, 32'sd1175731, -32'sd149097, 32'sd1763830, 32'sd510714, -32'sd99339, -32'sd1248074, -32'sd1040204, -32'sd282166, -32'sd1459461, -32'sd97694, 32'sd39309, -32'sd930592, 32'sd727552, 32'sd1240354, 32'sd2211131, 32'sd1796603, 32'sd1887713, 32'sd2274793, -32'sd660521, 32'sd155600, 32'sd2261356, -32'sd708442, 32'sd666903, 32'sd429219, 32'sd0, -32'sd202126, 32'sd2362786, -32'sd829971, -32'sd326426, 32'sd600526, -32'sd1031472, -32'sd680654, 32'sd329800, -32'sd299040, 32'sd1628711, 32'sd1275789, -32'sd831143, -32'sd1227082, -32'sd1637123, 32'sd731856, -32'sd894699, 32'sd1807405, -32'sd466494, 32'sd316123, 32'sd687985, 32'sd2089318, 32'sd1903277, -32'sd164324, 32'sd1409843, 32'sd425390, -32'sd166702, 32'sd304449, 32'sd0, 32'sd420424, 32'sd514056, -32'sd950979, 32'sd399806, 32'sd726219, -32'sd447320, -32'sd1135699, 32'sd146220, 32'sd483302, -32'sd210558, -32'sd436312, -32'sd567968, -32'sd413357, -32'sd609772, -32'sd1347482, 32'sd510463, 32'sd248639, 32'sd122771, -32'sd66745, 32'sd1175959, 32'sd417079, 32'sd192334, 32'sd12928, 32'sd1284891, 32'sd784873, 32'sd536887, -32'sd985410, 32'sd947976, -32'sd976640, 32'sd205696, 32'sd1147337, 32'sd393290, -32'sd23557, 32'sd99443, 32'sd188358, 32'sd1990545, -32'sd1488886, -32'sd62306, -32'sd1963996, -32'sd1140235, 32'sd1380182, -32'sd674288, 32'sd649087, -32'sd664962, -32'sd444922, 32'sd37711, -32'sd167659, -32'sd569715, -32'sd1032430, 32'sd2104204, -32'sd1474699, 32'sd68197, -32'sd347758, 32'sd1245290, 32'sd482589, 32'sd188168, 32'sd1218340, 32'sd716829, 32'sd1406053, 32'sd2881558, 32'sd1035221, -32'sd1430500, -32'sd157244, 32'sd830062, -32'sd758100, 32'sd794075, 32'sd787365, 32'sd324287, 32'sd1631435, 32'sd1159080, 32'sd95986, 32'sd757529, -32'sd2035024, -32'sd734861, 32'sd806033, 32'sd234976, -32'sd1587324, -32'sd1317910, 32'sd687866, 32'sd591508, -32'sd1119219, 32'sd505430, 32'sd365139, 32'sd621244, 32'sd435829, 32'sd111316, 32'sd1396216, 32'sd898688, -32'sd411663, -32'sd830073, 32'sd1085168, 32'sd1221849, 32'sd624009, 32'sd3333345, 32'sd763804, 32'sd2953275, 32'sd2835898, 32'sd2650262, 32'sd174891, 32'sd1829653, 32'sd1002766, 32'sd569096, 32'sd258802, 32'sd561902, -32'sd106607, -32'sd444667, 32'sd1994472, 32'sd736998, 32'sd83381, 32'sd2314653, 32'sd1238686, -32'sd863035, 32'sd365168, 32'sd1997619, 32'sd2662532, -32'sd257544, -32'sd294564, 32'sd1230572, 32'sd1351146, 32'sd943210, 32'sd1673653, 32'sd3515550, 32'sd3125270, 32'sd210524, -32'sd655908, -32'sd2177055, 32'sd315796, 32'sd5704, -32'sd1519588, 32'sd21987, -32'sd739709, 32'sd1638153, -32'sd24904, -32'sd1090649, 32'sd180605, -32'sd803021, 32'sd1204707, 32'sd2829719, -32'sd642082, 32'sd1116570, -32'sd576466, 32'sd1139262, 32'sd875645, -32'sd668978, 32'sd2257950, 32'sd1265992, 32'sd2279902, -32'sd874563, 32'sd2763991, 32'sd1172463, 32'sd1290901, -32'sd1497201, -32'sd4916624, -32'sd4194267, -32'sd385112, 32'sd2365876, -32'sd791028, -32'sd661765, 32'sd729611, -32'sd148690, 32'sd694288, -32'sd471241, -32'sd126300, -32'sd968486, 32'sd1279640, 32'sd1070971, 32'sd880712, 32'sd244361, -32'sd732022, 32'sd1096139, 32'sd1319208, 32'sd877228, 32'sd1466398, 32'sd926115, 32'sd2205826, -32'sd467421, -32'sd670655, -32'sd2677180, -32'sd1725660, -32'sd1294839, -32'sd4507566, -32'sd4931330, -32'sd2058139, -32'sd1101271, -32'sd140842, 32'sd426965, 32'sd964, 32'sd984824, -32'sd844529, -32'sd616846, -32'sd1330247, 32'sd1028149, 32'sd718283, -32'sd641195, -32'sd1046863, 32'sd996947, 32'sd802498, 32'sd321539, 32'sd349020, 32'sd271066, -32'sd1366356, -32'sd286714, -32'sd957948, -32'sd758489, -32'sd99166, -32'sd3277849, -32'sd2433022, -32'sd2009909, -32'sd2521702, -32'sd1928732, -32'sd1200464, -32'sd3225522, -32'sd385224, -32'sd1152423, 32'sd170511, -32'sd1049164, -32'sd460441, -32'sd1328966, 32'sd819087, 32'sd1596779, -32'sd812726, 32'sd1371482, 32'sd59562, 32'sd212568, -32'sd17216, 32'sd1372433, 32'sd128720, -32'sd57784, -32'sd748036, -32'sd2241109, -32'sd3280196, -32'sd5573111, -32'sd3945598, -32'sd1943139, -32'sd2724962, -32'sd3174096, -32'sd72635, -32'sd1777878, -32'sd1309102, -32'sd3768408, -32'sd1474646, -32'sd1796174, -32'sd915474, 32'sd662874, -32'sd673433, -32'sd736911, -32'sd1163810, -32'sd130660, -32'sd1017297, 32'sd111105, 32'sd192248, 32'sd774648, -32'sd463545, 32'sd685588, -32'sd1444588, -32'sd2352792, -32'sd2868549, -32'sd3731559, -32'sd2886156, -32'sd4616313, -32'sd3369676, -32'sd2127086, -32'sd2962873, -32'sd1412305, 32'sd1921066, -32'sd18464, -32'sd2568306, -32'sd2926050, -32'sd1903892, -32'sd1758113, -32'sd700060, -32'sd2160644, -32'sd2375743, -32'sd624184, -32'sd83544, 32'sd1068119, -32'sd260880, -32'sd319539, 32'sd629254, 32'sd1009692, 32'sd495897, 32'sd587683, -32'sd2182155, -32'sd3321267, -32'sd4159411, -32'sd4307180, -32'sd2610154, -32'sd2972545, -32'sd914658, -32'sd2012081, -32'sd179181, 32'sd1786486, 32'sd622650, 32'sd2800734, -32'sd197907, -32'sd112685, -32'sd1111573, -32'sd563438, -32'sd645414, -32'sd3759203, 32'sd37188, 32'sd1222173, 32'sd418752, -32'sd538535, 32'sd1387018, -32'sd275790, 32'sd1404969, 32'sd0, 32'sd1105443, -32'sd150035, -32'sd1534299, -32'sd298227, -32'sd1254423, -32'sd2187213, -32'sd2066260, -32'sd1075562, 32'sd1401179, 32'sd2312004, 32'sd1347736, 32'sd1923357, 32'sd2657369, 32'sd1132898, -32'sd906326, -32'sd217369, -32'sd1936006, -32'sd1582468, -32'sd1437705, -32'sd2466452, 32'sd918, -32'sd187648, 32'sd662122, 32'sd1930367, 32'sd3070525, -32'sd386601, 32'sd772041, 32'sd574404, -32'sd647116, 32'sd1521534, 32'sd499823, 32'sd1410921, -32'sd1468872, 32'sd446366, -32'sd1977032, 32'sd862053, 32'sd1132815, 32'sd3579413, -32'sd218230, 32'sd643341, 32'sd1695554, 32'sd912432, 32'sd2312296, -32'sd328052, -32'sd1026615, -32'sd848995, -32'sd104056, 32'sd187808, 32'sd727730, -32'sd636492, -32'sd2348922, -32'sd440676, 32'sd401647, 32'sd1818246, 32'sd199330, 32'sd782291, -32'sd911616, 32'sd210479, -32'sd98837, 32'sd1506450, -32'sd226964, -32'sd1473230, 32'sd1891598, 32'sd2955046, 32'sd2459239, 32'sd380196, 32'sd442779, 32'sd652934, 32'sd657970, 32'sd825244, 32'sd1540535, 32'sd2826219, 32'sd2581335, 32'sd1337872, 32'sd48695, 32'sd1343996, -32'sd787577, -32'sd565391, -32'sd518100, 32'sd1660536, 32'sd1760517, 32'sd1478034, 32'sd214064, 32'sd0, -32'sd68813, 32'sd180924, 32'sd772142, 32'sd32497, -32'sd418400, 32'sd962857, 32'sd1582054, 32'sd3445255, 32'sd1814322, 32'sd935700, -32'sd130836, 32'sd1490595, 32'sd2120465, 32'sd1842879, 32'sd2760754, 32'sd525439, 32'sd2758953, 32'sd169284, 32'sd1461506, -32'sd736794, 32'sd724126, -32'sd1782727, -32'sd916637, 32'sd460606, 32'sd320636, 32'sd1358036, 32'sd255081, 32'sd1106865, 32'sd709400, 32'sd171577, 32'sd2648924, 32'sd1313648, 32'sd2226543, 32'sd1999447, 32'sd776027, 32'sd520329, 32'sd1000007, 32'sd563937, 32'sd857900, -32'sd199397, 32'sd2095515, 32'sd1698584, 32'sd2661109, 32'sd2209182, 32'sd2514790, 32'sd2285258, 32'sd2239765, 32'sd305036, -32'sd1040346, -32'sd878197, 32'sd928361, 32'sd1764225, 32'sd1065339, 32'sd1880588, -32'sd987443, 32'sd73460, -32'sd225877, 32'sd491872, 32'sd715291, 32'sd1676191, 32'sd59848, 32'sd884951, 32'sd1374498, 32'sd573311, 32'sd404313, 32'sd582069, 32'sd799242, -32'sd866148, 32'sd1905522, -32'sd769776, 32'sd2473357, 32'sd1718633, 32'sd2588704, 32'sd1312319, 32'sd313593, -32'sd143013, -32'sd597232, -32'sd644183, 32'sd683172, -32'sd560482, 32'sd969376, 32'sd1216739, 32'sd697402, 32'sd0, 32'sd452274, 32'sd945358, 32'sd1071115, -32'sd85271, 32'sd1297017, 32'sd1590442, 32'sd700767, 32'sd1836364, 32'sd1424561, 32'sd1427871, -32'sd292325, 32'sd1958103, 32'sd1859979, -32'sd364605, 32'sd753068, 32'sd1901846, 32'sd326702, 32'sd868420, 32'sd318387, 32'sd1704035, -32'sd1085897, -32'sd585216, 32'sd837545, -32'sd788625, -32'sd1083609, -32'sd327018, 32'sd0, 32'sd0, 32'sd0, 32'sd262652, -32'sd1076421, 32'sd1412907, 32'sd439761, 32'sd765352, 32'sd655284, 32'sd1099723, 32'sd1473173, 32'sd1062668, 32'sd1078946, 32'sd116478, 32'sd1331812, -32'sd484851, 32'sd1161244, 32'sd1188974, 32'sd1070785, 32'sd1454472, 32'sd2453867, 32'sd1868076, -32'sd151458, 32'sd303207, -32'sd313649, 32'sd1281203, 32'sd550880, -32'sd1304267, 32'sd0, 32'sd0, 32'sd0, -32'sd1293993, -32'sd460739, -32'sd1123391, 32'sd926960, -32'sd60404, -32'sd5431, 32'sd788819, 32'sd1404457, -32'sd98270, 32'sd204671, 32'sd1399141, 32'sd1525001, 32'sd201999, -32'sd923681, 32'sd723038, 32'sd772001, 32'sd778583, 32'sd755148, -32'sd35810, 32'sd647178, -32'sd535569, -32'sd1393929, 32'sd637771, 32'sd101328, 32'sd578408, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd400980, -32'sd1371204, -32'sd303211, -32'sd258682, 32'sd1993730, 32'sd1662428, 32'sd780502, -32'sd690567, 32'sd475576, -32'sd997472, 32'sd1482610, 32'sd368967, 32'sd1261294, -32'sd37676, 32'sd643218, 32'sd165631, 32'sd1418060, -32'sd12568, -32'sd686182, 32'sd81626, -32'sd1620951, 32'sd976000, 32'sd373387, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1170613, 32'sd855750, 32'sd821088, -32'sd503455, -32'sd481015, 32'sd721683, 32'sd1700751, -32'sd171644, -32'sd955139, 32'sd2038436, 32'sd1193566, -32'sd604492, 32'sd1535371, 32'sd1566683, -32'sd117010, -32'sd1058784, 32'sd1457615, -32'sd912218, -32'sd146606, 32'sd584359, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1372774, 32'sd507677, 32'sd295159, -32'sd248529, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd295104, -32'sd677348, -32'sd614003, -32'sd1259137, 32'sd758222, -32'sd367307, -32'sd891494, 32'sd557312, 32'sd601828, -32'sd525912, -32'sd677212, 32'sd1035453, -32'sd920334, 32'sd2898, 32'sd833628, -32'sd251771, 32'sd449921, 32'sd1338996, -32'sd67066, 32'sd54485, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd183480, -32'sd308689, -32'sd297490, 32'sd99605, -32'sd96585, 32'sd233443, 32'sd817553, -32'sd318414, -32'sd1445183, -32'sd47879, 32'sd1526313, -32'sd658661, -32'sd1660129, -32'sd3275673, -32'sd2124880, -32'sd595467, -32'sd2263657, -32'sd1585929, -32'sd50693, -32'sd81959, -32'sd447110, 32'sd420047, 32'sd89004, -32'sd64024, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd276535, -32'sd36388, -32'sd754708, -32'sd2094686, -32'sd1440744, -32'sd766600, -32'sd1187121, 32'sd139854, 32'sd312690, 32'sd82572, -32'sd1226907, 32'sd760872, 32'sd1710238, 32'sd985742, -32'sd815979, 32'sd1145251, 32'sd1334559, 32'sd2490822, 32'sd1513627, -32'sd508499, 32'sd1416591, -32'sd510480, -32'sd562121, 32'sd965640, 32'sd1220938, 32'sd0, 32'sd0, -32'sd179039, -32'sd923312, 32'sd1152873, 32'sd965904, 32'sd807613, -32'sd245814, 32'sd241635, -32'sd1122528, -32'sd368596, -32'sd2693018, -32'sd409423, -32'sd1165030, 32'sd2876720, 32'sd1324577, 32'sd751503, 32'sd859886, 32'sd1777667, 32'sd1523531, 32'sd174823, 32'sd1211587, 32'sd942695, 32'sd743190, 32'sd723089, -32'sd1226208, -32'sd1831678, 32'sd1347346, -32'sd166842, 32'sd0, 32'sd995572, -32'sd367895, 32'sd644389, -32'sd2866125, -32'sd818957, -32'sd396884, -32'sd2253849, -32'sd1086353, 32'sd179089, -32'sd1727173, -32'sd3644455, -32'sd2228832, -32'sd482526, 32'sd512084, 32'sd1904817, 32'sd2300246, 32'sd66673, 32'sd1972525, 32'sd1301089, -32'sd621697, 32'sd1379205, 32'sd363813, -32'sd139585, -32'sd2175456, -32'sd1327278, 32'sd1351366, 32'sd1203754, 32'sd0, -32'sd122980, 32'sd610039, 32'sd586098, -32'sd261979, -32'sd1447888, -32'sd732815, -32'sd1159073, 32'sd796864, -32'sd786741, 32'sd42135, -32'sd1240896, -32'sd1528207, -32'sd913395, 32'sd532813, -32'sd515051, 32'sd894974, 32'sd1234732, 32'sd794277, 32'sd328494, -32'sd706264, -32'sd279422, 32'sd1116240, -32'sd961066, 32'sd100, -32'sd146998, 32'sd308753, 32'sd1586359, -32'sd306503, -32'sd521557, 32'sd1939248, 32'sd430588, -32'sd321247, 32'sd847448, 32'sd1636849, 32'sd655084, 32'sd725109, 32'sd1603635, -32'sd26201, -32'sd143824, -32'sd49195, -32'sd1125606, -32'sd49530, -32'sd1207004, 32'sd1760857, -32'sd807519, 32'sd279792, 32'sd2675601, 32'sd2740285, 32'sd1550377, 32'sd313277, 32'sd1615086, -32'sd71817, 32'sd5797, 32'sd176365, 32'sd1120125, -32'sd31144, 32'sd470875, 32'sd908229, -32'sd1640482, -32'sd315191, -32'sd177723, 32'sd1605050, 32'sd1317146, 32'sd1238083, 32'sd768404, 32'sd430194, -32'sd1798142, -32'sd1924224, -32'sd1061921, 32'sd452276, 32'sd2329134, 32'sd1468121, -32'sd1621227, -32'sd1560248, 32'sd1296807, 32'sd1169968, 32'sd522117, -32'sd125876, 32'sd658199, -32'sd811832, 32'sd666219, -32'sd1446489, 32'sd646270, 32'sd335120, -32'sd795175, -32'sd44430, 32'sd994174, 32'sd2041256, 32'sd470285, -32'sd1482921, -32'sd984768, 32'sd593677, 32'sd384224, -32'sd928583, -32'sd3113436, -32'sd3777856, 32'sd579203, 32'sd2228810, 32'sd1617144, -32'sd929129, -32'sd1884935, -32'sd706525, 32'sd1763550, 32'sd2159113, 32'sd614129, 32'sd756360, 32'sd1293293, -32'sd1272258, 32'sd1689214, -32'sd839448, 32'sd1281470, -32'sd1053135, -32'sd1570158, 32'sd1056639, -32'sd873170, -32'sd50268, -32'sd1236057, -32'sd1082076, -32'sd972836, -32'sd313438, 32'sd375745, -32'sd1555815, -32'sd2759044, -32'sd2277050, 32'sd2441826, 32'sd2254484, 32'sd1580373, 32'sd811906, 32'sd550148, -32'sd121432, 32'sd573565, 32'sd1931363, 32'sd185506, 32'sd3256928, 32'sd1791293, -32'sd1146897, 32'sd556040, -32'sd236920, -32'sd861044, 32'sd1033085, -32'sd908258, -32'sd619070, 32'sd1339219, -32'sd2673120, -32'sd1334505, -32'sd1627536, -32'sd902402, 32'sd396494, 32'sd450825, -32'sd2273370, -32'sd2393398, -32'sd2638360, -32'sd384644, 32'sd713689, 32'sd1458040, 32'sd178746, 32'sd620795, 32'sd1091538, -32'sd31892, 32'sd1026944, -32'sd25611, 32'sd2533921, -32'sd1448279, 32'sd65767, -32'sd1185558, 32'sd414986, 32'sd1137675, 32'sd574788, 32'sd849681, 32'sd427970, -32'sd1573430, -32'sd412524, -32'sd894589, 32'sd448407, -32'sd1052356, -32'sd97582, 32'sd75925, -32'sd3844814, -32'sd1427669, -32'sd2222773, -32'sd390375, 32'sd818210, 32'sd1140615, 32'sd1823710, -32'sd762212, -32'sd1173040, -32'sd1099218, 32'sd212787, -32'sd32920, 32'sd414344, -32'sd243871, 32'sd79844, -32'sd926126, -32'sd699236, 32'sd349760, -32'sd283659, -32'sd528250, -32'sd431777, 32'sd1130532, 32'sd15319, -32'sd91211, -32'sd1036333, 32'sd674499, -32'sd171325, -32'sd700680, -32'sd681650, -32'sd3794052, -32'sd2848007, 32'sd822333, 32'sd1706939, 32'sd1266388, 32'sd788161, 32'sd26861, 32'sd132546, 32'sd927266, 32'sd128886, 32'sd193437, 32'sd300086, 32'sd1828482, -32'sd876534, -32'sd1044315, -32'sd763131, -32'sd116684, -32'sd263249, 32'sd948395, -32'sd806698, -32'sd240208, -32'sd221298, 32'sd1512858, 32'sd815418, 32'sd1210375, 32'sd2357397, -32'sd1020515, -32'sd1754321, -32'sd1419466, -32'sd240386, -32'sd691532, 32'sd1022378, -32'sd825872, 32'sd91569, 32'sd759010, 32'sd1029153, 32'sd1129066, 32'sd2837225, 32'sd4143231, 32'sd2156793, 32'sd709764, 32'sd977002, -32'sd1587804, -32'sd732430, -32'sd542677, -32'sd252534, 32'sd533243, -32'sd439139, -32'sd986074, 32'sd598329, 32'sd1854317, 32'sd631573, 32'sd797711, -32'sd202228, -32'sd877035, -32'sd2992143, -32'sd920238, 32'sd689803, -32'sd229262, -32'sd130360, -32'sd1598412, 32'sd746885, 32'sd629560, -32'sd584810, -32'sd638998, 32'sd1721023, 32'sd522010, -32'sd87209, 32'sd738981, 32'sd522158, -32'sd3013828, 32'sd545039, -32'sd329555, -32'sd309596, 32'sd1502389, 32'sd404586, 32'sd1218217, -32'sd359438, 32'sd1101365, 32'sd1402441, 32'sd259784, 32'sd754780, -32'sd1358049, -32'sd2184462, -32'sd2435407, -32'sd27872, 32'sd674063, -32'sd657785, -32'sd472866, -32'sd1055670, -32'sd1038722, 32'sd125859, -32'sd1540484, 32'sd1617044, -32'sd71582, 32'sd660815, -32'sd1057725, 32'sd1422038, 32'sd82135, -32'sd1400678, -32'sd457755, 32'sd0, 32'sd1941735, 32'sd2324749, -32'sd580012, 32'sd1191675, 32'sd2057555, -32'sd517596, 32'sd1331064, 32'sd420496, -32'sd2051926, -32'sd3276308, -32'sd1847340, -32'sd573561, -32'sd1278374, -32'sd1589667, -32'sd338561, 32'sd499100, 32'sd912518, 32'sd441508, 32'sd43894, 32'sd239637, -32'sd951027, -32'sd532397, 32'sd949137, -32'sd1227795, -32'sd496643, 32'sd345421, -32'sd313166, 32'sd372342, -32'sd4383, 32'sd894867, -32'sd224937, -32'sd47243, 32'sd527088, 32'sd1280556, 32'sd1901767, 32'sd1896589, 32'sd1980964, 32'sd393037, -32'sd1236106, -32'sd1853401, 32'sd153832, -32'sd87946, 32'sd331792, -32'sd321471, -32'sd2804, 32'sd202450, -32'sd976665, -32'sd158042, -32'sd290559, 32'sd601281, 32'sd311057, -32'sd1538869, -32'sd1610226, 32'sd243335, -32'sd183923, 32'sd332428, 32'sd347327, -32'sd1551827, 32'sd580594, 32'sd1962383, 32'sd1669359, 32'sd2628116, 32'sd3138669, 32'sd1871744, 32'sd3605162, 32'sd1753372, -32'sd643704, 32'sd2393475, 32'sd151669, -32'sd25249, 32'sd1439690, -32'sd2558592, -32'sd1637491, -32'sd238070, 32'sd299727, 32'sd56934, -32'sd1587732, -32'sd774172, -32'sd136029, -32'sd581148, -32'sd970424, -32'sd460047, -32'sd154752, 32'sd0, 32'sd78228, -32'sd46140, 32'sd2202889, 32'sd1975101, 32'sd139811, 32'sd778206, 32'sd866834, 32'sd2283110, 32'sd2680843, 32'sd1899321, 32'sd891551, 32'sd1768497, 32'sd2626980, 32'sd50756, -32'sd2588841, -32'sd1401954, -32'sd2853587, -32'sd3041715, -32'sd1752893, 32'sd164811, 32'sd546886, -32'sd401286, -32'sd1768177, 32'sd414827, 32'sd1395287, -32'sd148060, 32'sd2035974, -32'sd392527, 32'sd817379, 32'sd71584, 32'sd637715, 32'sd1579184, -32'sd1703699, -32'sd402808, 32'sd1179129, 32'sd3079107, 32'sd3318717, 32'sd3343439, 32'sd3715363, 32'sd2478503, 32'sd1248097, 32'sd582744, -32'sd1385156, -32'sd904841, 32'sd645871, -32'sd1442121, 32'sd9763, 32'sd654453, -32'sd183305, -32'sd1941868, -32'sd1982728, -32'sd1404368, -32'sd535527, 32'sd1901272, 32'sd786851, -32'sd960405, 32'sd469017, 32'sd1608228, 32'sd1355916, 32'sd1502288, 32'sd325792, 32'sd362416, 32'sd227948, 32'sd2265804, 32'sd2498548, 32'sd4942884, 32'sd2124356, 32'sd3287936, 32'sd3346999, 32'sd1543147, 32'sd701178, 32'sd1571891, -32'sd8082, -32'sd1032203, 32'sd982119, 32'sd385540, 32'sd281601, 32'sd40714, -32'sd2235400, 32'sd455200, -32'sd69331, 32'sd494536, 32'sd1311949, 32'sd0, 32'sd768673, 32'sd1993913, 32'sd368203, -32'sd339364, 32'sd702309, 32'sd1808435, -32'sd318856, -32'sd909948, 32'sd1727196, 32'sd3027183, 32'sd3044641, 32'sd1235392, 32'sd1023795, 32'sd208825, -32'sd23762, 32'sd1021334, 32'sd1448140, -32'sd974028, -32'sd3745019, -32'sd2555902, -32'sd66556, -32'sd839924, -32'sd157323, -32'sd650763, -32'sd842300, -32'sd689372, 32'sd0, 32'sd0, 32'sd0, 32'sd260524, 32'sd1630770, 32'sd1824258, 32'sd547323, 32'sd1579150, 32'sd281478, 32'sd1889029, -32'sd1461637, -32'sd1706976, -32'sd3473180, -32'sd2124286, -32'sd1472824, -32'sd99812, 32'sd963607, -32'sd1569209, -32'sd1003305, -32'sd1369073, -32'sd2947793, 32'sd37071, -32'sd346292, 32'sd216579, -32'sd533206, 32'sd890152, 32'sd1087986, 32'sd1481199, 32'sd0, 32'sd0, 32'sd0, 32'sd1398174, -32'sd239636, 32'sd383615, -32'sd407268, -32'sd2298969, -32'sd2106101, 32'sd835775, 32'sd974817, -32'sd2126602, -32'sd2631066, -32'sd3692357, -32'sd1397765, -32'sd1165533, -32'sd980742, -32'sd1862601, -32'sd3224943, -32'sd1227951, -32'sd66340, -32'sd366194, -32'sd1176099, 32'sd435846, -32'sd116583, 32'sd1621567, -32'sd728137, 32'sd753907, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd268980, -32'sd873787, -32'sd1818170, -32'sd1154600, -32'sd580188, -32'sd2326606, -32'sd1598178, -32'sd552497, -32'sd688839, 32'sd1013474, -32'sd1097235, -32'sd767914, -32'sd1871102, -32'sd1515963, -32'sd666854, -32'sd1048895, -32'sd323707, -32'sd1351650, 32'sd150007, 32'sd505022, -32'sd1030492, 32'sd368597, 32'sd127462, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd562991, -32'sd621516, -32'sd328498, 32'sd149679, 32'sd589890, -32'sd310569, -32'sd648721, 32'sd143256, 32'sd1526204, 32'sd1278696, -32'sd685286, -32'sd912261, -32'sd1129017, -32'sd274971, 32'sd168396, 32'sd790632, 32'sd745914, -32'sd893658, 32'sd142077, -32'sd316570, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd879372, 32'sd887935, -32'sd218752, 32'sd1589868, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd140275, 32'sd452198, -32'sd461834, 32'sd858937, -32'sd1246048, 32'sd116584, -32'sd663102, -32'sd266130, -32'sd1013656, -32'sd957932, -32'sd450336, 32'sd1107870, -32'sd381770, 32'sd448580, -32'sd398607, -32'sd7760, 32'sd863091, 32'sd120513, 32'sd11379, 32'sd159295, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd827715, -32'sd33960, -32'sd1049025, -32'sd162370, -32'sd920105, 32'sd42243, -32'sd355687, -32'sd1684996, -32'sd348875, 32'sd8817, -32'sd1647823, -32'sd1879678, -32'sd1392856, -32'sd490853, -32'sd642226, -32'sd51657, -32'sd421395, -32'sd634028, -32'sd1380840, 32'sd504425, 32'sd804863, 32'sd696779, 32'sd1042745, -32'sd592057, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd591013, -32'sd59820, 32'sd633866, 32'sd1280600, -32'sd311806, -32'sd944099, -32'sd2248420, -32'sd710056, 32'sd752523, 32'sd816694, 32'sd1928458, 32'sd326873, -32'sd595204, -32'sd2241574, 32'sd488703, -32'sd469075, -32'sd2752601, -32'sd3800486, -32'sd2494254, -32'sd1115247, -32'sd1339659, -32'sd943875, 32'sd1124441, 32'sd476037, -32'sd1012493, 32'sd0, 32'sd0, -32'sd186973, 32'sd181184, 32'sd1160732, -32'sd1024890, 32'sd541741, 32'sd946139, 32'sd1361125, 32'sd213735, 32'sd636869, -32'sd344712, 32'sd936265, -32'sd971659, 32'sd322276, 32'sd443887, -32'sd355184, -32'sd203881, 32'sd393223, -32'sd566695, -32'sd2322567, -32'sd1044730, -32'sd1611844, -32'sd1214268, -32'sd1474435, 32'sd610703, -32'sd433715, -32'sd408932, 32'sd604045, 32'sd0, 32'sd372216, -32'sd296260, -32'sd1844138, -32'sd2565668, -32'sd505276, -32'sd613398, -32'sd1002781, -32'sd114079, 32'sd1825019, 32'sd1098629, 32'sd601142, 32'sd1367858, -32'sd91692, 32'sd66658, -32'sd396791, 32'sd2486, -32'sd75441, 32'sd2694408, 32'sd888873, -32'sd1038635, -32'sd1113957, -32'sd58557, -32'sd333669, -32'sd383414, -32'sd769006, 32'sd1541681, 32'sd414632, 32'sd0, 32'sd29830, -32'sd389070, -32'sd138768, 32'sd380951, -32'sd1659771, -32'sd1180758, 32'sd864257, 32'sd417566, 32'sd753184, 32'sd184131, -32'sd1062409, -32'sd793802, -32'sd42554, 32'sd122479, 32'sd610062, 32'sd2077677, 32'sd2127541, 32'sd1666403, 32'sd1524994, -32'sd368305, 32'sd1023361, -32'sd15864, -32'sd563896, -32'sd988847, 32'sd2046998, 32'sd278987, -32'sd1453774, 32'sd161313, 32'sd1036605, 32'sd545431, 32'sd2596, -32'sd150376, 32'sd747121, -32'sd1061319, -32'sd796839, 32'sd152531, -32'sd361449, -32'sd1165823, -32'sd1500645, -32'sd141164, 32'sd3204893, 32'sd1857652, 32'sd4085434, 32'sd2225034, -32'sd732676, 32'sd1833260, -32'sd577929, 32'sd258584, -32'sd139307, -32'sd51085, -32'sd557240, 32'sd742935, 32'sd1947599, -32'sd577896, 32'sd1104274, 32'sd1063778, 32'sd779604, -32'sd31641, -32'sd219593, 32'sd1398195, -32'sd1247866, -32'sd993330, -32'sd3226828, -32'sd1501870, -32'sd2317513, -32'sd1194503, 32'sd1102435, 32'sd1134613, 32'sd2373592, 32'sd134727, -32'sd222732, 32'sd1271150, -32'sd801204, -32'sd982378, 32'sd1443875, -32'sd876635, 32'sd1551203, -32'sd82675, -32'sd270958, 32'sd186899, -32'sd26572, 32'sd2165826, -32'sd103196, 32'sd173565, 32'sd387108, 32'sd112955, 32'sd652429, -32'sd1370910, -32'sd628850, -32'sd2469485, -32'sd2052291, -32'sd955956, -32'sd225153, -32'sd816879, 32'sd275416, 32'sd344137, -32'sd2137070, -32'sd2070964, -32'sd2350155, -32'sd2170809, 32'sd757421, -32'sd2247136, 32'sd837234, 32'sd549197, 32'sd502770, 32'sd235109, -32'sd761695, 32'sd98573, 32'sd2098, 32'sd1218183, 32'sd558440, 32'sd247696, -32'sd1027229, -32'sd708501, -32'sd2502401, -32'sd420684, -32'sd845520, -32'sd1461789, -32'sd357440, -32'sd777734, -32'sd449047, -32'sd1008298, -32'sd1763048, -32'sd3039559, -32'sd3834047, -32'sd3761012, -32'sd3072304, 32'sd355217, 32'sd926229, 32'sd678006, -32'sd413599, 32'sd3204, 32'sd1440461, -32'sd906468, -32'sd542656, -32'sd1250433, -32'sd883040, 32'sd171634, 32'sd1118837, 32'sd98600, -32'sd294645, -32'sd3653, 32'sd164878, 32'sd1127586, 32'sd1348756, 32'sd324518, 32'sd360763, 32'sd2390203, 32'sd1123400, -32'sd1960492, 32'sd970646, 32'sd188928, -32'sd1717290, 32'sd139635, -32'sd99616, 32'sd811628, 32'sd1360893, -32'sd234564, 32'sd513433, 32'sd757909, 32'sd352420, 32'sd893291, 32'sd1920797, -32'sd2892830, -32'sd1084068, -32'sd253881, 32'sd365316, -32'sd117141, -32'sd327174, 32'sd804091, 32'sd1695081, 32'sd39182, -32'sd253363, 32'sd1024494, 32'sd545660, 32'sd3096072, 32'sd630218, 32'sd698110, 32'sd594797, -32'sd696699, 32'sd1636704, -32'sd762608, -32'sd1271119, 32'sd1195287, 32'sd1702764, -32'sd148038, 32'sd978024, -32'sd568126, 32'sd1671206, 32'sd78405, 32'sd7532, -32'sd1563529, 32'sd793477, -32'sd367728, -32'sd195774, -32'sd259629, 32'sd161580, -32'sd774064, -32'sd407659, 32'sd484596, -32'sd5703, 32'sd1213510, -32'sd2027569, -32'sd729091, 32'sd586028, 32'sd656649, 32'sd128369, -32'sd116161, 32'sd1432232, -32'sd1097975, -32'sd1451613, 32'sd417882, -32'sd421823, -32'sd154391, -32'sd1967844, 32'sd886533, 32'sd956236, -32'sd49959, -32'sd1601861, -32'sd239205, 32'sd1397297, 32'sd1308318, 32'sd1695278, 32'sd887636, 32'sd985891, 32'sd672586, -32'sd160533, 32'sd970640, 32'sd1650747, 32'sd2333115, -32'sd727651, -32'sd3562460, -32'sd5036453, -32'sd2165320, -32'sd257632, 32'sd208061, 32'sd508168, -32'sd974282, -32'sd910582, -32'sd1288843, -32'sd2069078, -32'sd2223211, -32'sd1831031, 32'sd1083584, -32'sd114665, -32'sd3099673, -32'sd1814337, -32'sd631302, -32'sd1265598, -32'sd871714, 32'sd909876, 32'sd66560, 32'sd408186, -32'sd1997467, 32'sd38567, -32'sd544517, 32'sd815574, 32'sd3127410, 32'sd1442715, 32'sd377746, -32'sd3031977, -32'sd555801, -32'sd1134010, -32'sd2435901, -32'sd1913380, -32'sd2159008, -32'sd1368609, -32'sd1297880, -32'sd856389, -32'sd1263535, -32'sd2524127, -32'sd312184, -32'sd1615342, -32'sd1127491, -32'sd1269767, -32'sd1545167, -32'sd2812045, 32'sd887932, -32'sd419856, 32'sd207643, 32'sd712248, -32'sd690875, 32'sd332982, 32'sd660995, 32'sd458137, 32'sd810293, 32'sd829436, 32'sd1873747, 32'sd1062862, 32'sd1160127, 32'sd276292, -32'sd694454, -32'sd1300374, -32'sd1140547, -32'sd1250916, -32'sd1891805, -32'sd2299743, -32'sd1876334, -32'sd1745371, -32'sd245237, 32'sd547572, -32'sd1279322, -32'sd1989480, -32'sd2328384, -32'sd946070, -32'sd630941, -32'sd346277, 32'sd0, -32'sd90005, -32'sd1394493, 32'sd260510, -32'sd1186697, -32'sd719498, -32'sd1156990, -32'sd813077, 32'sd1259286, 32'sd1386820, 32'sd737666, 32'sd681976, 32'sd3538338, 32'sd2726623, 32'sd1303338, 32'sd2019919, 32'sd766843, -32'sd320285, -32'sd743917, -32'sd2844416, -32'sd1077940, -32'sd2500937, -32'sd2366355, -32'sd1126369, -32'sd797568, 32'sd2016340, -32'sd566497, 32'sd565133, -32'sd994190, -32'sd967101, -32'sd1730157, 32'sd14949, 32'sd1030183, 32'sd625555, 32'sd183804, 32'sd774766, 32'sd338020, 32'sd1499913, 32'sd1977431, 32'sd103021, 32'sd2431058, 32'sd780883, -32'sd638814, 32'sd1723049, -32'sd289082, -32'sd1648880, -32'sd1115181, 32'sd681065, -32'sd18374, -32'sd583782, -32'sd1206992, 32'sd417352, -32'sd649008, 32'sd118107, -32'sd955939, 32'sd923218, 32'sd777001, -32'sd1497016, -32'sd475403, -32'sd750173, -32'sd1310484, 32'sd1023169, 32'sd727368, 32'sd438759, -32'sd680454, 32'sd29007, 32'sd112433, -32'sd1178593, 32'sd672376, 32'sd58013, 32'sd310341, -32'sd1289362, -32'sd2339335, 32'sd439105, -32'sd310802, 32'sd390160, -32'sd64251, -32'sd18159, -32'sd1035883, -32'sd311191, 32'sd957612, 32'sd2274878, 32'sd167880, -32'sd1512844, 32'sd0, -32'sd24681, 32'sd840151, -32'sd541509, -32'sd1607774, -32'sd517615, 32'sd1241701, -32'sd953819, -32'sd1424206, 32'sd556791, -32'sd742214, 32'sd39026, 32'sd1152637, -32'sd413398, 32'sd887415, 32'sd427370, 32'sd463083, 32'sd1730631, 32'sd412968, 32'sd1938390, -32'sd320444, -32'sd740050, -32'sd1481274, -32'sd435159, 32'sd878604, 32'sd1854100, -32'sd310400, 32'sd736901, -32'sd100710, -32'sd1213148, 32'sd1689896, -32'sd2299450, -32'sd692296, 32'sd483502, 32'sd484193, -32'sd1050979, -32'sd2330061, -32'sd388847, -32'sd739633, -32'sd1700548, -32'sd1742958, 32'sd380755, -32'sd2235727, 32'sd857666, 32'sd2337860, 32'sd2098098, 32'sd774283, 32'sd189861, 32'sd1824516, 32'sd1963867, 32'sd2472355, 32'sd1219339, -32'sd50020, 32'sd2198077, 32'sd235878, 32'sd100772, -32'sd180308, -32'sd390928, -32'sd1095911, -32'sd1185682, -32'sd883589, 32'sd484482, 32'sd634591, 32'sd680219, -32'sd706106, -32'sd2578640, -32'sd234377, -32'sd258276, -32'sd76571, -32'sd2456470, -32'sd1432859, -32'sd747916, -32'sd164869, 32'sd1431807, 32'sd713139, -32'sd878282, 32'sd1206063, 32'sd1092144, 32'sd2776839, 32'sd961317, 32'sd1369535, -32'sd55304, -32'sd229917, -32'sd128816, 32'sd0, 32'sd537098, 32'sd275999, -32'sd2076758, -32'sd1015065, 32'sd121946, -32'sd211697, -32'sd58098, 32'sd856608, -32'sd1092812, -32'sd55763, 32'sd1367389, -32'sd1063151, -32'sd1514868, 32'sd1286751, 32'sd916677, 32'sd816747, 32'sd1993787, 32'sd1776806, -32'sd100000, -32'sd474042, 32'sd1097338, 32'sd1145714, 32'sd840681, -32'sd1793979, 32'sd1332998, -32'sd1213461, 32'sd0, 32'sd0, 32'sd0, 32'sd243267, 32'sd132205, -32'sd1333936, -32'sd1723965, -32'sd167732, 32'sd44962, 32'sd91645, -32'sd225725, -32'sd182716, -32'sd539851, 32'sd1773635, 32'sd3151527, 32'sd1858162, 32'sd999703, 32'sd2252137, 32'sd1498533, 32'sd1288150, 32'sd1175626, -32'sd663300, 32'sd448844, 32'sd964725, 32'sd1069356, -32'sd313496, 32'sd720257, 32'sd1074302, 32'sd0, 32'sd0, 32'sd0, -32'sd443925, -32'sd418563, -32'sd553864, -32'sd1233593, -32'sd319616, 32'sd891603, 32'sd1860316, -32'sd502240, -32'sd37416, 32'sd308991, 32'sd757706, 32'sd2827712, -32'sd702561, 32'sd2507923, 32'sd1515240, 32'sd3006880, 32'sd73384, -32'sd1215469, 32'sd389989, -32'sd958098, 32'sd1553999, 32'sd619966, -32'sd441942, -32'sd985048, -32'sd493199, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd593257, 32'sd687029, 32'sd744568, -32'sd724999, 32'sd1112185, 32'sd878681, 32'sd761889, -32'sd39128, 32'sd566029, 32'sd2819805, 32'sd970204, 32'sd1784984, 32'sd2302770, -32'sd235743, 32'sd1219084, 32'sd1054632, 32'sd393111, 32'sd980165, 32'sd84743, -32'sd287177, 32'sd1968743, 32'sd828108, 32'sd1290394, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd39573, 32'sd1416410, -32'sd441553, 32'sd257439, 32'sd120026, 32'sd248709, -32'sd1142904, 32'sd326566, 32'sd1344241, -32'sd205284, 32'sd644437, 32'sd1092608, 32'sd14245, -32'sd687382, 32'sd578422, 32'sd221445, -32'sd637780, 32'sd1582094, 32'sd3091042, -32'sd157450, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd164670, -32'sd901745, 32'sd1512551, 32'sd536967, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd511766, -32'sd1115086, -32'sd292327, 32'sd127109, 32'sd396610, -32'sd886265, -32'sd181931, -32'sd273721, -32'sd318384, -32'sd1409300, 32'sd683785, 32'sd204632, 32'sd1269469, -32'sd541337, 32'sd39293, -32'sd1221463, 32'sd1119229, 32'sd285373, -32'sd577528, 32'sd26795, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd416938, -32'sd400826, 32'sd357471, -32'sd487399, 32'sd193567, -32'sd742901, -32'sd1159405, -32'sd841465, -32'sd882974, -32'sd1518195, -32'sd2037102, -32'sd192291, 32'sd771205, 32'sd182275, 32'sd487308, 32'sd561135, -32'sd228824, -32'sd1699578, -32'sd1778896, -32'sd1121983, 32'sd839435, 32'sd395364, -32'sd1002769, -32'sd430616, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd105346, -32'sd1124543, -32'sd79359, -32'sd1446869, -32'sd1549088, 32'sd265627, -32'sd1501360, -32'sd2368352, -32'sd2278388, -32'sd1213612, -32'sd2090229, -32'sd2399823, -32'sd1623902, -32'sd814142, 32'sd814772, 32'sd3821599, 32'sd3026770, 32'sd734864, 32'sd133206, -32'sd868243, 32'sd654944, -32'sd550126, -32'sd472826, 32'sd665159, -32'sd687315, 32'sd0, 32'sd0, 32'sd288066, 32'sd517719, 32'sd1117117, -32'sd33508, 32'sd234130, -32'sd1322274, 32'sd43071, -32'sd2163208, -32'sd291314, 32'sd1085827, 32'sd356167, -32'sd123333, 32'sd495900, -32'sd1328843, -32'sd1041863, -32'sd280315, 32'sd1304756, 32'sd3329860, 32'sd1216775, -32'sd275459, -32'sd139152, -32'sd1251082, -32'sd475583, -32'sd348774, -32'sd868824, -32'sd1245482, 32'sd506299, 32'sd0, 32'sd531901, -32'sd132526, -32'sd941400, -32'sd71504, -32'sd132159, -32'sd682536, -32'sd2137096, -32'sd541035, -32'sd1889057, -32'sd150653, -32'sd205283, 32'sd385212, -32'sd1465149, -32'sd864439, -32'sd1536909, -32'sd492195, -32'sd1122860, 32'sd2543974, 32'sd3766661, 32'sd3621228, 32'sd615179, -32'sd804309, -32'sd1464750, 32'sd13617, -32'sd1320858, -32'sd1446443, -32'sd453991, 32'sd0, 32'sd953097, -32'sd1653059, 32'sd906239, -32'sd19968, 32'sd630937, -32'sd750070, -32'sd1606089, -32'sd1880891, -32'sd148072, -32'sd396741, 32'sd1550421, 32'sd1907919, -32'sd893435, -32'sd2634064, -32'sd244859, -32'sd615930, -32'sd1769567, 32'sd114955, 32'sd298329, 32'sd3943221, 32'sd360335, -32'sd1401934, 32'sd514007, 32'sd247968, -32'sd2675972, 32'sd362239, -32'sd591065, 32'sd125560, -32'sd771054, 32'sd1442890, 32'sd88184, 32'sd1310473, -32'sd597037, 32'sd1287937, 32'sd397194, -32'sd1500436, 32'sd996064, 32'sd582359, 32'sd814030, 32'sd1369450, -32'sd2138709, -32'sd1079090, -32'sd903051, 32'sd847094, -32'sd840780, 32'sd1054065, 32'sd1185522, 32'sd1051604, 32'sd1157213, 32'sd585693, -32'sd321815, 32'sd13330, -32'sd3428201, 32'sd223818, -32'sd335680, -32'sd20857, 32'sd377534, 32'sd1467332, 32'sd1700734, 32'sd1848611, 32'sd703361, 32'sd1406209, 32'sd41869, 32'sd1727508, 32'sd961942, -32'sd437029, -32'sd1244132, -32'sd1921393, -32'sd2404766, -32'sd2059882, -32'sd2553914, -32'sd946626, -32'sd740520, 32'sd1151044, 32'sd3742985, 32'sd1511031, 32'sd1557105, -32'sd549305, -32'sd1819500, -32'sd208204, -32'sd488330, -32'sd453694, -32'sd1573285, -32'sd468366, 32'sd707391, -32'sd58833, 32'sd1121686, 32'sd1409083, 32'sd1802840, 32'sd2805033, 32'sd1787675, 32'sd349303, -32'sd1902138, -32'sd4311482, -32'sd2226296, -32'sd2913155, -32'sd973892, -32'sd3109684, -32'sd547696, -32'sd1247511, 32'sd2028539, 32'sd4752913, 32'sd2704332, 32'sd2424174, -32'sd186622, -32'sd2034241, -32'sd311136, -32'sd3817932, -32'sd2899518, -32'sd738014, 32'sd690928, 32'sd29330, 32'sd428288, 32'sd368453, 32'sd566881, 32'sd189214, 32'sd737582, 32'sd1427066, -32'sd466643, 32'sd692642, -32'sd2110946, -32'sd3506250, -32'sd3024196, -32'sd6305, -32'sd2584121, -32'sd2319950, -32'sd2904568, -32'sd1097228, 32'sd2422204, 32'sd5167204, 32'sd2108897, 32'sd510145, 32'sd51353, -32'sd874731, -32'sd1773217, -32'sd2266642, 32'sd5130, 32'sd141967, 32'sd551034, 32'sd210594, -32'sd572947, -32'sd135840, -32'sd449801, 32'sd225478, 32'sd1445382, 32'sd841988, 32'sd857540, -32'sd2381085, -32'sd3282196, 32'sd159083, 32'sd579919, 32'sd431993, -32'sd2722639, -32'sd1792871, -32'sd51554, 32'sd1084088, 32'sd2039812, 32'sd2467754, 32'sd612878, -32'sd2123731, -32'sd2714432, -32'sd4393382, -32'sd2589139, -32'sd499200, 32'sd1757593, 32'sd907855, 32'sd781883, 32'sd130473, -32'sd364195, 32'sd357811, -32'sd553319, 32'sd63764, 32'sd776951, 32'sd912563, 32'sd1462588, -32'sd1846435, -32'sd2265316, 32'sd1128997, 32'sd58152, 32'sd1979218, -32'sd606275, 32'sd616682, -32'sd714014, 32'sd3565663, 32'sd1668979, 32'sd2448327, -32'sd1725320, -32'sd3043221, -32'sd3236351, -32'sd3603883, -32'sd999823, -32'sd1649635, -32'sd397444, -32'sd606765, 32'sd140514, 32'sd28525, -32'sd80510, -32'sd1442569, 32'sd728169, 32'sd1447409, -32'sd565108, 32'sd60578, 32'sd1671833, 32'sd1353444, 32'sd134113, 32'sd3107763, 32'sd3517167, 32'sd854260, 32'sd1531509, 32'sd333029, -32'sd250230, 32'sd2002441, 32'sd2559186, 32'sd1379685, -32'sd2198079, -32'sd2359374, -32'sd611821, -32'sd1598921, -32'sd1145650, -32'sd695369, -32'sd523567, 32'sd622390, -32'sd805672, -32'sd424860, 32'sd637995, -32'sd1716968, 32'sd1271025, -32'sd947382, 32'sd1096961, 32'sd1341076, 32'sd1848712, 32'sd2755748, 32'sd3245049, 32'sd3774890, 32'sd2243138, 32'sd993144, 32'sd325666, -32'sd457437, 32'sd1325650, 32'sd2168238, 32'sd2747910, -32'sd1230214, -32'sd991824, 32'sd1266529, 32'sd286503, -32'sd647051, 32'sd596003, -32'sd742058, -32'sd790648, -32'sd786105, -32'sd451034, -32'sd33628, 32'sd904261, 32'sd301957, 32'sd1251205, 32'sd683193, 32'sd321145, 32'sd114325, 32'sd685072, 32'sd2111654, 32'sd2765409, 32'sd2948856, 32'sd1328547, 32'sd2222237, 32'sd3829214, 32'sd880276, 32'sd1607726, -32'sd725717, 32'sd873533, -32'sd702575, 32'sd2086056, 32'sd1621261, -32'sd478145, 32'sd1548209, 32'sd1133176, -32'sd636757, 32'sd252515, -32'sd1695834, 32'sd177367, 32'sd366221, -32'sd827960, -32'sd546515, -32'sd998005, 32'sd1833631, -32'sd120992, -32'sd396503, 32'sd339331, 32'sd150647, 32'sd1604603, -32'sd1128275, 32'sd1544571, 32'sd2155355, 32'sd2084059, 32'sd1166272, 32'sd1491602, -32'sd473184, -32'sd29304, 32'sd2602076, 32'sd1407859, 32'sd1099871, 32'sd2504173, 32'sd610737, -32'sd251688, 32'sd1831829, 32'sd1226824, -32'sd2760768, 32'sd560051, 32'sd0, 32'sd697425, 32'sd218114, -32'sd97481, 32'sd107974, 32'sd183632, 32'sd969071, 32'sd624417, -32'sd614795, -32'sd2878889, -32'sd1308051, -32'sd1182948, 32'sd23061, 32'sd626130, 32'sd841837, 32'sd1865471, -32'sd1254894, -32'sd240327, 32'sd1533431, -32'sd558822, -32'sd141089, 32'sd1841954, 32'sd2148193, 32'sd278547, 32'sd1021922, -32'sd229439, -32'sd706623, -32'sd659944, 32'sd655072, -32'sd113881, 32'sd690210, 32'sd1985278, 32'sd512768, 32'sd1085761, -32'sd673976, -32'sd1023784, -32'sd1546916, -32'sd990652, -32'sd2561421, -32'sd650110, -32'sd804770, -32'sd1706580, -32'sd1105748, -32'sd950016, 32'sd800156, 32'sd1787087, 32'sd185288, -32'sd776742, -32'sd382488, 32'sd341512, 32'sd1555141, -32'sd2604543, -32'sd1670417, -32'sd1482129, -32'sd322317, -32'sd973413, -32'sd159102, -32'sd169012, 32'sd1292756, 32'sd2392269, 32'sd306655, 32'sd2551431, 32'sd1188802, -32'sd1690206, -32'sd2790437, -32'sd3133086, -32'sd2137727, -32'sd319945, -32'sd3105337, -32'sd1873276, 32'sd608097, 32'sd31890, 32'sd194502, 32'sd1379555, -32'sd228626, 32'sd267820, -32'sd541040, 32'sd678282, -32'sd571697, -32'sd323691, -32'sd1581743, -32'sd266372, 32'sd216688, -32'sd131475, 32'sd0, 32'sd1406814, 32'sd281379, 32'sd773264, -32'sd192635, 32'sd206886, -32'sd256745, -32'sd1435642, -32'sd1810412, -32'sd2034448, -32'sd3246799, -32'sd2698367, -32'sd2722939, -32'sd1814643, -32'sd2621287, -32'sd2154676, -32'sd2065145, 32'sd981038, -32'sd134558, 32'sd559613, 32'sd51617, -32'sd500418, 32'sd1779947, 32'sd134502, 32'sd1296025, -32'sd1089729, 32'sd230517, 32'sd466729, 32'sd667908, -32'sd353878, 32'sd675043, -32'sd409405, -32'sd815925, 32'sd2004019, 32'sd1339810, 32'sd1040040, 32'sd603749, -32'sd750590, -32'sd2475817, 32'sd332416, -32'sd539580, -32'sd1364327, -32'sd368199, 32'sd59451, 32'sd179176, 32'sd762779, 32'sd985016, 32'sd1280165, 32'sd224263, 32'sd1383627, 32'sd1275126, -32'sd133192, 32'sd2252783, 32'sd2221657, -32'sd207451, -32'sd151399, 32'sd141463, 32'sd1025928, 32'sd283293, 32'sd107609, -32'sd798340, -32'sd1614700, -32'sd641386, -32'sd276997, -32'sd514251, -32'sd1764570, -32'sd847898, 32'sd1388937, -32'sd403050, 32'sd747409, -32'sd1118066, -32'sd898909, 32'sd1574086, 32'sd2284232, 32'sd2209242, 32'sd1409829, 32'sd1763537, 32'sd500880, -32'sd542480, -32'sd1233491, 32'sd1016175, -32'sd310126, 32'sd1592455, 32'sd10636, 32'sd0, 32'sd823942, 32'sd341143, 32'sd1884192, 32'sd1158894, -32'sd391575, -32'sd503418, 32'sd1283890, -32'sd433290, -32'sd489725, 32'sd717081, 32'sd1608278, 32'sd68747, 32'sd2013317, 32'sd1365939, 32'sd185989, 32'sd677506, 32'sd729524, -32'sd701593, -32'sd264953, 32'sd869626, 32'sd190184, 32'sd469173, 32'sd357041, 32'sd369184, -32'sd844892, 32'sd1332381, 32'sd0, 32'sd0, 32'sd0, 32'sd952725, 32'sd1003337, 32'sd707179, -32'sd1084587, 32'sd850168, -32'sd391008, -32'sd1383194, -32'sd280122, 32'sd1143554, 32'sd762649, -32'sd497629, -32'sd682650, 32'sd178611, -32'sd400867, 32'sd209491, -32'sd808352, 32'sd740610, -32'sd18844, 32'sd662628, 32'sd519437, -32'sd674694, -32'sd1316170, 32'sd506125, -32'sd884964, -32'sd172997, 32'sd0, 32'sd0, 32'sd0, 32'sd454329, -32'sd1288955, -32'sd360268, -32'sd253557, 32'sd1677189, 32'sd990280, -32'sd968284, -32'sd1520466, -32'sd1014597, 32'sd45367, -32'sd2170609, -32'sd831758, 32'sd36224, -32'sd1506920, -32'sd981572, -32'sd47029, 32'sd2654751, 32'sd2149141, -32'sd675032, -32'sd1476957, -32'sd247586, 32'sd279481, -32'sd970553, 32'sd278306, -32'sd475100, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd639856, 32'sd161343, -32'sd1299531, -32'sd553009, 32'sd2144474, -32'sd1255283, -32'sd584935, -32'sd631494, 32'sd553600, 32'sd2155299, 32'sd975497, 32'sd569796, 32'sd588043, -32'sd863699, -32'sd1524576, -32'sd174598, -32'sd1880295, -32'sd551970, 32'sd23459, -32'sd1007124, -32'sd139496, -32'sd855295, 32'sd433719, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd326516, 32'sd187814, 32'sd1049623, 32'sd56581, -32'sd539734, -32'sd1066141, 32'sd115820, -32'sd376761, -32'sd184455, 32'sd41115, 32'sd135859, 32'sd727590, 32'sd77035, 32'sd745410, 32'sd1378005, -32'sd303922, -32'sd292343, -32'sd218081, -32'sd1030745, 32'sd169223, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1166351, 32'sd816495, -32'sd357634, 32'sd281261, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd406264, -32'sd600926, -32'sd234268, 32'sd582840, -32'sd400862, 32'sd717402, 32'sd150812, -32'sd581919, 32'sd107157, -32'sd275491, -32'sd493979, 32'sd767792, 32'sd191120, 32'sd2216, -32'sd1100503, 32'sd359088, -32'sd706202, -32'sd680241, -32'sd1360846, 32'sd423268, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd156954, -32'sd150161, 32'sd1377167, 32'sd211641, -32'sd947655, -32'sd185686, -32'sd272075, -32'sd1191063, 32'sd155245, 32'sd83531, -32'sd2759780, -32'sd2983081, -32'sd518513, -32'sd1060892, -32'sd851264, -32'sd459353, 32'sd1325764, 32'sd128217, 32'sd1582135, 32'sd1258376, 32'sd583117, 32'sd1009083, 32'sd159117, 32'sd217241, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd761219, -32'sd414065, 32'sd615075, 32'sd993934, 32'sd826405, 32'sd381055, 32'sd1151737, -32'sd1847708, -32'sd1075000, 32'sd545768, -32'sd1783965, -32'sd360460, -32'sd1345162, 32'sd352289, 32'sd1544502, 32'sd593848, -32'sd1252895, -32'sd2246376, 32'sd180988, -32'sd1936852, -32'sd1759895, -32'sd121748, 32'sd591734, -32'sd664010, -32'sd282144, 32'sd0, 32'sd0, 32'sd266440, 32'sd505499, -32'sd1972093, -32'sd852263, 32'sd1024273, -32'sd1363020, -32'sd555362, 32'sd893652, 32'sd907623, -32'sd1651411, 32'sd1889872, 32'sd851847, 32'sd443895, -32'sd686498, -32'sd1782725, 32'sd856003, 32'sd34794, -32'sd1400884, 32'sd146713, -32'sd184298, 32'sd480043, 32'sd842857, -32'sd63106, -32'sd627912, -32'sd309079, 32'sd601912, -32'sd441584, 32'sd0, -32'sd349112, -32'sd722765, -32'sd256855, -32'sd118537, 32'sd1218377, -32'sd604669, -32'sd614076, -32'sd97451, -32'sd1516994, -32'sd151639, 32'sd755449, 32'sd2258980, -32'sd860637, -32'sd96283, 32'sd1952551, 32'sd1767190, -32'sd478071, -32'sd1832099, -32'sd1558914, 32'sd499451, 32'sd294588, -32'sd557491, 32'sd172822, 32'sd558814, 32'sd682587, 32'sd488093, -32'sd692851, 32'sd0, 32'sd664263, 32'sd781248, -32'sd181130, -32'sd792058, 32'sd1542597, 32'sd63552, 32'sd454129, -32'sd532917, -32'sd1107527, -32'sd351033, 32'sd2065008, 32'sd168993, -32'sd84481, 32'sd1455096, -32'sd203294, 32'sd393783, -32'sd604361, -32'sd2672808, -32'sd2871159, -32'sd670632, 32'sd1402683, 32'sd617264, 32'sd2011883, -32'sd1212727, -32'sd2661071, 32'sd1721721, -32'sd1591661, 32'sd244494, -32'sd823734, -32'sd929624, -32'sd2349266, -32'sd741606, 32'sd1613482, -32'sd1322503, 32'sd1906492, 32'sd1047471, -32'sd935176, 32'sd1652413, 32'sd2801736, 32'sd1502693, 32'sd1576623, -32'sd714458, -32'sd3103551, -32'sd1856958, -32'sd1344708, -32'sd1891291, -32'sd1200678, -32'sd1368016, 32'sd365516, 32'sd521607, -32'sd763817, 32'sd423265, 32'sd384783, 32'sd90671, -32'sd1775018, 32'sd241518, -32'sd1348721, -32'sd557889, -32'sd623768, -32'sd1268617, -32'sd355775, -32'sd2008420, 32'sd858585, -32'sd461148, 32'sd244409, 32'sd786375, 32'sd1226296, 32'sd3332924, 32'sd316131, 32'sd578489, 32'sd237075, -32'sd2160168, -32'sd641702, -32'sd492255, -32'sd840275, 32'sd432007, 32'sd1433997, 32'sd1576516, 32'sd557955, -32'sd221880, 32'sd1505250, -32'sd856645, 32'sd34082, 32'sd88477, 32'sd1585239, 32'sd1757515, -32'sd85429, 32'sd213128, -32'sd1050434, -32'sd22128, -32'sd989287, 32'sd527418, 32'sd994011, 32'sd1585615, 32'sd381012, 32'sd265980, 32'sd2148447, -32'sd244851, -32'sd1926702, 32'sd387069, -32'sd562766, 32'sd1191571, 32'sd361540, 32'sd248322, 32'sd2645698, 32'sd1740603, 32'sd1850254, -32'sd849940, 32'sd323751, 32'sd1238360, -32'sd808833, 32'sd1626179, 32'sd1096932, 32'sd1982092, 32'sd1140038, -32'sd123959, 32'sd734946, -32'sd1119632, -32'sd1521635, -32'sd2055851, -32'sd2936598, -32'sd74112, 32'sd564603, 32'sd2403084, 32'sd464725, 32'sd935134, -32'sd847944, -32'sd1529533, -32'sd473532, 32'sd254832, 32'sd1480558, 32'sd2032230, 32'sd2497249, 32'sd1583934, 32'sd2468328, 32'sd786658, 32'sd2084707, 32'sd1280128, 32'sd1042108, -32'sd187228, 32'sd1047845, 32'sd964501, 32'sd1558818, 32'sd250017, 32'sd710219, 32'sd391364, -32'sd1337311, 32'sd190974, -32'sd1841185, -32'sd580374, 32'sd1031237, 32'sd1399300, -32'sd1501298, 32'sd450830, -32'sd2952612, -32'sd2009957, -32'sd1102981, -32'sd557394, 32'sd1170149, 32'sd1044766, 32'sd809287, -32'sd581803, -32'sd601553, -32'sd234503, -32'sd311002, -32'sd930914, -32'sd1956321, 32'sd208855, 32'sd1550604, 32'sd763614, 32'sd740216, 32'sd1663682, 32'sd1424125, -32'sd492098, 32'sd14450, 32'sd134545, -32'sd28939, 32'sd3229209, 32'sd1329910, 32'sd2770554, 32'sd1162906, -32'sd516220, -32'sd1862091, -32'sd284846, 32'sd199166, 32'sd1252983, -32'sd194478, 32'sd1165019, 32'sd1822025, 32'sd1540317, -32'sd451144, 32'sd753170, 32'sd979074, 32'sd966786, -32'sd1246057, 32'sd1028203, 32'sd1026295, 32'sd285192, 32'sd598901, 32'sd1057437, -32'sd998390, -32'sd513344, -32'sd138861, 32'sd157592, 32'sd3161026, 32'sd3957875, 32'sd3772349, 32'sd2907572, 32'sd265591, 32'sd317216, 32'sd943063, -32'sd337737, 32'sd1311123, 32'sd1900969, 32'sd338207, 32'sd1603966, 32'sd1349775, -32'sd199909, 32'sd64173, -32'sd599862, -32'sd435453, -32'sd978827, 32'sd294204, 32'sd11386, -32'sd85408, 32'sd747970, 32'sd383241, -32'sd458274, 32'sd929933, -32'sd1012507, -32'sd459206, 32'sd2082381, 32'sd3651900, 32'sd2453080, 32'sd3272619, 32'sd3541541, 32'sd3513018, 32'sd3245887, 32'sd3048956, 32'sd349738, 32'sd1493104, 32'sd783056, -32'sd18444, 32'sd14686, 32'sd2627194, 32'sd84615, -32'sd837903, 32'sd536573, -32'sd138461, -32'sd809840, 32'sd636539, -32'sd403018, -32'sd182091, 32'sd1353424, -32'sd414083, 32'sd513358, 32'sd273580, -32'sd1472171, -32'sd1056099, 32'sd222518, -32'sd193772, 32'sd2692544, 32'sd3374538, 32'sd2782468, 32'sd2900534, 32'sd2234450, 32'sd1257546, 32'sd1419077, 32'sd2234840, -32'sd608762, -32'sd309861, 32'sd331666, -32'sd102874, -32'sd10553, -32'sd1478073, -32'sd1272076, 32'sd69266, 32'sd793104, 32'sd201840, 32'sd363702, -32'sd397751, -32'sd1082514, 32'sd964191, 32'sd1319780, 32'sd219655, -32'sd771758, -32'sd1973967, -32'sd774006, -32'sd592715, 32'sd68866, 32'sd646076, 32'sd2790920, 32'sd3586402, 32'sd852957, 32'sd154712, -32'sd266556, -32'sd1421759, -32'sd1642105, -32'sd3660175, -32'sd1778019, 32'sd846167, 32'sd620057, -32'sd1036611, 32'sd1562474, -32'sd3068256, -32'sd260372, -32'sd266669, 32'sd0, 32'sd1356814, 32'sd215998, -32'sd1651311, -32'sd39781, -32'sd362671, -32'sd2864755, -32'sd871111, -32'sd3782543, -32'sd4851403, -32'sd5940954, -32'sd2962144, -32'sd1536732, 32'sd357430, 32'sd1082934, -32'sd878301, -32'sd640136, -32'sd797961, -32'sd2133976, -32'sd2734356, 32'sd421236, 32'sd225082, 32'sd1579092, 32'sd485862, 32'sd2113413, -32'sd840331, 32'sd1534716, -32'sd1068505, -32'sd305009, 32'sd1277450, -32'sd1473019, -32'sd171680, -32'sd909798, -32'sd2228852, -32'sd1860618, -32'sd2473234, -32'sd2521060, -32'sd5673791, -32'sd5319254, -32'sd2570163, -32'sd1699179, -32'sd111984, -32'sd532596, -32'sd1907219, -32'sd316609, -32'sd2664779, -32'sd3240371, -32'sd3698765, -32'sd2239870, 32'sd617546, 32'sd787884, 32'sd222831, -32'sd832807, 32'sd652589, 32'sd896868, -32'sd606268, 32'sd163292, 32'sd138795, -32'sd42308, 32'sd507366, 32'sd563424, -32'sd2869077, -32'sd3144578, -32'sd2667593, -32'sd4277602, -32'sd1661873, -32'sd2354154, -32'sd2353582, -32'sd3115599, -32'sd2143365, 32'sd101196, 32'sd85197, 32'sd629794, -32'sd127974, -32'sd1134354, -32'sd1292881, -32'sd2048156, 32'sd1726540, 32'sd1228292, -32'sd1235198, 32'sd226877, 32'sd1758559, 32'sd146828, -32'sd545213, 32'sd0, 32'sd1368126, 32'sd577704, -32'sd714840, 32'sd1264270, -32'sd2213554, -32'sd1797065, -32'sd1508869, -32'sd3048401, 32'sd1262893, 32'sd608804, 32'sd85049, -32'sd1652163, 32'sd523984, 32'sd1739917, -32'sd691046, -32'sd223191, 32'sd607996, -32'sd316614, -32'sd1296560, -32'sd1491017, -32'sd574084, 32'sd1964449, 32'sd1309894, -32'sd1092129, -32'sd978174, -32'sd342163, 32'sd412774, 32'sd953652, 32'sd735721, -32'sd670625, 32'sd112604, 32'sd2008806, -32'sd1360104, 32'sd1299231, 32'sd618590, 32'sd2105462, -32'sd41731, 32'sd725802, 32'sd1012516, 32'sd265322, -32'sd1475710, -32'sd1477362, -32'sd116181, -32'sd186517, -32'sd2386096, -32'sd139331, -32'sd2174519, -32'sd942447, 32'sd126856, -32'sd428159, 32'sd708782, 32'sd200197, -32'sd1708786, 32'sd773066, -32'sd191047, 32'sd595546, 32'sd1537155, -32'sd100021, -32'sd6082, 32'sd2914747, -32'sd445424, 32'sd148756, 32'sd2107971, 32'sd1869674, 32'sd428671, -32'sd81398, 32'sd1393428, 32'sd1708643, 32'sd1166151, 32'sd495322, 32'sd45953, -32'sd1247728, -32'sd142877, 32'sd127958, -32'sd394610, -32'sd416178, 32'sd213801, 32'sd857579, 32'sd953671, 32'sd750782, -32'sd2376234, -32'sd1970628, -32'sd592424, 32'sd0, 32'sd738035, -32'sd790699, -32'sd1158267, -32'sd730062, 32'sd385650, 32'sd1220083, -32'sd60053, 32'sd2642128, 32'sd740538, 32'sd1745973, 32'sd613762, 32'sd138404, 32'sd1972004, 32'sd1642244, -32'sd2125338, -32'sd576011, 32'sd908042, -32'sd1095595, -32'sd138709, -32'sd655149, -32'sd93221, 32'sd557854, 32'sd387807, -32'sd219114, 32'sd291125, -32'sd896282, 32'sd0, 32'sd0, 32'sd0, -32'sd381894, -32'sd158058, -32'sd167597, -32'sd799859, -32'sd1506210, 32'sd219903, -32'sd385624, -32'sd727454, 32'sd211159, 32'sd515256, 32'sd61947, 32'sd485310, 32'sd2746177, -32'sd1685105, -32'sd1848339, -32'sd958238, -32'sd500907, 32'sd1511548, -32'sd303519, 32'sd1148256, 32'sd84795, -32'sd1072527, 32'sd970003, -32'sd383934, 32'sd802191, 32'sd0, 32'sd0, 32'sd0, -32'sd538611, 32'sd26905, 32'sd1075653, 32'sd649345, -32'sd145586, -32'sd616122, 32'sd1159704, -32'sd244867, -32'sd968182, 32'sd134336, -32'sd1355225, -32'sd204688, 32'sd1047004, -32'sd1101318, -32'sd2537454, -32'sd1576940, 32'sd1596570, 32'sd787641, 32'sd614214, -32'sd1086832, -32'sd191912, 32'sd534943, 32'sd534608, 32'sd418885, -32'sd368093, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd26936, 32'sd1719704, -32'sd1224903, 32'sd886671, -32'sd101851, 32'sd233201, -32'sd287689, -32'sd563146, -32'sd1672063, -32'sd1072704, -32'sd646665, -32'sd2091978, -32'sd1121043, -32'sd110604, 32'sd371831, -32'sd1142816, -32'sd424356, 32'sd271027, -32'sd798431, -32'sd1569396, 32'sd927212, -32'sd562200, 32'sd380751, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd509621, -32'sd126145, -32'sd701210, -32'sd670196, 32'sd979497, 32'sd177072, 32'sd22637, -32'sd1133922, -32'sd1445044, 32'sd114851, -32'sd765976, 32'sd349290, -32'sd905795, -32'sd1274921, -32'sd495167, -32'sd437270, 32'sd752449, 32'sd1413934, -32'sd71422, 32'sd13301, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1524586, -32'sd591317, -32'sd303940, 32'sd230701, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd45605, -32'sd151178, -32'sd257009, -32'sd915482, -32'sd137607, -32'sd1856320, -32'sd697993, 32'sd323797, -32'sd187596, -32'sd309527, -32'sd750970, 32'sd21338, -32'sd926647, 32'sd453, 32'sd336306, 32'sd1153128, -32'sd293015, -32'sd682631, -32'sd947872, 32'sd773829, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd139658, -32'sd302890, -32'sd310305, -32'sd942337, -32'sd1004829, 32'sd456192, 32'sd687634, 32'sd645392, -32'sd1392546, -32'sd734987, 32'sd632607, 32'sd379036, -32'sd906152, -32'sd1479929, -32'sd1386713, -32'sd956905, 32'sd1183024, -32'sd960836, -32'sd254121, 32'sd2356581, 32'sd2698535, 32'sd1737107, 32'sd1215582, 32'sd214020, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1053085, -32'sd784566, -32'sd1315312, 32'sd102446, -32'sd2055383, -32'sd1891115, -32'sd1822570, -32'sd316983, 32'sd1214735, 32'sd420551, 32'sd1987411, 32'sd335653, -32'sd1224975, -32'sd1513364, -32'sd475431, 32'sd110565, 32'sd1053503, 32'sd190813, -32'sd806929, 32'sd1496941, -32'sd543874, 32'sd461551, -32'sd711241, -32'sd956371, 32'sd194207, 32'sd0, 32'sd0, 32'sd727750, 32'sd66618, -32'sd1041525, 32'sd317466, -32'sd386277, -32'sd183010, 32'sd1077501, 32'sd663075, -32'sd747376, 32'sd2605867, 32'sd1300584, 32'sd2139439, 32'sd2712444, 32'sd1849535, -32'sd483912, -32'sd2030957, -32'sd733631, -32'sd717161, 32'sd15448, 32'sd1470359, 32'sd1498509, -32'sd708883, 32'sd206301, 32'sd220274, 32'sd1067035, 32'sd990923, 32'sd1319379, 32'sd0, -32'sd835393, 32'sd1255336, -32'sd813251, 32'sd706096, 32'sd205541, 32'sd413796, 32'sd1612320, 32'sd1339131, -32'sd1020674, 32'sd1875241, 32'sd2568936, 32'sd1507746, 32'sd426790, 32'sd190727, 32'sd286335, -32'sd55586, 32'sd519291, 32'sd951303, -32'sd175216, 32'sd252004, 32'sd1509001, -32'sd1022021, 32'sd1733022, -32'sd1774607, 32'sd774524, 32'sd336240, 32'sd347321, 32'sd0, -32'sd367642, 32'sd380692, -32'sd1427110, -32'sd1190345, -32'sd3089593, -32'sd1356740, -32'sd314551, 32'sd535152, 32'sd683907, 32'sd2047124, 32'sd641778, -32'sd262057, -32'sd1890764, 32'sd91056, -32'sd444059, 32'sd1849433, 32'sd2398442, 32'sd647051, -32'sd1938980, -32'sd2885414, -32'sd1237332, -32'sd114659, 32'sd162234, -32'sd464754, -32'sd1027208, 32'sd1195633, -32'sd338058, -32'sd349230, -32'sd303799, -32'sd642072, -32'sd18090, 32'sd196723, -32'sd2376149, -32'sd1012825, -32'sd1487042, -32'sd479409, 32'sd877375, 32'sd3481336, -32'sd1196375, -32'sd2533198, -32'sd2795603, -32'sd226651, 32'sd941922, -32'sd141891, 32'sd1349111, -32'sd1859197, -32'sd3781004, -32'sd1456453, -32'sd1629674, 32'sd99865, -32'sd1389268, 32'sd1412922, 32'sd1639905, -32'sd259788, 32'sd872092, 32'sd95420, -32'sd1376769, 32'sd104480, 32'sd309004, 32'sd2012637, -32'sd2216892, 32'sd154727, -32'sd318685, 32'sd606519, 32'sd803804, 32'sd2382253, 32'sd1696433, -32'sd1120405, -32'sd1343623, -32'sd923062, 32'sd935592, -32'sd1319003, 32'sd928397, -32'sd1827838, -32'sd3362439, -32'sd2496948, -32'sd3557483, -32'sd1772099, 32'sd615851, 32'sd1101528, 32'sd1236885, 32'sd309410, -32'sd397126, 32'sd218958, 32'sd797290, 32'sd265406, 32'sd1262165, -32'sd348066, -32'sd914847, -32'sd538068, -32'sd2247189, -32'sd625770, 32'sd2090704, 32'sd1378501, -32'sd1299146, -32'sd948794, -32'sd2237223, -32'sd86956, -32'sd496111, -32'sd2766740, -32'sd2010987, -32'sd2200181, -32'sd1524999, -32'sd1598476, -32'sd1855052, 32'sd1553207, 32'sd1972532, 32'sd773265, 32'sd2413969, 32'sd420360, -32'sd764991, 32'sd86578, 32'sd477777, 32'sd1161174, 32'sd746419, 32'sd2891267, -32'sd1114328, 32'sd709539, 32'sd1424796, 32'sd408541, 32'sd969753, 32'sd1106653, -32'sd751614, -32'sd1869314, -32'sd1215773, 32'sd1302381, 32'sd1095867, -32'sd939836, -32'sd833027, 32'sd182788, -32'sd478047, -32'sd1352439, 32'sd513759, -32'sd171798, 32'sd387492, 32'sd1021151, -32'sd436344, -32'sd962439, 32'sd360695, -32'sd458020, -32'sd311021, 32'sd2031605, 32'sd655877, 32'sd595835, -32'sd1016217, 32'sd448591, 32'sd743381, 32'sd2071449, 32'sd2054849, -32'sd1163964, 32'sd59102, -32'sd884658, -32'sd1472475, 32'sd1958912, 32'sd971414, 32'sd768659, -32'sd893824, -32'sd1257118, 32'sd1390936, 32'sd545312, 32'sd1283855, -32'sd766957, 32'sd898104, 32'sd1697333, 32'sd1408247, 32'sd1162811, 32'sd776679, -32'sd925616, 32'sd1326262, 32'sd1531060, -32'sd781458, 32'sd133640, -32'sd1206118, 32'sd678818, 32'sd1287207, 32'sd221305, -32'sd202244, 32'sd2127670, 32'sd58707, -32'sd1160533, 32'sd67457, -32'sd393531, 32'sd141917, 32'sd875437, 32'sd194190, 32'sd723315, 32'sd889842, 32'sd3856050, 32'sd3779254, 32'sd2499532, 32'sd1014505, 32'sd1599202, 32'sd139055, 32'sd892221, 32'sd415270, -32'sd86730, -32'sd2368, 32'sd1050500, -32'sd567918, -32'sd1271777, -32'sd818912, -32'sd1815929, -32'sd138102, 32'sd1700361, 32'sd2216566, 32'sd629305, 32'sd1778853, 32'sd2089558, -32'sd235690, 32'sd622777, 32'sd2792527, 32'sd1223550, 32'sd11056, 32'sd1405310, 32'sd2876147, 32'sd3364542, 32'sd3357690, 32'sd1510968, -32'sd8616, 32'sd2385166, 32'sd665705, 32'sd976321, -32'sd144530, 32'sd1212250, -32'sd157539, 32'sd911263, 32'sd649863, -32'sd50848, -32'sd285576, -32'sd1196916, -32'sd1029482, 32'sd73242, -32'sd613981, 32'sd130375, 32'sd1182250, 32'sd653893, 32'sd283438, 32'sd1408778, 32'sd2728058, 32'sd2303358, -32'sd582088, 32'sd1212433, 32'sd2315032, 32'sd2482816, 32'sd1985386, 32'sd1275910, 32'sd314595, 32'sd1824645, 32'sd1935056, 32'sd289423, 32'sd1053174, 32'sd662022, 32'sd873861, 32'sd1438256, 32'sd1624838, 32'sd619677, 32'sd1051311, 32'sd937875, 32'sd945470, -32'sd1310115, -32'sd1170167, 32'sd1977578, 32'sd3024506, 32'sd1444751, 32'sd942685, 32'sd284409, 32'sd326265, -32'sd690665, -32'sd369546, 32'sd495167, -32'sd288851, -32'sd1127690, 32'sd417634, 32'sd1173599, -32'sd875303, -32'sd1863358, 32'sd910389, 32'sd503334, 32'sd1268069, 32'sd900443, 32'sd223599, -32'sd1206166, 32'sd1499897, -32'sd1704429, -32'sd141359, 32'sd872495, 32'sd464571, 32'sd473781, 32'sd2069985, 32'sd2685516, 32'sd630117, -32'sd760860, 32'sd1198381, 32'sd1019657, 32'sd322539, -32'sd1879592, -32'sd280949, 32'sd16182, -32'sd967002, -32'sd225873, 32'sd944197, -32'sd1380989, -32'sd186060, -32'sd1321487, -32'sd1096069, -32'sd1963391, -32'sd162437, 32'sd0, 32'sd567733, 32'sd129783, -32'sd655994, 32'sd542899, -32'sd157970, 32'sd318270, -32'sd1125989, 32'sd1193412, 32'sd1998396, 32'sd2138290, 32'sd224362, 32'sd602077, 32'sd1207360, 32'sd574579, -32'sd497618, -32'sd1666156, -32'sd3099107, -32'sd881593, -32'sd3074001, 32'sd599, 32'sd963194, 32'sd63987, 32'sd770989, 32'sd365269, -32'sd12510, -32'sd1618308, 32'sd575880, -32'sd928657, 32'sd528437, 32'sd514085, 32'sd31094, 32'sd708366, 32'sd2543148, 32'sd1624827, 32'sd249396, 32'sd717948, 32'sd2513246, 32'sd955532, -32'sd2056014, -32'sd1885084, -32'sd2269584, 32'sd390684, -32'sd1927770, -32'sd3090109, -32'sd650433, -32'sd1961328, -32'sd3373664, -32'sd1046893, 32'sd1027714, -32'sd1265519, 32'sd386845, 32'sd853246, 32'sd44258, -32'sd265457, 32'sd531611, -32'sd14434, -32'sd183086, 32'sd1374075, -32'sd1993027, 32'sd1369033, 32'sd17640, 32'sd2317062, 32'sd604767, 32'sd2815845, 32'sd354298, -32'sd2302060, -32'sd479350, -32'sd2539574, -32'sd2685060, -32'sd2834702, -32'sd1627311, -32'sd709673, -32'sd440740, -32'sd2404343, -32'sd2984698, -32'sd624439, -32'sd59195, 32'sd2151844, -32'sd581034, -32'sd375415, 32'sd15868, 32'sd611417, 32'sd1124177, 32'sd0, 32'sd1496131, 32'sd1720396, -32'sd595207, 32'sd2193, 32'sd1148614, 32'sd116982, 32'sd3281878, 32'sd3078051, 32'sd1121164, -32'sd2339820, -32'sd2846692, 32'sd201234, -32'sd1783912, -32'sd215971, 32'sd165975, -32'sd2346343, -32'sd806976, -32'sd1371673, -32'sd1751585, -32'sd1729087, 32'sd284919, 32'sd1941683, -32'sd653151, -32'sd2220607, -32'sd1558171, 32'sd1323808, -32'sd273037, 32'sd903276, -32'sd107536, 32'sd1373967, -32'sd486706, -32'sd1790765, -32'sd281434, 32'sd1575805, 32'sd3490526, 32'sd641104, 32'sd17562, 32'sd836876, 32'sd2054145, 32'sd1769204, 32'sd1419785, 32'sd804223, 32'sd41714, -32'sd1256247, 32'sd572803, -32'sd701914, -32'sd864298, -32'sd701182, 32'sd1278357, 32'sd870728, -32'sd18544, 32'sd828382, -32'sd1618666, 32'sd1511160, 32'sd369405, 32'sd970024, 32'sd430377, -32'sd705651, -32'sd1462360, -32'sd140973, -32'sd1238203, 32'sd2760805, 32'sd2962785, 32'sd1442992, 32'sd264565, 32'sd2746715, -32'sd427585, 32'sd1185483, -32'sd1719069, -32'sd2354191, -32'sd1354708, -32'sd1227816, -32'sd690112, -32'sd533095, 32'sd1264125, -32'sd99017, -32'sd695944, 32'sd456311, 32'sd759186, -32'sd95263, 32'sd843107, 32'sd214321, 32'sd459326, 32'sd0, 32'sd326323, -32'sd674520, 32'sd608634, -32'sd1734880, -32'sd1830644, -32'sd557777, 32'sd1408616, 32'sd1811596, -32'sd1409212, -32'sd596852, -32'sd873230, -32'sd221802, -32'sd2074920, -32'sd1098515, -32'sd2161416, -32'sd1096751, -32'sd3247675, -32'sd2933378, 32'sd497574, -32'sd1739616, -32'sd1807053, -32'sd396092, 32'sd681213, 32'sd98657, -32'sd1392612, -32'sd122764, 32'sd0, 32'sd0, 32'sd0, 32'sd333128, 32'sd550614, -32'sd623289, -32'sd2002199, 32'sd329204, 32'sd634727, -32'sd1126033, -32'sd1197103, 32'sd1125258, 32'sd194549, 32'sd260502, 32'sd2214007, 32'sd517347, -32'sd551874, -32'sd534647, 32'sd3035, -32'sd265401, -32'sd232427, -32'sd1121669, -32'sd1101014, 32'sd191069, 32'sd554864, -32'sd145345, -32'sd829531, -32'sd354319, 32'sd0, 32'sd0, 32'sd0, -32'sd1052935, 32'sd857270, 32'sd503425, -32'sd1991426, -32'sd494337, -32'sd1070698, 32'sd601568, 32'sd1123762, -32'sd52282, 32'sd572328, -32'sd327640, 32'sd1767254, 32'sd1838606, 32'sd2152936, 32'sd3390544, 32'sd1895496, 32'sd2788003, -32'sd1240778, 32'sd523794, -32'sd410393, -32'sd3714, 32'sd733810, 32'sd1118134, -32'sd237622, 32'sd135264, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd341495, -32'sd122778, -32'sd453646, -32'sd2637834, -32'sd684277, 32'sd1501917, 32'sd1497760, -32'sd293238, 32'sd2165587, 32'sd1289008, -32'sd920334, 32'sd242584, -32'sd744459, -32'sd1508651, -32'sd1164126, 32'sd60188, -32'sd1444048, 32'sd361407, 32'sd570044, 32'sd95342, -32'sd1334129, -32'sd591563, -32'sd449672, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd334094, 32'sd564764, -32'sd1308055, -32'sd721802, -32'sd826745, -32'sd1222247, -32'sd463945, -32'sd1393016, -32'sd1313042, -32'sd500823, -32'sd844365, 32'sd1229350, 32'sd111877, -32'sd171519, -32'sd1197508, -32'sd310726, 32'sd1075172, 32'sd1414118, -32'sd939282, -32'sd49797, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1188605, -32'sd537874, 32'sd570389, 32'sd1054405, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd326647, 32'sd1316580, 32'sd793127, 32'sd76470, 32'sd1795311, 32'sd423794, 32'sd1760860, 32'sd440188, -32'sd742843, 32'sd143009, -32'sd336092, 32'sd1004967, 32'sd1396737, 32'sd827002, 32'sd284327, 32'sd1099593, 32'sd454249, 32'sd466411, 32'sd608588, -32'sd292819, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd675892, 32'sd730424, -32'sd1880254, -32'sd626703, 32'sd678384, 32'sd797114, -32'sd1015879, 32'sd54934, 32'sd587155, 32'sd493849, 32'sd1033433, 32'sd1285040, 32'sd16667, 32'sd28351, -32'sd308767, 32'sd939841, 32'sd777339, 32'sd550984, 32'sd413967, -32'sd195528, -32'sd299255, -32'sd1684580, 32'sd2188502, 32'sd794403, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd576130, -32'sd468939, 32'sd455878, -32'sd2181620, -32'sd396422, -32'sd49327, -32'sd517488, -32'sd172224, 32'sd1378646, 32'sd964353, 32'sd972851, 32'sd735736, 32'sd1028617, 32'sd1349560, 32'sd795816, -32'sd1206314, -32'sd469550, -32'sd482278, -32'sd1909230, -32'sd1797140, -32'sd1110521, -32'sd1250931, -32'sd1346557, -32'sd89977, -32'sd272629, 32'sd0, 32'sd0, 32'sd460674, 32'sd1192241, 32'sd377439, 32'sd190466, -32'sd10897, -32'sd1013938, 32'sd869583, 32'sd1505213, 32'sd525755, 32'sd410349, 32'sd586633, 32'sd2067068, 32'sd993395, 32'sd2688866, 32'sd1066694, -32'sd408561, -32'sd1393099, -32'sd650337, -32'sd2082401, -32'sd3594565, -32'sd2752515, -32'sd18165, -32'sd1965562, -32'sd774846, 32'sd129849, -32'sd1030814, 32'sd377425, 32'sd0, 32'sd334929, 32'sd800372, -32'sd126297, 32'sd194429, 32'sd608205, 32'sd1247604, -32'sd100868, -32'sd1155579, -32'sd1130956, -32'sd56111, 32'sd1155173, 32'sd1407590, 32'sd2707751, 32'sd1689918, 32'sd1704048, -32'sd161821, -32'sd1563907, 32'sd716943, -32'sd5494, -32'sd946229, -32'sd4091521, -32'sd1580851, -32'sd518731, -32'sd120751, -32'sd228978, -32'sd190462, 32'sd796755, 32'sd0, 32'sd311223, -32'sd305848, -32'sd1236336, -32'sd132557, 32'sd1236555, -32'sd722994, -32'sd345376, -32'sd1628114, -32'sd1468798, -32'sd1578470, -32'sd1385495, 32'sd375189, 32'sd354954, 32'sd314186, 32'sd684854, 32'sd152791, 32'sd741227, -32'sd453320, 32'sd233529, -32'sd724259, -32'sd1503984, -32'sd726395, -32'sd1436080, -32'sd872814, 32'sd1283899, -32'sd829360, -32'sd777890, 32'sd485524, -32'sd54862, 32'sd649810, 32'sd349954, -32'sd245098, -32'sd1682615, -32'sd978653, -32'sd846747, -32'sd3429598, -32'sd499585, -32'sd51287, 32'sd179180, -32'sd1169071, -32'sd267375, 32'sd1876883, 32'sd721828, 32'sd2238838, 32'sd972921, -32'sd1091165, 32'sd565705, 32'sd257984, 32'sd408159, -32'sd1435245, -32'sd1236643, -32'sd1681848, 32'sd493558, -32'sd293450, -32'sd344671, 32'sd1075888, -32'sd91177, 32'sd1413231, 32'sd343536, 32'sd1427363, -32'sd729311, -32'sd18265, -32'sd871820, -32'sd1694447, -32'sd1466886, -32'sd342269, -32'sd3031529, -32'sd1723166, -32'sd1231801, 32'sd2197676, 32'sd2099235, 32'sd1661859, 32'sd1684794, -32'sd150770, -32'sd283410, -32'sd685946, -32'sd1538630, -32'sd551222, -32'sd2219674, -32'sd1859913, -32'sd1545340, -32'sd1120679, 32'sd1681521, 32'sd1914719, 32'sd97257, -32'sd279182, -32'sd1256565, -32'sd681558, -32'sd1399925, -32'sd851219, -32'sd723604, -32'sd1096242, -32'sd838051, -32'sd126708, -32'sd2194151, -32'sd1060014, 32'sd1720327, 32'sd3562186, 32'sd2689808, 32'sd2278459, 32'sd2228082, 32'sd48462, 32'sd851920, -32'sd2488644, -32'sd2842089, -32'sd465642, -32'sd1510717, -32'sd907008, -32'sd1313684, -32'sd892586, 32'sd769977, 32'sd203009, 32'sd1290043, 32'sd1284036, -32'sd228636, -32'sd1775564, -32'sd2220090, -32'sd721829, -32'sd690300, 32'sd624271, -32'sd294930, 32'sd194528, -32'sd1624779, 32'sd1705702, 32'sd1773966, 32'sd3366085, 32'sd3588728, 32'sd2165377, -32'sd388482, -32'sd2549322, -32'sd1470040, -32'sd2437379, -32'sd1590064, 32'sd612657, -32'sd2170934, -32'sd1266641, 32'sd179577, 32'sd655550, -32'sd922656, 32'sd850470, 32'sd46972, 32'sd2510986, 32'sd446747, -32'sd138997, -32'sd2333857, 32'sd308327, 32'sd215775, 32'sd58370, -32'sd627496, 32'sd1199159, -32'sd825631, 32'sd2281518, 32'sd1810409, 32'sd1503880, 32'sd2184896, 32'sd1330610, -32'sd1002513, -32'sd1275144, -32'sd1594031, -32'sd304923, 32'sd54949, 32'sd334051, -32'sd285285, -32'sd1303904, 32'sd2787095, -32'sd747798, 32'sd575508, 32'sd728228, 32'sd2418815, 32'sd1743378, 32'sd147396, -32'sd1517192, -32'sd2131483, 32'sd896560, 32'sd134503, 32'sd406987, 32'sd2977803, 32'sd2768696, -32'sd856350, 32'sd943993, 32'sd2422398, 32'sd1838407, 32'sd1377839, 32'sd879542, -32'sd740552, -32'sd1316169, -32'sd2662940, -32'sd1415352, -32'sd1901731, -32'sd2106077, -32'sd251797, -32'sd22459, -32'sd49049, -32'sd694730, -32'sd300681, 32'sd133605, 32'sd2477553, 32'sd1666135, -32'sd961461, 32'sd845110, -32'sd1557577, 32'sd2770141, 32'sd1427949, -32'sd2349601, 32'sd252101, 32'sd1417476, -32'sd308158, -32'sd285217, 32'sd1130872, 32'sd2498766, 32'sd2744770, 32'sd319607, -32'sd50210, -32'sd2240623, -32'sd2985538, -32'sd51010, -32'sd1673099, -32'sd370303, 32'sd343147, 32'sd844216, 32'sd564017, -32'sd212176, 32'sd198760, -32'sd38636, 32'sd251133, 32'sd1184151, -32'sd219109, 32'sd289989, -32'sd591645, -32'sd57251, -32'sd417244, -32'sd1750589, -32'sd1894792, -32'sd2243742, -32'sd2809450, 32'sd363371, 32'sd948632, 32'sd3365430, 32'sd3493853, 32'sd522232, 32'sd697839, -32'sd1953486, -32'sd1460916, 32'sd861160, 32'sd904963, -32'sd176288, 32'sd1784255, 32'sd367854, 32'sd1152521, -32'sd1896316, -32'sd458805, -32'sd142658, 32'sd1530623, 32'sd227081, -32'sd1779665, 32'sd2142689, -32'sd596553, -32'sd684576, 32'sd953366, -32'sd387759, -32'sd557430, -32'sd2558075, -32'sd2036974, -32'sd1856251, 32'sd1707673, 32'sd1968322, -32'sd425416, 32'sd1238763, -32'sd1556681, -32'sd1781542, -32'sd1353903, -32'sd1142029, -32'sd931682, 32'sd1385403, 32'sd1457087, 32'sd1157827, 32'sd1972571, -32'sd1543378, 32'sd892969, 32'sd411232, 32'sd990136, 32'sd1909797, -32'sd143975, 32'sd1503754, -32'sd542205, 32'sd456018, 32'sd472213, -32'sd119065, -32'sd1492761, -32'sd1546501, -32'sd95523, -32'sd499955, 32'sd2344158, 32'sd840932, 32'sd218207, -32'sd870538, -32'sd1644943, -32'sd2013045, -32'sd2621040, -32'sd1238227, 32'sd246663, -32'sd944427, 32'sd1314569, 32'sd585988, -32'sd1441682, -32'sd526937, 32'sd93365, 32'sd0, 32'sd739453, -32'sd51492, 32'sd687287, 32'sd154979, -32'sd1266739, -32'sd1018968, 32'sd234418, 32'sd143216, -32'sd213230, -32'sd1183193, -32'sd341816, -32'sd2123169, 32'sd1359279, 32'sd302503, 32'sd1228380, -32'sd1593227, -32'sd1495021, -32'sd1191166, -32'sd197420, -32'sd483603, 32'sd16484, 32'sd238139, -32'sd92427, 32'sd1838655, -32'sd67917, 32'sd8214, 32'sd655794, 32'sd693182, 32'sd1096708, 32'sd85616, -32'sd169960, -32'sd321069, 32'sd575509, 32'sd823082, -32'sd453707, 32'sd1654963, -32'sd1283493, -32'sd145737, -32'sd700360, -32'sd2614412, 32'sd390445, 32'sd738462, -32'sd115581, -32'sd925106, -32'sd1108265, -32'sd1531861, -32'sd368729, -32'sd1675, -32'sd287306, -32'sd773591, 32'sd1612184, 32'sd442545, 32'sd1265235, 32'sd969357, 32'sd1418395, 32'sd502916, 32'sd179966, 32'sd627176, -32'sd1599704, 32'sd1064856, 32'sd572347, -32'sd993314, 32'sd1499043, -32'sd613393, -32'sd1205681, -32'sd1700960, -32'sd2369508, -32'sd1448904, 32'sd225101, 32'sd823984, -32'sd399758, -32'sd1535321, -32'sd987783, -32'sd1678598, 32'sd1209732, 32'sd473136, -32'sd1693957, -32'sd312972, -32'sd779683, -32'sd1637092, 32'sd1637904, 32'sd414401, 32'sd1435459, 32'sd0, -32'sd52524, 32'sd320276, -32'sd1110215, -32'sd654443, -32'sd752011, -32'sd1535115, -32'sd148500, 32'sd699546, -32'sd115217, -32'sd1320047, -32'sd988763, 32'sd1400435, -32'sd1577405, -32'sd205444, -32'sd1715857, -32'sd560257, 32'sd195273, -32'sd563031, 32'sd472210, -32'sd1194892, -32'sd310275, -32'sd1493602, 32'sd1570810, 32'sd769053, 32'sd2011188, 32'sd992253, 32'sd1543843, 32'sd1421838, 32'sd704898, 32'sd1117691, 32'sd794867, -32'sd585537, -32'sd2507148, -32'sd1756749, -32'sd706365, 32'sd1126029, 32'sd535285, 32'sd578165, -32'sd465542, 32'sd335801, -32'sd501364, -32'sd1779065, -32'sd545614, -32'sd1436195, -32'sd2016861, -32'sd1707779, 32'sd85664, 32'sd634375, -32'sd123330, 32'sd209613, -32'sd1482563, -32'sd37893, 32'sd1243259, 32'sd758135, 32'sd842579, 32'sd638929, 32'sd1240023, 32'sd574563, 32'sd1937634, 32'sd1159570, -32'sd1221838, 32'sd148485, 32'sd299289, -32'sd540587, 32'sd2130980, 32'sd2177095, 32'sd599421, -32'sd2189536, -32'sd839233, 32'sd2315754, 32'sd1202328, -32'sd1172342, 32'sd856640, 32'sd1544446, 32'sd1383812, 32'sd1842403, -32'sd52019, -32'sd889544, -32'sd1432253, -32'sd1240689, 32'sd455996, 32'sd880250, 32'sd1488975, 32'sd0, 32'sd751289, -32'sd334039, 32'sd1780570, 32'sd111308, -32'sd1521104, -32'sd1645082, 32'sd137450, 32'sd87537, 32'sd826181, 32'sd1346214, 32'sd78493, 32'sd253793, 32'sd535326, -32'sd152846, 32'sd2179320, -32'sd1148464, 32'sd1551283, 32'sd368039, 32'sd612361, 32'sd1193103, 32'sd536266, 32'sd569632, 32'sd1029198, -32'sd1600775, -32'sd644818, 32'sd19343, 32'sd0, 32'sd0, 32'sd0, -32'sd22621, 32'sd2239709, 32'sd1126936, -32'sd679801, -32'sd1574125, -32'sd1535844, 32'sd1015506, 32'sd561590, -32'sd453349, -32'sd817637, -32'sd1092450, -32'sd1553600, 32'sd89372, 32'sd1278387, -32'sd416712, 32'sd112269, 32'sd167076, 32'sd1504005, 32'sd445007, 32'sd1401741, 32'sd1088264, -32'sd307519, 32'sd1213970, -32'sd949096, 32'sd855464, 32'sd0, 32'sd0, 32'sd0, 32'sd776058, -32'sd1424493, 32'sd712262, -32'sd12762, -32'sd2062705, 32'sd797437, 32'sd3727094, 32'sd1938944, 32'sd1658937, -32'sd902490, -32'sd1821882, 32'sd207921, 32'sd867351, 32'sd1535221, -32'sd705096, 32'sd855019, -32'sd2737680, -32'sd1145240, 32'sd2117800, -32'sd265784, -32'sd774650, 32'sd243465, 32'sd388629, -32'sd421257, 32'sd209063, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd755304, -32'sd1389863, 32'sd483403, 32'sd1921330, 32'sd2757386, 32'sd1587760, 32'sd933836, 32'sd417498, 32'sd1269820, 32'sd1384926, -32'sd2251016, -32'sd11646, -32'sd493648, -32'sd550168, 32'sd113318, -32'sd1686272, -32'sd113658, 32'sd621258, 32'sd1182425, -32'sd1802842, 32'sd1067206, 32'sd2024908, 32'sd1439687, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1956563, -32'sd661166, 32'sd1134523, -32'sd974093, 32'sd537028, 32'sd455554, 32'sd77496, 32'sd772725, 32'sd1623087, 32'sd365303, 32'sd443910, 32'sd573920, 32'sd933384, 32'sd595504, -32'sd31594, 32'sd752729, -32'sd505501, 32'sd2565179, 32'sd1784273, 32'sd2554705, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd199122, -32'sd864578, -32'sd421380, -32'sd68504, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd720239, -32'sd193562, 32'sd378086, 32'sd14385, 32'sd886839, -32'sd159348, -32'sd701141, -32'sd1220573, 32'sd930476, -32'sd601652, 32'sd443339, -32'sd515724, 32'sd15889, -32'sd730115, -32'sd1964854, 32'sd934049, 32'sd152208, 32'sd540776, -32'sd767058, 32'sd663290, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd174457, 32'sd376569, 32'sd726762, -32'sd785864, -32'sd373905, -32'sd759085, -32'sd910893, -32'sd19629, -32'sd1933051, -32'sd2079164, -32'sd2110340, -32'sd982730, -32'sd964747, -32'sd193986, -32'sd359267, 32'sd77122, 32'sd442517, 32'sd1564359, 32'sd862188, -32'sd1290011, -32'sd1706861, -32'sd1150064, 32'sd486728, -32'sd694578, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd351988, -32'sd470449, 32'sd1509171, 32'sd1676526, -32'sd870230, 32'sd694163, -32'sd682780, -32'sd1762653, 32'sd140438, 32'sd105260, 32'sd203065, -32'sd1267674, 32'sd1570027, -32'sd667820, 32'sd1749665, 32'sd824409, 32'sd582929, 32'sd85052, 32'sd1589321, 32'sd43429, 32'sd613541, 32'sd113121, 32'sd26030, 32'sd1390191, -32'sd54383, 32'sd0, 32'sd0, -32'sd165681, -32'sd774376, 32'sd462460, 32'sd495583, 32'sd66948, 32'sd210283, -32'sd365927, -32'sd441634, -32'sd1337682, -32'sd1706658, -32'sd1077478, 32'sd780135, 32'sd1353449, 32'sd994371, -32'sd649205, 32'sd1654682, -32'sd755863, -32'sd2460919, -32'sd907842, -32'sd2150157, -32'sd2319583, 32'sd38961, 32'sd709821, 32'sd1074357, 32'sd1288643, 32'sd327495, 32'sd722063, 32'sd0, 32'sd169954, 32'sd1775475, 32'sd2550945, 32'sd902858, -32'sd170661, -32'sd624136, -32'sd640542, 32'sd414140, 32'sd446104, 32'sd1008182, -32'sd2522265, -32'sd1661799, -32'sd161891, 32'sd436486, 32'sd1458223, -32'sd421860, -32'sd371709, -32'sd823858, 32'sd586502, 32'sd57912, -32'sd1659976, 32'sd302604, -32'sd721556, -32'sd269209, -32'sd349380, 32'sd816138, -32'sd1007153, 32'sd0, 32'sd325460, 32'sd102401, 32'sd267642, 32'sd478293, 32'sd65376, -32'sd363908, -32'sd494167, -32'sd233467, -32'sd372119, -32'sd1262447, -32'sd2229422, -32'sd2053023, 32'sd1491161, 32'sd2214603, 32'sd3907117, 32'sd2949820, 32'sd2156860, 32'sd3250530, 32'sd1210144, -32'sd469538, 32'sd2269385, -32'sd1094906, 32'sd782517, 32'sd250901, 32'sd194365, -32'sd295839, 32'sd829815, 32'sd190388, -32'sd692389, -32'sd382927, -32'sd1686805, -32'sd962839, -32'sd1266929, -32'sd70138, 32'sd1238250, 32'sd88838, -32'sd1147109, -32'sd1735696, 32'sd343317, 32'sd1466857, -32'sd783614, 32'sd2090913, 32'sd4041190, 32'sd2323858, 32'sd2449129, 32'sd4274388, 32'sd1198282, 32'sd2426543, 32'sd2093201, 32'sd204119, -32'sd2657206, 32'sd1482145, 32'sd2428498, 32'sd991771, -32'sd806828, 32'sd819049, 32'sd363085, -32'sd413943, -32'sd820807, -32'sd299009, 32'sd1637371, 32'sd940219, -32'sd937275, -32'sd2185105, -32'sd94437, 32'sd360257, 32'sd1291317, -32'sd793704, 32'sd1465625, 32'sd309012, 32'sd2427076, 32'sd4468896, 32'sd2365097, 32'sd4271559, 32'sd973980, 32'sd1526087, 32'sd1960061, -32'sd1112737, 32'sd515387, 32'sd2250928, 32'sd2129438, 32'sd1245402, 32'sd767497, -32'sd114478, 32'sd1123900, 32'sd1171483, -32'sd124981, 32'sd780044, -32'sd70764, -32'sd1560978, -32'sd232498, -32'sd125905, 32'sd1544896, 32'sd721459, 32'sd803824, 32'sd723578, 32'sd632986, 32'sd3192591, 32'sd2376255, 32'sd470520, 32'sd3556702, 32'sd1511942, 32'sd2188301, 32'sd2239398, 32'sd109561, -32'sd1470096, -32'sd499249, 32'sd1725839, 32'sd1550157, 32'sd458217, 32'sd1219591, -32'sd345502, -32'sd90029, 32'sd1073592, 32'sd209120, 32'sd764924, -32'sd355307, 32'sd916031, 32'sd367426, 32'sd508265, -32'sd861695, -32'sd357511, 32'sd29659, -32'sd1491596, 32'sd323003, 32'sd169895, -32'sd1090724, -32'sd591612, -32'sd1393661, 32'sd141366, 32'sd832857, 32'sd265412, -32'sd115406, -32'sd296186, -32'sd640742, -32'sd809295, 32'sd835515, 32'sd801902, -32'sd997743, -32'sd103973, 32'sd1113711, 32'sd1554862, 32'sd1405069, 32'sd214774, -32'sd1383194, 32'sd509665, 32'sd1412681, 32'sd965718, -32'sd1334735, -32'sd435169, 32'sd1913886, -32'sd2785513, 32'sd317023, 32'sd2654157, 32'sd186223, -32'sd2224140, -32'sd399075, -32'sd933071, -32'sd1450925, 32'sd1237920, -32'sd1915666, -32'sd2075543, -32'sd32930, 32'sd343085, -32'sd458670, -32'sd1575347, -32'sd1765302, 32'sd312471, 32'sd206927, -32'sd714877, 32'sd740492, 32'sd143851, -32'sd1543238, -32'sd2841970, -32'sd1226625, -32'sd1464602, -32'sd265906, -32'sd656682, -32'sd860434, -32'sd2659724, -32'sd1395205, -32'sd1030405, 32'sd2272211, -32'sd980017, 32'sd994672, 32'sd507539, -32'sd213216, 32'sd154135, -32'sd951168, -32'sd1099367, -32'sd1452844, -32'sd1165361, -32'sd1665470, -32'sd2474970, -32'sd1070230, -32'sd374544, -32'sd824915, 32'sd85821, -32'sd1287291, 32'sd843686, -32'sd763874, -32'sd264991, -32'sd60863, 32'sd709005, -32'sd578385, -32'sd2933255, -32'sd2162671, -32'sd1978039, -32'sd2477725, 32'sd777996, -32'sd455468, -32'sd1718445, -32'sd922676, 32'sd581778, 32'sd96191, -32'sd1464049, -32'sd332132, -32'sd2941314, -32'sd2219111, -32'sd1391025, -32'sd94787, -32'sd34568, -32'sd1029243, 32'sd419924, -32'sd70927, -32'sd124831, 32'sd462898, -32'sd1300541, -32'sd1057379, 32'sd970845, 32'sd244740, -32'sd2047946, -32'sd2872337, -32'sd2131429, -32'sd4109288, -32'sd2607596, -32'sd1166369, -32'sd767002, 32'sd1013263, 32'sd215659, -32'sd841312, 32'sd1957363, 32'sd1389731, 32'sd482432, -32'sd1997268, -32'sd1551626, -32'sd3988280, -32'sd1364094, 32'sd1051548, 32'sd73909, -32'sd133604, 32'sd883867, 32'sd11426, 32'sd1154769, -32'sd1026629, -32'sd1293305, 32'sd1075908, -32'sd1302624, 32'sd272635, -32'sd1270650, -32'sd3330346, -32'sd632881, -32'sd2769949, -32'sd967512, -32'sd614079, -32'sd1018857, 32'sd1685250, -32'sd111500, -32'sd1761503, 32'sd49549, -32'sd1078027, -32'sd381320, -32'sd2181785, -32'sd2703034, -32'sd2394008, -32'sd3147, 32'sd121424, -32'sd826039, -32'sd464115, 32'sd828412, -32'sd489974, 32'sd354949, 32'sd595231, -32'sd1348813, -32'sd1637250, -32'sd725666, -32'sd1049033, 32'sd1189619, 32'sd24291, -32'sd1018092, -32'sd2548191, -32'sd742032, -32'sd1833681, -32'sd2223710, -32'sd130061, -32'sd581788, -32'sd583517, 32'sd370675, 32'sd10454, -32'sd1294771, -32'sd3873604, -32'sd1482006, -32'sd1271682, 32'sd1810481, 32'sd1103967, -32'sd2114119, -32'sd1125261, 32'sd0, 32'sd528220, 32'sd1165033, 32'sd960515, -32'sd1255001, -32'sd2174772, -32'sd1801829, 32'sd763644, 32'sd1373853, -32'sd741145, -32'sd2366936, -32'sd1468538, -32'sd277252, -32'sd447765, -32'sd2163495, 32'sd306602, -32'sd840123, 32'sd1774518, 32'sd1567281, 32'sd652407, -32'sd2077298, -32'sd3357633, -32'sd2316707, -32'sd2322266, 32'sd533452, 32'sd1986085, -32'sd593924, -32'sd350007, -32'sd801417, -32'sd919094, -32'sd360929, -32'sd1773368, -32'sd2966886, 32'sd198594, 32'sd594197, 32'sd1018750, 32'sd1317179, -32'sd2162, -32'sd499464, -32'sd330438, 32'sd1711937, 32'sd706112, -32'sd981782, 32'sd541647, 32'sd2003043, 32'sd3940554, 32'sd423155, -32'sd703138, -32'sd3071489, -32'sd1170833, -32'sd755640, -32'sd655058, 32'sd1124110, -32'sd159455, -32'sd308087, -32'sd1022771, 32'sd144676, 32'sd921911, 32'sd1668721, -32'sd2163119, 32'sd566243, 32'sd1473605, 32'sd1929416, -32'sd544592, -32'sd1583162, -32'sd831910, 32'sd645009, 32'sd549451, 32'sd2641761, -32'sd1117326, 32'sd488929, -32'sd150836, 32'sd349929, 32'sd2246258, 32'sd1044533, -32'sd1269673, -32'sd2270868, -32'sd1909111, -32'sd1061920, -32'sd2128226, 32'sd1701910, 32'sd1103372, -32'sd884494, -32'sd675255, 32'sd0, -32'sd315987, 32'sd828378, -32'sd433537, 32'sd376800, 32'sd242842, 32'sd1767984, 32'sd1042291, -32'sd239403, -32'sd2070633, 32'sd618460, 32'sd456542, -32'sd860249, -32'sd1343040, 32'sd464374, -32'sd113917, 32'sd1587881, 32'sd3845737, -32'sd118245, -32'sd374403, -32'sd2854064, -32'sd974656, -32'sd649751, 32'sd299499, 32'sd425756, -32'sd739181, -32'sd542875, 32'sd329931, -32'sd984964, -32'sd950200, 32'sd120096, -32'sd933265, -32'sd1090815, -32'sd403682, 32'sd502192, -32'sd774318, -32'sd2684777, -32'sd2238563, -32'sd972454, -32'sd997356, -32'sd1100757, 32'sd330480, -32'sd212540, -32'sd197667, 32'sd1376264, 32'sd1736154, -32'sd2319577, -32'sd2083796, -32'sd2299980, -32'sd1670272, -32'sd2299885, -32'sd743341, -32'sd26661, 32'sd653329, -32'sd702964, 32'sd560239, -32'sd187129, -32'sd772635, -32'sd205231, -32'sd309009, -32'sd622544, -32'sd2313269, 32'sd1562397, -32'sd913868, -32'sd1597891, -32'sd2194011, 32'sd497526, -32'sd90193, 32'sd2685773, 32'sd1588979, 32'sd2317548, 32'sd399240, -32'sd1274346, 32'sd339067, -32'sd2668837, -32'sd3190087, -32'sd2811767, -32'sd2704202, -32'sd3398477, -32'sd1380279, -32'sd1012381, -32'sd626076, 32'sd22765, 32'sd199718, 32'sd0, 32'sd506295, 32'sd684406, -32'sd1691417, -32'sd723950, -32'sd1675980, -32'sd2438319, -32'sd1244149, -32'sd2805701, -32'sd2312143, -32'sd649553, 32'sd576100, 32'sd51711, 32'sd2305406, -32'sd821070, -32'sd1921077, -32'sd735774, -32'sd1513842, -32'sd1932181, -32'sd3117377, -32'sd1382057, -32'sd1319407, 32'sd1270165, 32'sd737569, -32'sd584963, 32'sd566888, -32'sd1302304, 32'sd0, 32'sd0, 32'sd0, 32'sd537265, 32'sd37371, -32'sd648582, 32'sd2205182, 32'sd864038, -32'sd1217430, -32'sd379556, -32'sd997731, 32'sd68620, 32'sd1683277, 32'sd2605359, 32'sd1661202, -32'sd31846, 32'sd238828, 32'sd612789, 32'sd28869, -32'sd3585085, -32'sd2217412, -32'sd354183, -32'sd4453807, -32'sd1601296, -32'sd203702, -32'sd1713308, 32'sd394556, -32'sd479795, 32'sd0, 32'sd0, 32'sd0, 32'sd879408, -32'sd737781, -32'sd1639353, 32'sd831647, -32'sd289501, 32'sd1826780, 32'sd1814061, -32'sd1375835, 32'sd1790356, -32'sd317025, 32'sd2062449, 32'sd675601, 32'sd1401473, -32'sd361466, -32'sd723253, 32'sd1261343, -32'sd1476628, -32'sd683722, -32'sd1818446, -32'sd664278, 32'sd1612503, -32'sd1198456, 32'sd201052, 32'sd718217, 32'sd269849, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd79428, -32'sd1147368, 32'sd103540, -32'sd1473174, 32'sd1454984, 32'sd1041463, 32'sd3203064, 32'sd1676511, 32'sd423869, 32'sd564323, 32'sd135839, -32'sd189168, 32'sd1374096, -32'sd397208, 32'sd790055, 32'sd1407400, 32'sd544041, -32'sd811349, -32'sd922205, 32'sd1263109, 32'sd165956, -32'sd1564334, -32'sd452284, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd706192, 32'sd86634, -32'sd205004, 32'sd1327674, -32'sd869626, 32'sd1144833, 32'sd1241723, 32'sd783385, -32'sd1553191, -32'sd953142, 32'sd600195, 32'sd598776, 32'sd1663214, 32'sd2150417, 32'sd485060, -32'sd209882, -32'sd567538, -32'sd425783, -32'sd611416, -32'sd435730, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd857091, 32'sd783414, -32'sd579532, -32'sd1343445, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2421677, 32'sd103186, 32'sd1266518, -32'sd237628, 32'sd1393482, 32'sd70412, 32'sd704654, 32'sd335017, 32'sd347941, 32'sd1254638, 32'sd1443572, 32'sd824669, 32'sd119427, 32'sd1023646, 32'sd393854, -32'sd257146, 32'sd1372760, 32'sd523164, 32'sd777347, 32'sd91257, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1131219, 32'sd83887, 32'sd375890, 32'sd1104500, -32'sd843207, -32'sd465054, -32'sd593619, 32'sd157159, -32'sd1974027, -32'sd763337, -32'sd433034, 32'sd1688067, 32'sd1641928, 32'sd376570, -32'sd608821, -32'sd1898387, 32'sd1881562, 32'sd316374, 32'sd1884786, 32'sd1572439, 32'sd1941872, -32'sd91613, -32'sd305576, 32'sd1100839, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1284902, 32'sd1296246, 32'sd458279, -32'sd1079688, 32'sd232064, -32'sd1457702, 32'sd3032606, 32'sd1458462, 32'sd1575899, -32'sd803918, -32'sd469067, -32'sd299696, 32'sd201806, 32'sd1286180, -32'sd65609, -32'sd976817, 32'sd1963099, 32'sd2334735, 32'sd2067707, 32'sd24636, -32'sd765065, -32'sd1741879, -32'sd1756011, 32'sd8191, 32'sd1266013, 32'sd0, 32'sd0, 32'sd1046735, 32'sd171355, 32'sd614136, -32'sd1198377, 32'sd573869, -32'sd136380, -32'sd1325004, 32'sd1063027, 32'sd1337822, 32'sd928556, 32'sd1797778, 32'sd55344, 32'sd1067957, 32'sd1957633, 32'sd2691918, 32'sd1333042, -32'sd973491, 32'sd1403140, -32'sd237332, 32'sd1314662, 32'sd213658, -32'sd1779959, 32'sd448140, -32'sd621405, 32'sd460908, 32'sd1302883, 32'sd244663, 32'sd0, 32'sd155649, 32'sd582587, 32'sd164214, 32'sd5538, -32'sd702473, -32'sd1781252, -32'sd393228, -32'sd77555, 32'sd259595, -32'sd31117, -32'sd202621, -32'sd2514501, -32'sd1895288, -32'sd1253081, 32'sd1109498, -32'sd62183, -32'sd100687, -32'sd282947, 32'sd807001, 32'sd1030144, -32'sd940524, -32'sd1598918, -32'sd216461, 32'sd836277, 32'sd230747, 32'sd1061221, -32'sd931997, 32'sd0, 32'sd64046, -32'sd418376, 32'sd1528635, 32'sd874908, 32'sd1403738, 32'sd1903244, -32'sd763511, 32'sd390565, -32'sd2026242, -32'sd1121220, -32'sd942399, -32'sd427841, -32'sd1034454, 32'sd24654, 32'sd644418, 32'sd648100, -32'sd1638903, -32'sd1060812, -32'sd471568, -32'sd97694, -32'sd430622, -32'sd1781107, 32'sd338435, 32'sd1147826, 32'sd295714, 32'sd809003, 32'sd882069, 32'sd177500, 32'sd1053473, 32'sd1125337, 32'sd186962, -32'sd1309540, -32'sd1738733, -32'sd1258208, -32'sd644033, 32'sd741406, -32'sd1827570, -32'sd836503, 32'sd129280, 32'sd1430511, 32'sd637504, 32'sd2659515, 32'sd775572, -32'sd1054423, 32'sd230525, -32'sd3019973, -32'sd3540827, -32'sd1923625, -32'sd1625106, -32'sd1079962, -32'sd2800919, -32'sd1993634, 32'sd225460, 32'sd77650, -32'sd1308836, 32'sd431764, -32'sd698367, 32'sd945202, 32'sd1405975, -32'sd1168864, -32'sd1553430, -32'sd2421286, -32'sd1820841, -32'sd226919, -32'sd719838, -32'sd2208715, -32'sd241452, 32'sd360400, -32'sd501117, -32'sd484937, -32'sd1575189, -32'sd2391623, -32'sd1277203, -32'sd2926083, -32'sd2375548, -32'sd2130042, 32'sd246644, -32'sd496819, -32'sd339899, -32'sd364533, 32'sd670129, 32'sd1470965, 32'sd937906, 32'sd647546, -32'sd2122837, -32'sd539105, 32'sd1454120, -32'sd308296, -32'sd2867029, -32'sd246870, -32'sd843013, -32'sd1276542, -32'sd1217885, -32'sd846997, -32'sd1187501, 32'sd276584, 32'sd935963, 32'sd160626, -32'sd807639, 32'sd1306637, 32'sd2051026, -32'sd36630, -32'sd262910, -32'sd413917, 32'sd1194055, 32'sd2010887, 32'sd48416, 32'sd2008902, 32'sd1502353, -32'sd453663, -32'sd182504, 32'sd199010, -32'sd1672787, -32'sd790636, 32'sd332843, 32'sd819025, -32'sd481241, -32'sd1916609, -32'sd876150, -32'sd1144412, -32'sd1879391, -32'sd1823799, -32'sd1015954, 32'sd1568416, 32'sd2291123, 32'sd2269700, 32'sd1168855, 32'sd1116399, 32'sd2641405, 32'sd1599834, 32'sd952026, 32'sd342968, -32'sd371837, -32'sd894238, 32'sd2475825, 32'sd2146653, -32'sd784720, 32'sd1167321, 32'sd1405003, -32'sd842955, 32'sd573642, 32'sd1091442, 32'sd326573, 32'sd480773, -32'sd2002863, -32'sd1360476, -32'sd1983479, -32'sd895395, 32'sd88058, 32'sd1535392, -32'sd1179221, 32'sd242345, 32'sd631534, 32'sd684742, -32'sd936445, 32'sd1203574, 32'sd4454121, 32'sd856094, 32'sd1420065, 32'sd18201, -32'sd376666, -32'sd628786, 32'sd730850, -32'sd974491, -32'sd179768, 32'sd145228, 32'sd1176552, 32'sd582759, 32'sd1022443, -32'sd373105, 32'sd1766568, 32'sd41645, -32'sd294964, 32'sd269795, -32'sd343468, -32'sd891866, 32'sd59556, -32'sd1161492, -32'sd1928202, -32'sd648981, -32'sd358134, 32'sd929768, -32'sd1299236, 32'sd491776, -32'sd103928, -32'sd1547785, -32'sd17882, -32'sd1215127, -32'sd1683923, 32'sd1001643, 32'sd316698, -32'sd1703026, -32'sd2354040, -32'sd724632, 32'sd38804, 32'sd1364460, 32'sd346380, -32'sd307397, 32'sd1142111, -32'sd162486, -32'sd1953065, -32'sd1126546, 32'sd223135, -32'sd750966, 32'sd698923, -32'sd208027, -32'sd624623, -32'sd2060349, -32'sd1085366, 32'sd192573, 32'sd720603, 32'sd440021, -32'sd3255104, -32'sd2361284, -32'sd48851, 32'sd389763, -32'sd715002, 32'sd479874, 32'sd2121472, -32'sd3242467, -32'sd1216136, -32'sd161863, 32'sd400035, 32'sd1912011, 32'sd488126, -32'sd974627, 32'sd1378371, 32'sd1388691, -32'sd2596158, -32'sd2521360, -32'sd470753, -32'sd1028252, 32'sd2186980, -32'sd775861, -32'sd2736044, -32'sd1613940, -32'sd962741, -32'sd601241, -32'sd738537, -32'sd937144, -32'sd4041586, -32'sd3848781, -32'sd1235594, -32'sd188323, 32'sd1032583, 32'sd1247569, -32'sd28304, -32'sd618633, -32'sd973553, 32'sd291807, -32'sd688992, 32'sd805448, 32'sd893226, 32'sd1516923, 32'sd755949, 32'sd1667291, -32'sd209919, -32'sd509731, -32'sd1533478, 32'sd368410, 32'sd867898, -32'sd1249753, 32'sd636357, -32'sd629335, 32'sd330848, 32'sd307517, -32'sd2799305, -32'sd1383081, -32'sd2855299, -32'sd1383949, -32'sd975212, 32'sd552997, 32'sd684189, -32'sd426139, -32'sd147731, -32'sd1829109, 32'sd360500, 32'sd1295128, -32'sd279003, 32'sd85292, 32'sd1114646, 32'sd1165795, -32'sd73864, -32'sd18439, 32'sd372497, 32'sd1022636, -32'sd1615664, -32'sd857135, -32'sd892928, 32'sd69178, -32'sd198895, -32'sd594265, -32'sd735273, 32'sd206245, -32'sd2891151, -32'sd190826, -32'sd3662578, -32'sd458511, -32'sd2047612, -32'sd454690, -32'sd408440, 32'sd547809, 32'sd175821, -32'sd115762, -32'sd168501, 32'sd1141509, 32'sd1003557, 32'sd0, 32'sd302552, 32'sd1414268, -32'sd52438, -32'sd577839, 32'sd1924744, 32'sd1876070, 32'sd1275298, 32'sd1514417, -32'sd1057575, 32'sd640435, -32'sd1085007, -32'sd2142493, -32'sd23264, -32'sd1238497, -32'sd815896, -32'sd1646588, -32'sd2236083, -32'sd1146229, -32'sd2182771, -32'sd1111322, -32'sd443162, 32'sd53635, 32'sd1505327, -32'sd1352871, -32'sd2192684, -32'sd783359, -32'sd1577002, -32'sd143109, 32'sd313814, 32'sd1271216, 32'sd97096, -32'sd137252, 32'sd729294, 32'sd2106216, 32'sd774617, 32'sd1663182, -32'sd166999, 32'sd1041643, -32'sd1262845, -32'sd154202, 32'sd126540, 32'sd259497, -32'sd779812, -32'sd329803, -32'sd1736603, -32'sd1591949, -32'sd2595382, -32'sd2174566, -32'sd708459, -32'sd198210, -32'sd641169, 32'sd931720, 32'sd460780, -32'sd809442, -32'sd616591, 32'sd294700, -32'sd1354490, 32'sd178307, -32'sd498047, -32'sd18270, -32'sd383023, 32'sd2315403, 32'sd2150228, 32'sd1768650, -32'sd548234, -32'sd568293, 32'sd698721, 32'sd1380882, -32'sd367926, 32'sd1239648, 32'sd1285059, -32'sd537649, -32'sd1388868, -32'sd690041, -32'sd1414780, 32'sd191224, -32'sd1106735, -32'sd2627936, 32'sd265693, -32'sd395177, 32'sd1079484, -32'sd872976, -32'sd789397, 32'sd0, 32'sd645993, -32'sd69884, -32'sd620934, -32'sd544786, 32'sd2032088, 32'sd2631120, 32'sd151544, 32'sd747921, 32'sd2821459, 32'sd765014, -32'sd473371, 32'sd1932751, 32'sd1410184, 32'sd2878923, 32'sd2373702, 32'sd1667298, -32'sd866030, -32'sd260233, -32'sd1432546, 32'sd16193, -32'sd359913, 32'sd403217, -32'sd501771, 32'sd94363, 32'sd690225, -32'sd1612336, 32'sd1934192, -32'sd283395, -32'sd730556, -32'sd1373979, -32'sd2146238, -32'sd3053677, -32'sd524727, 32'sd1416302, -32'sd183939, 32'sd739977, 32'sd877989, 32'sd1953455, 32'sd1821062, 32'sd2597446, -32'sd102245, 32'sd2983067, 32'sd656614, 32'sd337690, 32'sd1517480, 32'sd1395894, -32'sd1285414, 32'sd117313, 32'sd97015, 32'sd493576, 32'sd317244, 32'sd225898, -32'sd680982, -32'sd729377, -32'sd121410, 32'sd1979852, 32'sd1963922, 32'sd1405156, 32'sd1487936, -32'sd2437807, -32'sd1976947, -32'sd1197527, -32'sd2159610, -32'sd191285, -32'sd780612, 32'sd2523723, 32'sd1454849, -32'sd129830, 32'sd1559284, 32'sd863224, -32'sd244095, -32'sd244126, 32'sd860668, -32'sd53679, 32'sd665783, -32'sd158692, 32'sd1813172, -32'sd2774441, 32'sd893727, -32'sd572381, 32'sd202745, -32'sd213231, 32'sd440511, 32'sd0, 32'sd194826, -32'sd666567, -32'sd731314, -32'sd1029103, -32'sd388074, -32'sd1151895, -32'sd2388304, -32'sd551919, 32'sd219806, 32'sd157134, -32'sd447885, 32'sd1756121, -32'sd319744, -32'sd995419, 32'sd255239, 32'sd949730, -32'sd297199, -32'sd1468622, -32'sd83321, 32'sd408376, -32'sd1714180, -32'sd1334906, 32'sd916389, 32'sd156293, -32'sd129829, 32'sd1812338, 32'sd0, 32'sd0, 32'sd0, 32'sd1426456, 32'sd106060, -32'sd678401, -32'sd622527, 32'sd203331, 32'sd473835, -32'sd1139045, 32'sd904030, 32'sd670485, -32'sd1802306, 32'sd419423, -32'sd1923983, -32'sd1242523, -32'sd1387422, 32'sd1130048, -32'sd1262535, -32'sd821589, -32'sd723869, -32'sd322082, 32'sd3074065, -32'sd1005007, -32'sd1857652, -32'sd28513, 32'sd585697, -32'sd600030, 32'sd0, 32'sd0, 32'sd0, 32'sd672902, -32'sd1055696, 32'sd83037, -32'sd1085394, -32'sd909858, -32'sd493378, -32'sd569749, -32'sd539465, -32'sd218521, -32'sd962830, -32'sd259556, -32'sd802084, 32'sd1493176, -32'sd633823, -32'sd167449, -32'sd1375020, 32'sd2843855, 32'sd1223351, 32'sd219115, 32'sd770010, -32'sd277896, -32'sd701844, -32'sd585429, 32'sd453080, 32'sd282730, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1210811, 32'sd395108, -32'sd580857, -32'sd749474, 32'sd22627, -32'sd1541828, -32'sd888782, -32'sd3097763, -32'sd1084718, -32'sd975345, -32'sd664741, -32'sd1898215, 32'sd1965129, 32'sd1136245, -32'sd2237102, -32'sd118871, -32'sd694699, 32'sd977875, 32'sd1113064, 32'sd417965, -32'sd721422, 32'sd137225, 32'sd665662, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1065452, 32'sd834239, 32'sd269190, -32'sd299814, 32'sd1420059, 32'sd1151411, 32'sd867586, 32'sd1316096, 32'sd966963, -32'sd1367313, -32'sd294554, 32'sd1779757, 32'sd1500995, 32'sd112017, 32'sd167394, 32'sd406232, 32'sd491553, 32'sd1481647, -32'sd773113, 32'sd853530, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd748538, -32'sd404006, -32'sd277026, 32'sd171429, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd727535, 32'sd106062, -32'sd992676, 32'sd208576, 32'sd518625, -32'sd1179719, 32'sd10234, -32'sd1428149, -32'sd1068788, -32'sd366880, -32'sd712988, -32'sd310241, -32'sd1464523, 32'sd77141, 32'sd913202, -32'sd2090495, -32'sd938294, -32'sd1425924, -32'sd1198036, -32'sd483875, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd606625, -32'sd174815, 32'sd85302, 32'sd199073, -32'sd980780, -32'sd1630985, -32'sd1741970, 32'sd756359, -32'sd1169612, -32'sd2536528, -32'sd828399, -32'sd2802112, -32'sd2423431, -32'sd600952, -32'sd2534283, 32'sd620821, 32'sd2761791, -32'sd1987090, 32'sd586222, -32'sd249707, 32'sd1903886, -32'sd1791387, -32'sd834660, -32'sd1139219, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1047766, -32'sd1303022, 32'sd425893, -32'sd614, -32'sd1529073, -32'sd1708208, -32'sd1696693, -32'sd456876, -32'sd1298608, 32'sd935977, -32'sd2180139, -32'sd2928732, -32'sd1303262, -32'sd1162751, -32'sd2439873, 32'sd132779, 32'sd1580736, -32'sd1049177, 32'sd1016882, 32'sd1688754, 32'sd1712890, 32'sd268451, 32'sd1589717, -32'sd1791248, -32'sd3407, 32'sd0, 32'sd0, 32'sd246250, 32'sd659136, -32'sd1154210, -32'sd835889, -32'sd208116, 32'sd29777, 32'sd472080, -32'sd401826, -32'sd4370857, -32'sd3304393, -32'sd2308214, -32'sd1489103, -32'sd1741601, -32'sd2373810, 32'sd285757, 32'sd381315, 32'sd1521074, 32'sd478031, -32'sd2525890, -32'sd1589703, -32'sd26086, 32'sd594849, 32'sd1360514, 32'sd64101, -32'sd1221109, -32'sd1280184, -32'sd194458, 32'sd0, -32'sd321741, -32'sd705340, -32'sd985489, 32'sd788081, -32'sd569968, -32'sd837396, -32'sd1017436, -32'sd757461, -32'sd1585557, -32'sd1756210, -32'sd27464, 32'sd1211370, 32'sd879682, 32'sd452775, -32'sd443881, -32'sd508174, -32'sd196844, -32'sd243799, 32'sd1185251, 32'sd958263, -32'sd1940950, -32'sd1846370, -32'sd1477734, -32'sd1034235, 32'sd371504, 32'sd911025, -32'sd585359, 32'sd0, 32'sd828315, 32'sd686556, -32'sd659537, -32'sd1782958, -32'sd2711303, 32'sd280255, -32'sd1381055, -32'sd533600, 32'sd652507, 32'sd1182127, 32'sd472714, 32'sd1193075, 32'sd121754, 32'sd1510607, 32'sd481258, 32'sd509564, 32'sd788604, -32'sd406851, 32'sd1696492, 32'sd3582507, 32'sd1209711, 32'sd397750, -32'sd1254538, -32'sd166002, 32'sd544332, 32'sd1171686, -32'sd1101682, -32'sd124942, -32'sd1453154, 32'sd332467, 32'sd159700, -32'sd1050402, 32'sd122549, 32'sd272104, -32'sd1258450, -32'sd24913, -32'sd1058151, 32'sd473906, 32'sd79639, 32'sd1113955, 32'sd745308, -32'sd344797, 32'sd121055, -32'sd108751, 32'sd1787487, 32'sd2669174, 32'sd2247271, 32'sd2529894, 32'sd1927431, 32'sd1944547, 32'sd368444, 32'sd766098, 32'sd960447, 32'sd372137, 32'sd451965, -32'sd387268, 32'sd95153, -32'sd1506457, -32'sd920859, -32'sd200807, 32'sd54407, 32'sd372950, -32'sd560268, -32'sd1542039, -32'sd1597343, -32'sd2277016, -32'sd2541015, -32'sd2143426, -32'sd1130084, -32'sd660531, 32'sd115148, 32'sd848793, 32'sd2830403, 32'sd3545494, 32'sd539796, 32'sd1718371, 32'sd1341812, 32'sd836789, 32'sd1226142, 32'sd2522276, 32'sd1443787, -32'sd523042, -32'sd231379, -32'sd872276, 32'sd212237, 32'sd1392105, -32'sd1155374, -32'sd2389289, -32'sd47419, -32'sd779310, -32'sd1192254, 32'sd347337, -32'sd564802, 32'sd118177, 32'sd648876, -32'sd484903, 32'sd4886, -32'sd701429, 32'sd884345, 32'sd2121070, 32'sd1249806, 32'sd1783037, 32'sd1400987, 32'sd1659717, 32'sd1480578, 32'sd532762, 32'sd902783, -32'sd144351, 32'sd938101, -32'sd9746, 32'sd373644, -32'sd163874, 32'sd180284, -32'sd1039872, 32'sd110130, 32'sd540373, 32'sd1678689, 32'sd151490, 32'sd1668559, -32'sd1829264, 32'sd1046787, 32'sd1084980, -32'sd326203, -32'sd878878, -32'sd1647506, -32'sd932370, -32'sd11640, -32'sd1517435, -32'sd3590370, -32'sd1689391, -32'sd303892, -32'sd653537, 32'sd470355, 32'sd240459, 32'sd1006955, 32'sd1177640, 32'sd1443539, -32'sd555496, -32'sd1008894, 32'sd641288, -32'sd71396, -32'sd1942457, 32'sd54535, 32'sd1924454, 32'sd1939283, 32'sd152405, -32'sd489466, 32'sd845866, 32'sd2573864, -32'sd600370, -32'sd2344192, -32'sd2282958, -32'sd2454915, -32'sd2868564, -32'sd477658, -32'sd4138330, -32'sd3960263, -32'sd2499519, -32'sd1476282, -32'sd960347, 32'sd175239, 32'sd1951906, 32'sd453517, -32'sd2391822, 32'sd1054139, 32'sd534669, -32'sd1104945, -32'sd795622, -32'sd481499, 32'sd744910, 32'sd1483347, 32'sd1907955, 32'sd98104, 32'sd2606689, 32'sd2463707, 32'sd2638141, 32'sd784432, -32'sd1186578, -32'sd3389283, -32'sd475442, -32'sd2063513, -32'sd4017266, -32'sd477163, -32'sd2564225, -32'sd3654832, -32'sd1119689, -32'sd723369, 32'sd828341, 32'sd1345818, 32'sd1851525, 32'sd137854, -32'sd1598807, 32'sd109414, -32'sd3002564, 32'sd326709, 32'sd543231, -32'sd227168, 32'sd394586, 32'sd1138940, 32'sd1457820, 32'sd699795, 32'sd303508, 32'sd3140169, 32'sd3202979, 32'sd1440149, 32'sd1415448, -32'sd1184623, -32'sd1042352, -32'sd63659, -32'sd145808, -32'sd1865929, -32'sd2697803, -32'sd2602334, -32'sd2689082, -32'sd593210, 32'sd1374137, 32'sd1390793, -32'sd836276, -32'sd1390935, 32'sd441806, 32'sd1265988, 32'sd452833, -32'sd242401, -32'sd475540, -32'sd248341, -32'sd635066, 32'sd1455529, -32'sd58623, 32'sd1239265, 32'sd1143518, 32'sd1705828, 32'sd536764, 32'sd1021345, 32'sd3771304, 32'sd1285576, -32'sd1575177, 32'sd1642994, 32'sd2104977, 32'sd1689918, -32'sd459573, -32'sd282344, -32'sd1840407, 32'sd41738, 32'sd863698, 32'sd122537, -32'sd312971, -32'sd2443766, 32'sd597953, 32'sd514510, -32'sd1165971, -32'sd510409, 32'sd954704, -32'sd1338562, 32'sd47559, 32'sd1814911, 32'sd1384330, 32'sd668903, 32'sd2365499, -32'sd781143, 32'sd1084247, 32'sd1372750, 32'sd2382925, -32'sd153312, 32'sd1833516, 32'sd905458, 32'sd326484, 32'sd1139901, 32'sd280625, -32'sd442423, 32'sd1054845, -32'sd1291515, 32'sd378241, -32'sd1605957, -32'sd1018821, 32'sd31282, -32'sd1065102, -32'sd1668443, -32'sd206263, -32'sd355089, 32'sd121542, -32'sd1919524, 32'sd138737, -32'sd512667, -32'sd866952, 32'sd1374508, -32'sd932304, -32'sd475500, -32'sd947550, 32'sd2534535, 32'sd2251246, 32'sd2275823, 32'sd1943116, 32'sd2299969, 32'sd713047, 32'sd1388224, 32'sd1877756, 32'sd582938, -32'sd346607, 32'sd116024, 32'sd466405, -32'sd2168774, -32'sd1708521, -32'sd958951, -32'sd2859291, -32'sd1952760, 32'sd1610864, -32'sd542513, 32'sd0, 32'sd526772, 32'sd75811, 32'sd1552630, -32'sd1305795, -32'sd825438, -32'sd76566, -32'sd1685751, 32'sd11054, 32'sd718804, 32'sd2898449, 32'sd3881614, 32'sd4612350, 32'sd3384600, 32'sd2430875, 32'sd3148943, 32'sd1417046, 32'sd2408287, 32'sd1865660, 32'sd423738, -32'sd587502, 32'sd106300, -32'sd1025089, -32'sd3246887, -32'sd3074511, -32'sd415318, -32'sd161073, -32'sd2007126, -32'sd288315, 32'sd416741, 32'sd1416185, 32'sd1401509, -32'sd956094, -32'sd1397528, -32'sd1253769, -32'sd717550, -32'sd2753669, -32'sd2154633, 32'sd907317, 32'sd3037211, 32'sd1157266, 32'sd1992881, 32'sd1257340, 32'sd1273214, 32'sd3070710, 32'sd1975155, 32'sd261729, 32'sd1997145, 32'sd225022, -32'sd412980, -32'sd795044, -32'sd2952442, -32'sd1261132, 32'sd1761435, 32'sd605333, -32'sd309305, -32'sd760299, -32'sd233623, 32'sd821323, 32'sd828697, 32'sd794518, -32'sd2360579, -32'sd2910396, -32'sd3110094, -32'sd3093161, -32'sd4435684, -32'sd508967, -32'sd600866, -32'sd1384158, 32'sd297599, 32'sd357268, 32'sd210886, 32'sd3048918, 32'sd1674082, 32'sd2259891, 32'sd352377, -32'sd30038, -32'sd659665, -32'sd1131175, 32'sd89377, -32'sd427438, -32'sd614286, 32'sd445544, -32'sd1083684, 32'sd0, -32'sd387345, -32'sd408007, -32'sd1137904, 32'sd807974, 32'sd998552, 32'sd191721, -32'sd2982716, -32'sd3018714, -32'sd3262408, -32'sd3087578, -32'sd2074435, -32'sd3040721, -32'sd1373118, -32'sd834857, 32'sd1531905, 32'sd2837649, 32'sd2828729, 32'sd1937992, -32'sd255766, 32'sd172324, 32'sd751048, 32'sd1550283, 32'sd890707, 32'sd718299, 32'sd1593393, -32'sd1027067, 32'sd897013, 32'sd350609, -32'sd219852, 32'sd1305523, -32'sd256451, 32'sd404953, 32'sd912553, -32'sd562782, -32'sd226198, -32'sd69308, -32'sd1946891, -32'sd2565478, -32'sd2386976, -32'sd3960435, -32'sd2619285, 32'sd652604, 32'sd1615580, 32'sd3913276, 32'sd1982204, 32'sd1297740, -32'sd718544, 32'sd171107, 32'sd1131821, 32'sd172497, 32'sd807953, 32'sd1885158, 32'sd460774, -32'sd982594, -32'sd420527, -32'sd654463, 32'sd732797, 32'sd888477, -32'sd1258536, 32'sd336109, 32'sd138245, -32'sd390883, -32'sd1090290, -32'sd971874, 32'sd1770398, 32'sd765890, -32'sd784858, -32'sd596892, -32'sd116259, 32'sd1497075, 32'sd2329612, 32'sd290618, 32'sd157007, -32'sd690946, -32'sd1836592, 32'sd1706455, 32'sd1548254, 32'sd629340, 32'sd464032, 32'sd1116814, -32'sd3192089, -32'sd643365, -32'sd269778, 32'sd0, -32'sd569733, -32'sd906577, 32'sd795222, 32'sd1188483, 32'sd1080317, -32'sd841393, 32'sd516462, 32'sd1322114, -32'sd462903, 32'sd1225588, 32'sd627154, 32'sd985677, 32'sd3002933, -32'sd345756, 32'sd597912, 32'sd339098, -32'sd2757704, -32'sd1985936, -32'sd506197, -32'sd337073, 32'sd2664196, 32'sd1821293, 32'sd1173866, -32'sd1229824, -32'sd1682261, -32'sd594585, 32'sd0, 32'sd0, 32'sd0, -32'sd611529, -32'sd18743, 32'sd1449931, 32'sd279774, -32'sd137087, 32'sd1203423, 32'sd657976, 32'sd224851, 32'sd1584023, 32'sd1400612, 32'sd1567599, 32'sd2364123, 32'sd2423272, 32'sd2571182, -32'sd795427, -32'sd382173, 32'sd138589, 32'sd341620, 32'sd1897685, 32'sd1992836, 32'sd1860947, -32'sd524719, -32'sd1097705, -32'sd1633554, -32'sd552540, 32'sd0, 32'sd0, 32'sd0, -32'sd1222548, -32'sd1457117, 32'sd1060539, -32'sd416528, 32'sd1587295, -32'sd469902, 32'sd764270, -32'sd73592, 32'sd1086203, 32'sd2314520, 32'sd291096, 32'sd936027, -32'sd2016321, 32'sd881441, 32'sd144153, 32'sd505917, -32'sd464708, 32'sd639793, 32'sd785849, -32'sd528665, 32'sd150446, -32'sd200042, -32'sd72830, 32'sd615985, 32'sd666487, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd690242, -32'sd469449, -32'sd554783, 32'sd481985, 32'sd1958377, 32'sd112658, 32'sd551999, 32'sd1324522, 32'sd1858574, 32'sd1740214, 32'sd3018791, -32'sd276627, 32'sd20480, 32'sd209535, -32'sd728707, -32'sd1654804, -32'sd2689546, -32'sd367225, 32'sd1521334, -32'sd1018203, 32'sd1247414, 32'sd1412905, 32'sd726870, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd294913, 32'sd870904, -32'sd400054, -32'sd780587, 32'sd190955, 32'sd355753, 32'sd479403, 32'sd922714, 32'sd1227554, 32'sd1141463, 32'sd1137065, -32'sd365639, -32'sd2063679, -32'sd1701996, 32'sd60979, -32'sd1810267, -32'sd728450, -32'sd1422608, 32'sd374495, -32'sd779759, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd782471, 32'sd1102381, 32'sd714255, -32'sd1280640, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd941354, 32'sd647584, -32'sd1810542, -32'sd390648, -32'sd294553, 32'sd221084, -32'sd621014, 32'sd1386204, -32'sd145805, 32'sd2017958, -32'sd839987, 32'sd733245, -32'sd1175535, 32'sd378275, 32'sd1634568, 32'sd2027237, 32'sd794624, 32'sd301798, 32'sd1447045, 32'sd1659432, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1684839, 32'sd602908, 32'sd1425683, 32'sd389438, -32'sd332250, -32'sd1307952, -32'sd40021, -32'sd1583693, -32'sd690296, -32'sd1031695, -32'sd935395, -32'sd677695, -32'sd1783371, -32'sd218687, -32'sd265038, -32'sd127686, -32'sd134251, -32'sd765438, -32'sd461972, 32'sd1655441, 32'sd2153355, -32'sd525063, 32'sd683060, 32'sd2553436, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1191731, 32'sd2141310, 32'sd999635, -32'sd786501, -32'sd2197709, 32'sd184576, -32'sd362377, -32'sd982024, 32'sd1134469, -32'sd1390805, -32'sd113340, 32'sd414531, -32'sd1173217, -32'sd767822, -32'sd368517, 32'sd2686196, 32'sd1141899, 32'sd1324569, 32'sd239286, 32'sd1607291, 32'sd955210, 32'sd251535, 32'sd610285, 32'sd660152, 32'sd1613793, 32'sd0, 32'sd0, 32'sd1008634, -32'sd35784, 32'sd1223706, 32'sd575406, 32'sd253631, -32'sd2078827, -32'sd979394, 32'sd382684, -32'sd592554, -32'sd2694264, -32'sd1374223, -32'sd1262594, -32'sd747663, -32'sd950087, -32'sd165925, -32'sd634408, 32'sd438422, -32'sd264103, 32'sd381417, -32'sd1195684, 32'sd122111, 32'sd467932, 32'sd1393255, -32'sd1404198, 32'sd843508, 32'sd399507, -32'sd422669, 32'sd0, 32'sd653083, 32'sd24168, -32'sd1091990, 32'sd1701770, 32'sd2093219, 32'sd1681709, 32'sd691926, -32'sd418175, -32'sd2156825, -32'sd2634275, -32'sd2092933, -32'sd385619, -32'sd1357085, -32'sd437805, -32'sd490709, -32'sd1236599, -32'sd624553, -32'sd573709, -32'sd1646513, -32'sd117346, -32'sd251758, 32'sd640065, 32'sd221704, 32'sd442295, 32'sd1132901, -32'sd63049, 32'sd1173152, 32'sd0, -32'sd192988, 32'sd436501, -32'sd1467855, 32'sd1367744, 32'sd269011, 32'sd827369, 32'sd1599587, -32'sd319733, -32'sd1368137, -32'sd3228760, -32'sd1970580, -32'sd265399, 32'sd1488283, 32'sd483519, -32'sd142851, 32'sd450249, 32'sd2087392, 32'sd394543, 32'sd1046527, 32'sd1754002, 32'sd182632, 32'sd35764, 32'sd113158, 32'sd1455953, 32'sd356405, -32'sd111727, 32'sd44831, 32'sd1981215, 32'sd1211607, -32'sd350215, 32'sd561568, 32'sd1320222, 32'sd100807, -32'sd946738, -32'sd507584, -32'sd2015322, -32'sd399869, 32'sd318636, -32'sd1647455, 32'sd320743, -32'sd321304, 32'sd2546209, 32'sd2504816, 32'sd2087815, 32'sd2057850, -32'sd1132388, -32'sd1754779, -32'sd228977, 32'sd99552, -32'sd87348, 32'sd1817376, 32'sd212478, 32'sd1180342, 32'sd1044020, -32'sd273470, 32'sd333475, 32'sd29294, -32'sd128374, 32'sd1323942, 32'sd1034178, -32'sd137671, 32'sd1285694, 32'sd1154654, 32'sd1507356, -32'sd620596, -32'sd867201, -32'sd1315849, -32'sd999581, 32'sd1635685, 32'sd3579050, 32'sd2403084, -32'sd246443, 32'sd708538, 32'sd725659, 32'sd38154, -32'sd799458, -32'sd278921, 32'sd387488, -32'sd593426, 32'sd1583955, 32'sd541758, -32'sd472753, 32'sd510854, 32'sd1951604, 32'sd1513185, 32'sd953479, -32'sd483617, -32'sd76104, -32'sd35288, 32'sd506008, 32'sd1380049, 32'sd1492493, 32'sd99486, -32'sd3115487, -32'sd4060791, -32'sd3646458, 32'sd620785, 32'sd3632581, 32'sd1054013, -32'sd1425156, -32'sd1033589, 32'sd883446, -32'sd529970, -32'sd1592039, -32'sd421771, -32'sd1632946, 32'sd8307, 32'sd1502657, 32'sd1687603, -32'sd1011949, 32'sd1125077, 32'sd1400290, -32'sd494791, 32'sd906518, 32'sd116309, -32'sd1272606, -32'sd2683979, -32'sd1457213, 32'sd58662, 32'sd1532331, 32'sd58344, -32'sd2959212, -32'sd3998159, -32'sd1770107, 32'sd2525205, 32'sd1542656, 32'sd1529395, -32'sd460851, -32'sd1173749, 32'sd2131008, 32'sd1342215, -32'sd681504, 32'sd514092, 32'sd2048838, 32'sd79297, 32'sd930190, 32'sd1139299, -32'sd140021, 32'sd454976, 32'sd1184746, -32'sd75689, 32'sd1405786, 32'sd390927, 32'sd1154550, -32'sd2709518, -32'sd30433, 32'sd729002, 32'sd632037, -32'sd939015, -32'sd660909, -32'sd2696130, -32'sd1849312, 32'sd3656196, 32'sd2777307, -32'sd96666, -32'sd232536, 32'sd1271025, 32'sd299807, 32'sd156092, -32'sd1293471, 32'sd96324, 32'sd162018, 32'sd1287135, 32'sd1533190, -32'sd31703, 32'sd782514, 32'sd74488, 32'sd2109522, -32'sd819736, -32'sd839485, 32'sd7360, -32'sd1134059, -32'sd1088691, -32'sd11665, -32'sd207686, 32'sd1262928, 32'sd527441, -32'sd1422881, -32'sd1591458, -32'sd1249099, 32'sd3131834, 32'sd2188387, 32'sd128010, -32'sd385100, -32'sd656589, 32'sd725150, -32'sd348675, 32'sd42728, -32'sd1764297, 32'sd273244, -32'sd1307274, -32'sd2065619, 32'sd454421, 32'sd453402, 32'sd1599974, 32'sd1252375, -32'sd1515996, -32'sd62872, -32'sd1373494, 32'sd968861, 32'sd241002, 32'sd1208763, 32'sd194253, -32'sd1480993, 32'sd1427103, 32'sd1239445, -32'sd741286, 32'sd333379, -32'sd462437, 32'sd2399744, 32'sd1500363, -32'sd298598, -32'sd720150, -32'sd2632561, -32'sd578896, -32'sd354180, -32'sd646004, -32'sd1388792, -32'sd2173265, -32'sd2129104, 32'sd493107, -32'sd331038, -32'sd619646, 32'sd2788396, 32'sd349973, 32'sd1118268, 32'sd1109440, 32'sd126822, -32'sd766908, 32'sd380001, 32'sd457588, 32'sd1457465, 32'sd546953, 32'sd319852, 32'sd781807, 32'sd56090, 32'sd304288, 32'sd1514842, 32'sd988493, -32'sd1289218, -32'sd674973, -32'sd947546, -32'sd695727, 32'sd1451144, 32'sd1436227, -32'sd1369100, -32'sd4116828, -32'sd3678453, 32'sd59490, 32'sd222507, 32'sd127685, 32'sd1309552, 32'sd416568, 32'sd1420518, -32'sd80582, -32'sd1027471, 32'sd895503, 32'sd1102632, 32'sd2620881, 32'sd1783795, 32'sd1667951, -32'sd129786, 32'sd62102, -32'sd1094142, -32'sd449940, 32'sd2318900, 32'sd2245678, -32'sd1205881, 32'sd395126, -32'sd377311, 32'sd527964, 32'sd2667818, 32'sd583287, -32'sd1516186, -32'sd1600558, -32'sd1557181, 32'sd993802, -32'sd544815, -32'sd230587, 32'sd1153533, -32'sd906815, 32'sd441332, -32'sd1330370, 32'sd594929, 32'sd1565432, -32'sd1149501, -32'sd426519, 32'sd1299272, 32'sd128533, -32'sd520830, -32'sd1356770, -32'sd1068597, 32'sd1716974, 32'sd2929316, -32'sd56357, 32'sd475931, -32'sd1173077, -32'sd131560, 32'sd771749, 32'sd994903, -32'sd879873, -32'sd2172793, -32'sd464322, -32'sd1660530, -32'sd882896, -32'sd119211, -32'sd807114, 32'sd0, 32'sd92972, 32'sd1164002, 32'sd37575, 32'sd65912, -32'sd165837, -32'sd2016552, -32'sd569363, -32'sd576540, 32'sd1571638, -32'sd1097174, -32'sd1011178, -32'sd1191850, 32'sd1432494, 32'sd758043, 32'sd1761538, 32'sd1243500, -32'sd162964, -32'sd997730, -32'sd901813, 32'sd558821, -32'sd3120251, -32'sd1243940, -32'sd447535, -32'sd978134, 32'sd387985, 32'sd207011, 32'sd595881, -32'sd549640, 32'sd487921, 32'sd1643915, 32'sd347940, -32'sd2019253, -32'sd1328297, -32'sd389366, -32'sd284610, 32'sd1323982, -32'sd962428, 32'sd100366, -32'sd877659, 32'sd1626289, 32'sd3029089, 32'sd1412931, 32'sd1646436, -32'sd1739885, -32'sd1620262, -32'sd2205005, -32'sd1635344, -32'sd3025846, -32'sd2116508, -32'sd2569064, -32'sd290641, -32'sd912361, 32'sd1231787, 32'sd123204, 32'sd716299, 32'sd1148607, -32'sd120525, -32'sd971776, -32'sd807843, -32'sd165068, -32'sd522113, -32'sd27813, 32'sd257523, 32'sd497244, 32'sd1530373, 32'sd101699, -32'sd758697, 32'sd3103267, 32'sd3221589, 32'sd2005091, -32'sd57687, -32'sd1429099, -32'sd3220737, -32'sd3392282, -32'sd1937878, -32'sd2132381, -32'sd4488427, -32'sd3323458, -32'sd2776133, 32'sd560420, 32'sd768060, 32'sd1050385, 32'sd615115, 32'sd0, -32'sd136775, -32'sd1999657, -32'sd1848809, -32'sd1557583, 32'sd1132984, -32'sd364091, -32'sd1425537, -32'sd345304, -32'sd1202380, 32'sd754288, 32'sd548398, 32'sd1125895, 32'sd2496434, 32'sd889196, -32'sd2106436, -32'sd2878454, -32'sd2101956, -32'sd1312656, 32'sd123110, -32'sd2644575, -32'sd2333935, -32'sd2722372, -32'sd1902752, -32'sd53796, -32'sd524023, 32'sd846496, 32'sd1029113, 32'sd360272, 32'sd607792, -32'sd1713053, -32'sd617434, -32'sd882563, 32'sd432207, -32'sd308815, 32'sd1238796, 32'sd1021223, 32'sd718022, 32'sd833522, 32'sd1603844, 32'sd2064662, 32'sd887616, 32'sd1627202, -32'sd2050697, -32'sd1544364, -32'sd812717, -32'sd2070284, -32'sd1745123, -32'sd418240, -32'sd553151, -32'sd1497243, 32'sd296100, 32'sd1252084, -32'sd801016, -32'sd522884, 32'sd818584, 32'sd1917330, 32'sd1614957, -32'sd1582569, -32'sd64666, -32'sd1593887, 32'sd58667, 32'sd409095, -32'sd68676, 32'sd1057693, 32'sd1677273, 32'sd1534652, 32'sd830688, 32'sd966463, 32'sd2587998, -32'sd16812, -32'sd1038732, -32'sd3092921, -32'sd1693309, -32'sd814446, -32'sd1188752, -32'sd820034, 32'sd521945, 32'sd946829, 32'sd176266, -32'sd121444, 32'sd4173, 32'sd314906, 32'sd1247247, 32'sd0, 32'sd1445514, -32'sd540431, -32'sd2253340, -32'sd338423, -32'sd251416, -32'sd220046, -32'sd786534, -32'sd1166758, -32'sd331301, 32'sd180050, 32'sd134579, 32'sd999075, -32'sd1095268, -32'sd1854728, -32'sd2079130, -32'sd2375512, -32'sd2246616, -32'sd2074706, -32'sd1983138, 32'sd712284, -32'sd1805318, -32'sd645472, -32'sd897428, 32'sd406109, 32'sd1238243, 32'sd30095, 32'sd0, 32'sd0, 32'sd0, -32'sd669814, 32'sd523745, -32'sd143056, 32'sd702646, 32'sd998610, -32'sd101573, -32'sd202773, 32'sd432663, -32'sd325772, 32'sd787376, 32'sd470661, -32'sd2934415, -32'sd1026934, 32'sd156027, -32'sd1190142, -32'sd1412887, -32'sd2710763, -32'sd2796116, -32'sd650642, -32'sd544579, -32'sd373509, -32'sd225525, -32'sd401232, -32'sd1121430, 32'sd543808, 32'sd0, 32'sd0, 32'sd0, -32'sd381860, 32'sd657473, -32'sd769828, 32'sd802885, -32'sd813701, 32'sd957170, 32'sd814721, 32'sd1460569, 32'sd859548, 32'sd18282, -32'sd835489, -32'sd1610663, 32'sd784127, 32'sd2264666, -32'sd165124, -32'sd428297, -32'sd1938222, -32'sd1968346, -32'sd102803, -32'sd649106, 32'sd685069, 32'sd954544, -32'sd895717, -32'sd386510, 32'sd223480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2174367, -32'sd1749948, -32'sd1123600, -32'sd152838, 32'sd1152897, 32'sd30898, -32'sd87006, 32'sd361751, 32'sd1529519, -32'sd236208, 32'sd1261089, -32'sd479626, -32'sd134158, -32'sd304778, 32'sd1997760, 32'sd1119233, -32'sd567129, 32'sd1204628, -32'sd754742, 32'sd1085328, -32'sd14120, 32'sd1839530, 32'sd1341989, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1036960, -32'sd805955, 32'sd1261710, 32'sd332177, -32'sd1302258, 32'sd123737, 32'sd1013750, -32'sd169949, 32'sd1605609, 32'sd1531839, 32'sd963394, 32'sd75752, 32'sd1510344, 32'sd196807, -32'sd641066, 32'sd293485, 32'sd1424970, -32'sd416938, -32'sd49529, 32'sd1804618, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1217925, 32'sd393794, 32'sd890587, 32'sd1736743, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd477530, -32'sd45496, -32'sd404566, -32'sd293464, 32'sd1257239, -32'sd1364494, 32'sd557623, -32'sd1468450, 32'sd702531, -32'sd1317141, 32'sd1852391, 32'sd582740, -32'sd83132, 32'sd1361015, -32'sd1007963, -32'sd178897, -32'sd1985, 32'sd47000, 32'sd209113, 32'sd1050136, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd743481, -32'sd916617, 32'sd375219, -32'sd424114, -32'sd871378, -32'sd1010154, -32'sd1235731, -32'sd574492, 32'sd1742430, 32'sd761640, 32'sd23681, 32'sd548392, 32'sd877578, -32'sd1379975, 32'sd556395, 32'sd376838, -32'sd394986, 32'sd2493726, 32'sd1553398, -32'sd457787, 32'sd1455629, -32'sd1103887, 32'sd1215173, 32'sd1507650, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1151367, 32'sd985681, -32'sd717131, 32'sd322675, 32'sd751695, -32'sd832765, 32'sd1649233, 32'sd946747, -32'sd1505689, 32'sd1083796, -32'sd2358156, -32'sd2784387, -32'sd277158, -32'sd782825, -32'sd54481, 32'sd1675492, 32'sd822000, 32'sd729994, 32'sd1600915, 32'sd509938, 32'sd472824, -32'sd471969, -32'sd1366660, -32'sd883148, 32'sd634957, 32'sd0, 32'sd0, 32'sd1689358, -32'sd120333, 32'sd635131, 32'sd789603, 32'sd54940, 32'sd64329, 32'sd57962, -32'sd1014802, -32'sd1019739, -32'sd289820, -32'sd356835, -32'sd1224429, -32'sd538949, -32'sd160761, 32'sd892139, 32'sd1299410, 32'sd688419, 32'sd1047322, 32'sd1120050, 32'sd973526, 32'sd1712603, 32'sd1023027, -32'sd375733, -32'sd662162, -32'sd101752, -32'sd1006538, 32'sd1348861, 32'sd0, 32'sd1721350, -32'sd1028671, 32'sd1455541, 32'sd558171, -32'sd945129, 32'sd351040, -32'sd134420, 32'sd137490, 32'sd794332, 32'sd921865, 32'sd39050, 32'sd2106399, 32'sd900275, -32'sd1365766, -32'sd1187264, 32'sd1420898, 32'sd2453586, 32'sd668581, -32'sd422738, 32'sd64483, 32'sd202994, -32'sd2084224, -32'sd866851, -32'sd357112, -32'sd130387, 32'sd244531, -32'sd1352163, 32'sd0, 32'sd757748, 32'sd1475482, -32'sd1025038, 32'sd672544, 32'sd810418, 32'sd893881, 32'sd1470800, 32'sd93170, 32'sd59325, -32'sd1131309, -32'sd1366182, 32'sd1387300, -32'sd1734211, -32'sd718406, -32'sd1730511, 32'sd1704207, 32'sd2071448, 32'sd1837324, 32'sd2475555, -32'sd284866, -32'sd1337812, -32'sd1105767, 32'sd340979, -32'sd997041, 32'sd151772, -32'sd455589, 32'sd616466, 32'sd855924, 32'sd617520, -32'sd909054, -32'sd591370, 32'sd1349428, 32'sd770818, 32'sd2190788, 32'sd3592517, 32'sd1626018, 32'sd90222, 32'sd445975, -32'sd1782144, -32'sd1748161, -32'sd2562590, -32'sd4473613, -32'sd1809360, -32'sd171112, 32'sd2925609, 32'sd3105180, 32'sd1433749, -32'sd1899193, -32'sd1665104, -32'sd1135551, -32'sd2495958, -32'sd568736, 32'sd1920431, -32'sd641651, 32'sd524815, 32'sd69402, 32'sd877370, 32'sd867330, 32'sd1171494, -32'sd456007, 32'sd556105, 32'sd70753, 32'sd2267487, 32'sd851025, 32'sd2281263, 32'sd215687, -32'sd1608195, -32'sd628010, -32'sd2242583, -32'sd4454222, -32'sd1847481, 32'sd2048061, 32'sd3581771, 32'sd1259465, -32'sd1575508, -32'sd3506089, -32'sd4662108, -32'sd2062860, -32'sd300367, 32'sd1259270, 32'sd2076029, 32'sd1611372, 32'sd229705, -32'sd334345, 32'sd995351, 32'sd227419, -32'sd440843, 32'sd912190, 32'sd1478837, 32'sd1070017, 32'sd1316349, 32'sd1432767, -32'sd613572, -32'sd417552, 32'sd1046540, 32'sd833240, -32'sd1544478, -32'sd336597, 32'sd2251992, 32'sd5454302, 32'sd4258820, 32'sd1174803, -32'sd3580045, -32'sd3952625, -32'sd3263974, 32'sd156785, 32'sd1011229, -32'sd54514, 32'sd1028423, -32'sd1012219, 32'sd58794, 32'sd1570965, 32'sd1028302, -32'sd365730, -32'sd442472, 32'sd1247601, -32'sd1590513, 32'sd906394, 32'sd1450455, 32'sd1596601, -32'sd74404, -32'sd656169, 32'sd1372812, 32'sd421046, 32'sd212248, 32'sd946386, 32'sd2387961, 32'sd4224654, 32'sd1679930, -32'sd2584364, -32'sd4324475, -32'sd2227215, -32'sd2019617, 32'sd367514, 32'sd2663859, -32'sd2343536, 32'sd1136275, 32'sd1052052, 32'sd328639, 32'sd1895335, 32'sd155311, -32'sd1167012, 32'sd202500, 32'sd1369886, 32'sd1117909, -32'sd627150, -32'sd677453, 32'sd2016197, 32'sd1273591, 32'sd942943, 32'sd1807157, 32'sd1474429, 32'sd1153932, 32'sd2707802, 32'sd3570729, 32'sd1768504, -32'sd2286431, -32'sd4174500, -32'sd3007853, -32'sd1186661, -32'sd273985, -32'sd24120, 32'sd425769, -32'sd2758152, 32'sd107496, -32'sd1170161, -32'sd398642, 32'sd580000, 32'sd340091, 32'sd1501490, -32'sd430163, 32'sd359457, 32'sd1217233, 32'sd1125951, 32'sd634963, 32'sd934155, 32'sd1096416, 32'sd5101923, 32'sd2706709, 32'sd1590406, 32'sd355912, 32'sd606370, 32'sd1743758, 32'sd1231103, -32'sd1907927, -32'sd2432504, -32'sd534008, 32'sd33879, 32'sd343671, -32'sd44039, 32'sd803166, -32'sd298494, 32'sd245309, -32'sd1774080, -32'sd160550, 32'sd881615, -32'sd373559, 32'sd1715384, -32'sd1300096, -32'sd1731259, 32'sd212286, -32'sd505214, 32'sd311093, 32'sd1316525, 32'sd2037505, 32'sd487421, 32'sd1456345, 32'sd200519, 32'sd497428, 32'sd545797, 32'sd1080067, 32'sd145744, -32'sd783969, 32'sd1487100, -32'sd633332, 32'sd1958163, 32'sd555208, -32'sd1027156, 32'sd370500, 32'sd1309192, 32'sd2399024, 32'sd714159, -32'sd354141, -32'sd164086, 32'sd836746, 32'sd359634, -32'sd129442, -32'sd464012, 32'sd382983, -32'sd457022, -32'sd1575519, 32'sd69724, -32'sd1009170, -32'sd1263408, 32'sd382604, 32'sd212886, 32'sd2851919, 32'sd1927258, 32'sd1779127, -32'sd720451, -32'sd2519297, -32'sd13140, 32'sd1950630, -32'sd1001699, 32'sd463689, 32'sd1196704, -32'sd247033, -32'sd965449, -32'sd354819, 32'sd800637, 32'sd718221, 32'sd955727, 32'sd1335409, 32'sd520776, 32'sd501503, -32'sd1130821, -32'sd958007, 32'sd1186821, -32'sd527867, -32'sd2689227, -32'sd2382963, -32'sd1676088, 32'sd121887, -32'sd1435902, -32'sd335888, 32'sd1431000, 32'sd3758423, 32'sd619907, -32'sd817855, -32'sd289575, -32'sd1004855, 32'sd1206949, -32'sd422063, 32'sd1767073, -32'sd333093, -32'sd569413, -32'sd1774680, 32'sd768743, -32'sd80630, 32'sd1285509, 32'sd1222985, -32'sd725903, -32'sd1029172, -32'sd2113291, 32'sd542867, 32'sd2041858, 32'sd1396008, -32'sd1509539, -32'sd1230229, 32'sd1062939, 32'sd661117, 32'sd473617, -32'sd40765, -32'sd480056, 32'sd3274640, -32'sd1892497, -32'sd41185, 32'sd472876, -32'sd887042, -32'sd402171, 32'sd946821, 32'sd168269, -32'sd152709, -32'sd397143, -32'sd1762649, 32'sd26155, -32'sd693117, 32'sd0, -32'sd622650, 32'sd63541, -32'sd1567270, 32'sd998631, 32'sd1187923, -32'sd1698863, 32'sd638853, -32'sd503774, 32'sd639840, -32'sd636857, -32'sd1509480, -32'sd1094903, 32'sd1244112, 32'sd36625, 32'sd383642, -32'sd273466, 32'sd1352293, -32'sd1485710, -32'sd31201, -32'sd898947, 32'sd2019080, 32'sd1954981, 32'sd158900, 32'sd1890323, -32'sd2045857, 32'sd487007, 32'sd891655, 32'sd1212296, 32'sd1291264, -32'sd1838905, -32'sd1317812, 32'sd1032327, 32'sd396773, -32'sd235707, -32'sd1433357, 32'sd817173, -32'sd687910, -32'sd730848, -32'sd1553296, -32'sd1399110, -32'sd1553435, 32'sd130337, -32'sd1495908, -32'sd2144523, 32'sd433823, 32'sd616565, 32'sd1020890, 32'sd1911953, 32'sd1948924, 32'sd329245, 32'sd263883, 32'sd1884989, -32'sd1152964, -32'sd404757, 32'sd193675, 32'sd328868, 32'sd1131175, -32'sd973338, 32'sd2017111, 32'sd1004296, -32'sd436215, -32'sd462975, -32'sd65338, 32'sd625155, 32'sd1207923, 32'sd137994, -32'sd476357, -32'sd2349636, -32'sd2035464, -32'sd1404503, -32'sd3724430, -32'sd581015, -32'sd518737, 32'sd1234438, 32'sd361815, 32'sd672157, 32'sd1804930, -32'sd47757, -32'sd886873, 32'sd1619243, 32'sd565443, -32'sd1600396, -32'sd1033260, 32'sd0, -32'sd377580, -32'sd427787, 32'sd1647513, -32'sd882470, -32'sd1879733, 32'sd1066088, 32'sd923046, -32'sd226785, -32'sd931185, 32'sd222018, 32'sd219499, -32'sd818011, -32'sd656930, 32'sd405866, -32'sd216385, -32'sd371774, 32'sd104362, 32'sd1179976, 32'sd305105, -32'sd891947, -32'sd568974, -32'sd916249, 32'sd749599, 32'sd1161488, -32'sd387808, 32'sd468844, 32'sd502305, 32'sd1839581, 32'sd298027, 32'sd247645, -32'sd92483, -32'sd2416655, -32'sd1951434, -32'sd1627685, -32'sd431826, -32'sd1707706, -32'sd473202, -32'sd114510, 32'sd596961, -32'sd1181081, 32'sd230411, -32'sd676168, -32'sd64546, 32'sd298740, -32'sd1183666, 32'sd1230185, -32'sd1124399, 32'sd664443, -32'sd1045326, 32'sd320212, -32'sd605905, -32'sd529699, 32'sd1294301, -32'sd1301880, -32'sd541233, -32'sd104426, 32'sd2083945, -32'sd907595, -32'sd250201, 32'sd9383, -32'sd355949, -32'sd949556, -32'sd1594393, -32'sd368034, 32'sd525657, 32'sd647830, -32'sd1178261, -32'sd310974, -32'sd954642, -32'sd1280365, -32'sd73001, 32'sd401929, -32'sd54220, -32'sd602, 32'sd1809951, 32'sd1299327, -32'sd1085079, 32'sd248150, -32'sd801371, 32'sd1746550, 32'sd1066198, 32'sd213302, 32'sd679211, 32'sd0, -32'sd378929, 32'sd951461, 32'sd1140291, -32'sd237395, 32'sd54774, -32'sd699773, 32'sd1229588, 32'sd1660634, 32'sd970739, 32'sd2269299, -32'sd997685, -32'sd2405685, -32'sd211484, -32'sd1109491, 32'sd171458, -32'sd186553, -32'sd1156525, 32'sd1305400, 32'sd1286605, -32'sd979114, -32'sd467158, 32'sd962321, 32'sd1742089, -32'sd137189, -32'sd719941, -32'sd431235, 32'sd0, 32'sd0, 32'sd0, 32'sd169909, 32'sd855177, 32'sd847722, -32'sd1425856, -32'sd45581, 32'sd836283, -32'sd702941, 32'sd812938, -32'sd393692, 32'sd974128, -32'sd870658, 32'sd83668, 32'sd1591600, -32'sd1361792, -32'sd1275632, -32'sd1213415, -32'sd103636, 32'sd764902, -32'sd896547, -32'sd263152, 32'sd1159520, 32'sd56671, 32'sd407680, 32'sd198694, 32'sd248438, 32'sd0, 32'sd0, 32'sd0, 32'sd234684, -32'sd34570, -32'sd632455, -32'sd1942035, 32'sd1647751, 32'sd269595, -32'sd288153, -32'sd45089, -32'sd359096, -32'sd259001, 32'sd609417, 32'sd391079, -32'sd1264143, -32'sd110844, -32'sd175221, -32'sd408882, 32'sd1100464, -32'sd229249, -32'sd1066279, 32'sd651121, -32'sd332984, -32'sd251034, 32'sd991213, 32'sd353409, 32'sd1023809, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd295159, -32'sd517166, -32'sd43228, 32'sd837476, 32'sd920827, -32'sd611241, -32'sd2727746, 32'sd1124181, 32'sd410009, 32'sd160973, 32'sd612322, 32'sd1917455, -32'sd710685, -32'sd766121, -32'sd2954889, -32'sd1518979, 32'sd734529, -32'sd1378174, 32'sd705195, -32'sd712190, 32'sd65229, 32'sd394990, 32'sd1153489, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd672490, 32'sd1051285, 32'sd1433571, 32'sd700428, -32'sd798847, 32'sd36173, -32'sd411371, 32'sd64690, -32'sd155822, -32'sd725922, 32'sd1190692, 32'sd562860, -32'sd32211, -32'sd471737, 32'sd1018983, -32'sd708693, 32'sd55081, -32'sd263554, 32'sd930114, 32'sd1826362, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd796665, 32'sd2027974, 32'sd728759, 32'sd1024712, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1140307, 32'sd1470809, -32'sd381466, -32'sd549261, -32'sd291843, -32'sd2495728, -32'sd829758, -32'sd234466, 32'sd1439928, 32'sd2124207, -32'sd669080, 32'sd419851, -32'sd132722, 32'sd488867, 32'sd1296283, 32'sd904623, 32'sd356100, 32'sd2080194, -32'sd345826, 32'sd1212434, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1198713, 32'sd1133926, 32'sd987366, -32'sd382797, 32'sd488084, -32'sd1428436, -32'sd364374, -32'sd1591565, -32'sd2050664, 32'sd899453, 32'sd851842, 32'sd1162910, 32'sd1487580, -32'sd230466, 32'sd173834, 32'sd1466240, -32'sd320845, 32'sd199320, 32'sd1155647, 32'sd1993346, 32'sd2313788, 32'sd1301372, 32'sd1353929, 32'sd867641, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd276074, 32'sd702447, 32'sd99901, 32'sd861142, -32'sd268748, 32'sd577826, -32'sd1863203, -32'sd1942696, -32'sd42834, 32'sd991190, 32'sd238817, -32'sd20925, 32'sd1578211, 32'sd2142872, 32'sd1484670, -32'sd1564337, 32'sd398288, 32'sd634040, -32'sd9676, 32'sd657116, -32'sd784801, 32'sd506046, -32'sd2485087, 32'sd686495, 32'sd43601, 32'sd0, 32'sd0, -32'sd30461, 32'sd145150, 32'sd7107, 32'sd667649, 32'sd756569, 32'sd431332, -32'sd189373, -32'sd1052433, -32'sd629949, -32'sd1517654, 32'sd1187021, 32'sd571083, 32'sd2023600, 32'sd566833, 32'sd683723, -32'sd121819, -32'sd673076, -32'sd93325, 32'sd1198395, 32'sd1405802, 32'sd319001, -32'sd1134815, -32'sd2615556, -32'sd2383716, -32'sd1360890, -32'sd784482, 32'sd1355324, 32'sd0, -32'sd8209, 32'sd670900, 32'sd810215, -32'sd790645, 32'sd529244, -32'sd774472, -32'sd1551119, -32'sd1307737, -32'sd2437902, -32'sd3093106, -32'sd781329, -32'sd841990, 32'sd276329, 32'sd1158475, 32'sd1978059, 32'sd344878, 32'sd1826112, 32'sd1104769, 32'sd1700161, 32'sd236437, -32'sd1683894, -32'sd1009977, -32'sd2832476, -32'sd1313327, 32'sd1328521, 32'sd1518731, 32'sd597398, 32'sd0, 32'sd839849, 32'sd1281908, -32'sd664116, 32'sd1126753, -32'sd559255, 32'sd50240, -32'sd1997772, -32'sd1820139, -32'sd2192647, -32'sd2076764, -32'sd3258566, -32'sd3126356, 32'sd486035, 32'sd387695, 32'sd3703005, 32'sd2570268, -32'sd15682, -32'sd407715, -32'sd2428645, -32'sd2266981, -32'sd799861, -32'sd881327, 32'sd329312, -32'sd2567, -32'sd819094, 32'sd150518, 32'sd1504683, 32'sd722398, 32'sd321332, 32'sd202660, 32'sd2058451, 32'sd1616509, -32'sd899328, -32'sd2160326, -32'sd1420638, -32'sd2254339, -32'sd3491640, -32'sd2554703, -32'sd1942045, -32'sd1711797, -32'sd1144592, 32'sd2853271, 32'sd2011265, 32'sd130023, -32'sd1844750, -32'sd94598, -32'sd1375212, -32'sd695732, 32'sd1204028, -32'sd770905, 32'sd626643, 32'sd226971, -32'sd198568, -32'sd777688, 32'sd165687, 32'sd1078025, -32'sd469376, 32'sd1143715, -32'sd725404, -32'sd195698, 32'sd644728, -32'sd1167642, -32'sd2049995, -32'sd3055006, -32'sd2191441, -32'sd1710657, -32'sd898220, -32'sd1022416, 32'sd2224477, 32'sd3738632, 32'sd1643406, 32'sd546410, -32'sd3732858, -32'sd2105894, 32'sd1298269, -32'sd352275, 32'sd308119, -32'sd714762, -32'sd60656, 32'sd916635, -32'sd1381605, 32'sd75876, 32'sd164239, 32'sd400787, 32'sd613527, 32'sd416126, 32'sd156121, -32'sd635426, -32'sd1026412, -32'sd1598507, -32'sd2013825, -32'sd3100561, -32'sd1269005, -32'sd468678, -32'sd46669, 32'sd354164, 32'sd2023784, 32'sd2872545, -32'sd94464, -32'sd3862498, -32'sd4535246, -32'sd453994, 32'sd196028, 32'sd787546, -32'sd491506, -32'sd1952804, 32'sd1808140, -32'sd700704, -32'sd2179682, 32'sd581473, -32'sd152067, 32'sd318828, -32'sd162672, -32'sd369042, 32'sd2266790, -32'sd1044172, 32'sd1277489, -32'sd722036, -32'sd1452364, -32'sd2833032, -32'sd996419, 32'sd727299, 32'sd380845, 32'sd1593205, 32'sd2864115, 32'sd1743521, -32'sd2756693, -32'sd3907520, -32'sd1167752, 32'sd661350, 32'sd1310326, -32'sd29334, -32'sd1139099, -32'sd970148, -32'sd288604, 32'sd50770, -32'sd168968, -32'sd1127963, -32'sd617894, -32'sd779292, 32'sd1410314, -32'sd1848458, -32'sd693979, 32'sd106443, -32'sd435139, -32'sd133852, -32'sd2627933, -32'sd2201597, 32'sd1237074, 32'sd1348074, 32'sd973001, 32'sd608543, 32'sd1407409, -32'sd1044188, -32'sd1713662, -32'sd353146, 32'sd1772389, 32'sd342666, 32'sd754002, 32'sd562171, 32'sd421253, -32'sd357771, -32'sd777164, -32'sd1768995, 32'sd577549, -32'sd2169344, 32'sd124544, 32'sd1454030, 32'sd389508, -32'sd1405182, -32'sd1023794, -32'sd322385, -32'sd781436, -32'sd104631, -32'sd1651953, -32'sd2730639, 32'sd825693, 32'sd538115, -32'sd701083, 32'sd545937, 32'sd714320, 32'sd518944, -32'sd791394, -32'sd425747, -32'sd1222602, 32'sd1041247, 32'sd331445, -32'sd923284, -32'sd206124, 32'sd1334971, -32'sd740537, -32'sd598970, -32'sd977175, -32'sd180677, 32'sd146355, 32'sd297044, -32'sd534463, -32'sd1930871, -32'sd1843783, 32'sd1978767, -32'sd426373, -32'sd1681559, 32'sd281243, -32'sd756328, 32'sd976406, 32'sd112494, -32'sd2850240, -32'sd964410, -32'sd1205471, -32'sd1032838, -32'sd2144970, 32'sd544651, 32'sd287514, 32'sd692628, 32'sd2497005, 32'sd683955, 32'sd1810263, 32'sd1301978, 32'sd232357, -32'sd927346, 32'sd372873, 32'sd253127, 32'sd109267, 32'sd74005, 32'sd634012, -32'sd1104672, -32'sd1017125, 32'sd1724033, -32'sd629944, 32'sd457366, 32'sd272402, 32'sd994953, 32'sd1699969, 32'sd1659482, 32'sd90018, -32'sd988939, -32'sd2663497, 32'sd590405, -32'sd1524564, -32'sd107123, -32'sd1294684, 32'sd571866, -32'sd506248, 32'sd702064, 32'sd2319868, 32'sd2706714, 32'sd1526457, -32'sd233742, -32'sd651215, -32'sd143062, -32'sd1110498, 32'sd554465, 32'sd801335, -32'sd1198526, 32'sd98040, 32'sd984477, -32'sd1005585, 32'sd925563, -32'sd1408313, -32'sd955385, -32'sd796858, -32'sd387774, -32'sd956099, -32'sd132858, -32'sd1534265, -32'sd1544283, -32'sd1966085, -32'sd1536527, 32'sd468166, -32'sd625848, 32'sd494629, 32'sd2093286, 32'sd665307, 32'sd1271565, 32'sd2661212, 32'sd1347805, 32'sd572171, -32'sd7821, -32'sd574079, 32'sd594067, -32'sd859423, 32'sd485247, -32'sd2492281, 32'sd1370861, -32'sd786547, 32'sd464926, 32'sd2156818, -32'sd899114, 32'sd732369, -32'sd1000176, 32'sd1988917, 32'sd490027, -32'sd596533, 32'sd2763362, 32'sd337912, 32'sd105493, 32'sd382329, 32'sd1873701, 32'sd480945, 32'sd1065772, -32'sd620255, 32'sd653869, 32'sd166191, -32'sd607, 32'sd1296853, 32'sd456945, 32'sd1086743, 32'sd0, 32'sd115396, -32'sd565319, -32'sd1368221, -32'sd26024, 32'sd871312, -32'sd484487, -32'sd835514, 32'sd1350875, 32'sd949230, 32'sd1393669, 32'sd3606769, 32'sd2773199, -32'sd83272, 32'sd2330048, 32'sd1692996, 32'sd2048643, 32'sd1871341, -32'sd73253, 32'sd806811, -32'sd119820, 32'sd392850, 32'sd187348, 32'sd1358508, 32'sd409154, -32'sd329207, 32'sd121565, 32'sd512540, 32'sd1070192, 32'sd804956, -32'sd867311, -32'sd1454731, 32'sd1743451, -32'sd941066, -32'sd1364364, -32'sd1098493, 32'sd245807, 32'sd2970132, 32'sd1695541, 32'sd2222667, 32'sd225986, 32'sd444243, -32'sd149836, 32'sd1295165, 32'sd100248, -32'sd387358, 32'sd1270182, -32'sd101229, -32'sd2056314, 32'sd290299, 32'sd391367, 32'sd2157023, 32'sd892024, -32'sd416697, 32'sd808278, 32'sd891460, 32'sd1002027, 32'sd767201, -32'sd1535504, 32'sd1340377, 32'sd785543, 32'sd1251081, -32'sd1283489, -32'sd2021607, -32'sd512826, 32'sd1770349, 32'sd849401, 32'sd1784097, -32'sd1000983, -32'sd914963, 32'sd189851, 32'sd1670166, 32'sd311553, -32'sd1633371, 32'sd1102115, 32'sd1912209, 32'sd1464464, -32'sd507113, 32'sd605658, 32'sd1361232, 32'sd573588, -32'sd284108, -32'sd552984, 32'sd810894, 32'sd0, 32'sd1165419, -32'sd1532382, -32'sd648275, 32'sd18922, 32'sd84358, 32'sd281470, 32'sd588374, -32'sd1785988, 32'sd644130, 32'sd157734, 32'sd216390, -32'sd1304020, 32'sd719556, 32'sd1385272, -32'sd531771, -32'sd454293, -32'sd1321540, -32'sd2376373, 32'sd1125170, 32'sd1173237, 32'sd418524, 32'sd130487, 32'sd52781, -32'sd537608, 32'sd159076, -32'sd2158987, -32'sd229808, -32'sd109999, -32'sd525875, -32'sd1942560, 32'sd1253902, 32'sd2151098, -32'sd558546, 32'sd203434, 32'sd1684981, -32'sd545500, -32'sd890926, -32'sd439336, -32'sd91687, 32'sd1855890, 32'sd277009, 32'sd2046848, 32'sd1496913, -32'sd690652, 32'sd942156, 32'sd1090501, -32'sd1317900, 32'sd121089, -32'sd104463, -32'sd685913, 32'sd506765, -32'sd1643644, 32'sd370243, 32'sd425240, 32'sd142870, 32'sd602590, -32'sd44795, 32'sd1467765, 32'sd941052, 32'sd1236888, 32'sd1293415, 32'sd1180974, 32'sd1142372, -32'sd799038, -32'sd301064, 32'sd943012, -32'sd2447815, 32'sd2709980, 32'sd424177, -32'sd363919, 32'sd1947262, 32'sd1728402, 32'sd1027284, -32'sd419188, 32'sd35712, 32'sd564616, 32'sd40706, -32'sd1312170, -32'sd289501, -32'sd1101094, 32'sd26633, 32'sd111433, 32'sd930026, 32'sd0, 32'sd1259900, -32'sd453149, 32'sd837001, -32'sd1232940, -32'sd283677, 32'sd623851, 32'sd1457166, 32'sd2168036, 32'sd1704096, 32'sd89766, -32'sd477958, -32'sd1319761, -32'sd810072, 32'sd794163, 32'sd1825167, 32'sd367257, -32'sd1533101, -32'sd723666, 32'sd1167558, -32'sd397693, 32'sd546932, -32'sd536677, -32'sd559386, 32'sd302862, -32'sd677470, 32'sd119252, 32'sd0, 32'sd0, 32'sd0, -32'sd423493, -32'sd292606, -32'sd283670, 32'sd14040, 32'sd568697, 32'sd2654086, 32'sd1680341, 32'sd347625, -32'sd1904563, 32'sd71825, 32'sd1607129, -32'sd487139, -32'sd1173999, 32'sd2321044, 32'sd785212, 32'sd414372, -32'sd873685, -32'sd1256860, -32'sd473124, 32'sd744216, 32'sd1056708, 32'sd847621, 32'sd855720, 32'sd1293354, 32'sd1337808, 32'sd0, 32'sd0, 32'sd0, 32'sd1745196, 32'sd741660, 32'sd540210, 32'sd636025, -32'sd26454, -32'sd269029, 32'sd1405101, -32'sd1079386, -32'sd123375, 32'sd1513250, 32'sd475336, 32'sd644300, -32'sd623804, -32'sd1277790, 32'sd983775, 32'sd12334, -32'sd741789, 32'sd1376660, -32'sd962952, -32'sd134569, 32'sd274405, 32'sd958472, 32'sd567847, 32'sd416787, -32'sd204606, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd462017, 32'sd1039024, 32'sd537002, 32'sd1379159, 32'sd897427, 32'sd347846, -32'sd1620542, -32'sd1490122, -32'sd266391, -32'sd926479, -32'sd2245976, 32'sd90375, -32'sd2449275, -32'sd2929603, -32'sd1038609, 32'sd1839705, 32'sd1698756, 32'sd66880, 32'sd284894, 32'sd421113, -32'sd198447, 32'sd1424751, 32'sd294619, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1356864, 32'sd559698, 32'sd693288, 32'sd569436, 32'sd160054, 32'sd585645, -32'sd261055, -32'sd777203, -32'sd872599, 32'sd1097314, -32'sd73972, 32'sd1387913, -32'sd941872, 32'sd552963, 32'sd1555614, 32'sd2028969, 32'sd1040240, 32'sd271094, 32'sd999435, 32'sd986632, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd973816, -32'sd1561557, -32'sd434891, -32'sd129554, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd592176, -32'sd813986, -32'sd1268536, -32'sd1238902, -32'sd2225750, -32'sd224564, -32'sd119991, 32'sd333829, 32'sd339677, 32'sd1117793, 32'sd478997, -32'sd571193, 32'sd36107, -32'sd1317369, -32'sd17770, -32'sd1207148, -32'sd1856549, -32'sd1693015, 32'sd114564, 32'sd238636, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd700703, 32'sd296846, -32'sd1117865, -32'sd702090, 32'sd26720, -32'sd439259, 32'sd583057, 32'sd636732, 32'sd1947236, 32'sd342448, 32'sd938080, 32'sd951846, 32'sd933139, -32'sd1602999, -32'sd1490193, 32'sd229564, -32'sd1805071, -32'sd834593, -32'sd569330, -32'sd1292868, 32'sd680612, -32'sd860969, 32'sd23910, -32'sd942355, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd198021, -32'sd183603, -32'sd902133, 32'sd926998, -32'sd643381, 32'sd1418410, -32'sd5093, 32'sd472238, 32'sd1316187, 32'sd1019297, 32'sd841871, 32'sd1709516, 32'sd1261844, -32'sd1967903, -32'sd1126469, -32'sd1251144, -32'sd189718, 32'sd16220, -32'sd1102805, -32'sd1159071, -32'sd43549, -32'sd215684, 32'sd1797188, 32'sd685033, -32'sd370215, 32'sd0, 32'sd0, -32'sd1111313, -32'sd71430, 32'sd163758, -32'sd761229, -32'sd826207, 32'sd2217611, 32'sd3532285, 32'sd2806045, -32'sd863062, 32'sd1015448, 32'sd2345300, 32'sd1832428, 32'sd1012242, 32'sd1406342, 32'sd553816, 32'sd11275, -32'sd1116380, 32'sd296356, -32'sd60241, -32'sd163483, -32'sd619703, 32'sd798775, -32'sd30046, 32'sd627949, -32'sd1211820, -32'sd356808, -32'sd1474312, 32'sd0, 32'sd841782, 32'sd157360, 32'sd2314610, 32'sd1374375, -32'sd124771, -32'sd856139, -32'sd135580, -32'sd728420, 32'sd19019, 32'sd111817, -32'sd261350, 32'sd705631, 32'sd2570367, 32'sd1271946, 32'sd615666, 32'sd2264297, 32'sd1617222, 32'sd2406803, 32'sd2017574, -32'sd1370515, -32'sd792018, -32'sd1525332, -32'sd1277521, -32'sd577452, 32'sd945900, 32'sd1093608, 32'sd169514, 32'sd0, -32'sd1531778, -32'sd1326822, 32'sd1530579, 32'sd1559497, -32'sd77490, -32'sd2616805, -32'sd2450461, -32'sd1363411, -32'sd2560034, 32'sd329595, -32'sd460418, 32'sd1177195, 32'sd859918, 32'sd1596959, 32'sd1773303, 32'sd3440627, -32'sd614363, 32'sd2712855, -32'sd42782, -32'sd1148850, -32'sd3453322, -32'sd2901417, -32'sd2562246, -32'sd1402976, 32'sd1104834, -32'sd1135955, -32'sd169107, -32'sd238263, 32'sd603392, -32'sd1386093, -32'sd466842, -32'sd284290, -32'sd986118, -32'sd1637441, -32'sd849112, -32'sd278303, -32'sd2025029, -32'sd950794, -32'sd1230718, -32'sd552772, -32'sd1018209, 32'sd579570, 32'sd2493012, 32'sd943864, 32'sd23691, 32'sd1638875, -32'sd451491, 32'sd487966, -32'sd1411962, -32'sd796705, -32'sd781491, -32'sd1898710, -32'sd217940, -32'sd1853867, 32'sd82898, -32'sd1494858, 32'sd778219, -32'sd1005784, -32'sd58619, 32'sd317921, -32'sd1207722, -32'sd1193229, -32'sd925795, 32'sd821962, -32'sd1438339, -32'sd818899, -32'sd2467959, -32'sd2251442, -32'sd1959604, -32'sd116097, -32'sd1641924, 32'sd168356, 32'sd1544715, 32'sd2093029, 32'sd984608, -32'sd630919, -32'sd1870385, -32'sd1021553, -32'sd1285417, -32'sd1534245, -32'sd2187911, -32'sd326679, -32'sd1800752, -32'sd1747034, -32'sd971056, -32'sd835017, 32'sd1095241, -32'sd1255336, 32'sd563417, 32'sd235493, 32'sd208417, 32'sd1189691, -32'sd385062, -32'sd2502954, -32'sd728678, -32'sd2514851, -32'sd2452951, -32'sd2912878, -32'sd700420, -32'sd379624, 32'sd1254557, 32'sd2815510, 32'sd1966933, 32'sd1437795, -32'sd1222689, -32'sd1848358, -32'sd1979152, -32'sd3156029, -32'sd1278795, -32'sd289449, 32'sd385363, -32'sd978176, 32'sd76364, 32'sd798377, -32'sd7700, 32'sd741994, 32'sd1187812, 32'sd1811644, 32'sd774362, -32'sd129509, -32'sd1635807, -32'sd2010728, -32'sd3374654, -32'sd1917779, -32'sd1368030, 32'sd184067, -32'sd989804, -32'sd1009006, 32'sd1499596, 32'sd1801437, 32'sd715828, 32'sd450828, 32'sd1230572, -32'sd1032666, -32'sd755425, -32'sd1687586, 32'sd724318, -32'sd1259680, -32'sd1233152, -32'sd1228151, -32'sd754579, -32'sd1913195, -32'sd110019, -32'sd791447, 32'sd1011300, 32'sd56564, -32'sd364083, -32'sd3640643, -32'sd1978351, -32'sd1352335, -32'sd25451, -32'sd378115, 32'sd945593, -32'sd340759, -32'sd1043175, -32'sd732177, 32'sd1401325, 32'sd292838, -32'sd523897, 32'sd131233, -32'sd618990, -32'sd1355682, -32'sd1301909, -32'sd2780359, 32'sd349639, 32'sd297184, -32'sd1739690, -32'sd893241, -32'sd1235367, 32'sd95028, -32'sd1907031, 32'sd587785, -32'sd2819320, -32'sd846112, -32'sd1503596, -32'sd3084051, -32'sd574215, -32'sd691375, -32'sd1729039, -32'sd1580782, -32'sd1292938, 32'sd1160377, -32'sd1393333, -32'sd242060, 32'sd854812, -32'sd3156497, 32'sd288243, 32'sd49140, -32'sd1918382, -32'sd2370321, -32'sd1631364, -32'sd1324764, 32'sd757353, -32'sd2033474, -32'sd1411189, -32'sd585804, -32'sd366390, -32'sd813840, 32'sd864608, -32'sd1090483, -32'sd1537407, -32'sd2311175, -32'sd405012, 32'sd1618649, 32'sd893188, -32'sd2048006, -32'sd2382292, -32'sd1650993, -32'sd1575749, 32'sd1702594, -32'sd1968276, -32'sd627414, 32'sd1122485, -32'sd1054129, 32'sd2226105, 32'sd1745449, -32'sd769655, -32'sd1042044, -32'sd850043, -32'sd58651, 32'sd1661819, -32'sd679979, -32'sd514775, -32'sd1235590, -32'sd1767983, -32'sd1580095, -32'sd78495, 32'sd691763, -32'sd1472685, -32'sd1565692, -32'sd840015, -32'sd667126, -32'sd1107302, -32'sd1591922, -32'sd1835455, -32'sd1544985, -32'sd740294, 32'sd1733557, -32'sd1298229, -32'sd728782, -32'sd761882, 32'sd533917, 32'sd154793, 32'sd698715, -32'sd989134, -32'sd1604286, -32'sd1385273, -32'sd2108525, 32'sd697091, 32'sd1241183, 32'sd61351, -32'sd217013, -32'sd100347, -32'sd396636, 32'sd2013882, -32'sd913048, 32'sd358238, -32'sd1131700, -32'sd1194713, -32'sd1938527, 32'sd532289, -32'sd1550206, 32'sd182667, -32'sd642117, 32'sd1285709, 32'sd2237540, -32'sd514552, 32'sd819871, -32'sd472189, 32'sd761437, -32'sd1821274, -32'sd1648517, 32'sd58352, 32'sd1743527, 32'sd1432888, -32'sd37134, 32'sd488097, -32'sd223573, 32'sd500887, -32'sd862731, -32'sd1370447, -32'sd2883231, 32'sd55624, -32'sd170802, -32'sd1596891, -32'sd785413, -32'sd2335658, -32'sd487084, -32'sd706881, -32'sd957183, -32'sd1743268, 32'sd386078, 32'sd714971, -32'sd742026, -32'sd2252683, -32'sd1417061, 32'sd350008, -32'sd125058, 32'sd601249, -32'sd859809, -32'sd92139, 32'sd644104, 32'sd131344, -32'sd54394, 32'sd299382, -32'sd33719, -32'sd1758562, 32'sd0, -32'sd1827177, -32'sd2282887, -32'sd3335, -32'sd602643, -32'sd225687, -32'sd550075, 32'sd192387, -32'sd449573, -32'sd1216547, -32'sd366907, -32'sd452750, -32'sd1091053, -32'sd1241919, -32'sd1631037, -32'sd196966, 32'sd497122, -32'sd212832, -32'sd132245, 32'sd340346, -32'sd2028008, -32'sd43074, 32'sd621264, -32'sd1046377, 32'sd1699242, 32'sd1543688, -32'sd960861, -32'sd1598556, -32'sd618643, -32'sd1231672, -32'sd965788, -32'sd57184, 32'sd950301, -32'sd567221, 32'sd387346, -32'sd2386148, 32'sd1026633, 32'sd1481928, 32'sd1467919, -32'sd507618, -32'sd2530167, -32'sd1173732, -32'sd1047782, 32'sd448146, 32'sd749602, 32'sd764988, 32'sd862824, -32'sd625689, 32'sd189780, -32'sd471921, -32'sd1389356, -32'sd368038, 32'sd430084, 32'sd1240619, -32'sd306530, -32'sd1543646, -32'sd508355, -32'sd809957, -32'sd947169, -32'sd15455, -32'sd764877, -32'sd381345, -32'sd712268, -32'sd177909, -32'sd1583419, 32'sd1461958, 32'sd680870, -32'sd1685787, -32'sd1271012, -32'sd301130, -32'sd576349, 32'sd1475669, 32'sd1737010, 32'sd1674103, 32'sd868673, 32'sd161840, -32'sd1322926, -32'sd103995, -32'sd1017069, -32'sd1485646, -32'sd1053232, -32'sd1470981, 32'sd1197658, -32'sd527812, 32'sd0, 32'sd372072, -32'sd388924, 32'sd1110874, -32'sd1045812, 32'sd164421, -32'sd392463, -32'sd507950, 32'sd97446, 32'sd1889757, 32'sd1019661, 32'sd500237, 32'sd558487, 32'sd1314551, 32'sd893725, 32'sd2002381, 32'sd1415690, -32'sd40118, 32'sd1715326, -32'sd435233, 32'sd412880, -32'sd1438924, -32'sd1386412, -32'sd235649, -32'sd753100, -32'sd876721, -32'sd1036167, -32'sd1306118, -32'sd410998, 32'sd1576873, -32'sd10377, 32'sd1213218, 32'sd338718, -32'sd1453128, -32'sd781193, 32'sd1426902, -32'sd598144, 32'sd97350, 32'sd1826691, 32'sd180440, 32'sd1049317, 32'sd3450163, 32'sd2410127, 32'sd394721, -32'sd91957, 32'sd404088, 32'sd414165, 32'sd1147123, -32'sd1127630, -32'sd1226614, -32'sd330943, 32'sd18141, 32'sd320661, 32'sd19062, 32'sd301166, -32'sd394929, -32'sd657542, 32'sd523515, -32'sd703580, -32'sd2018433, 32'sd180943, -32'sd446762, -32'sd1752401, -32'sd1474564, -32'sd513641, 32'sd1324989, -32'sd604297, 32'sd1648825, 32'sd606591, 32'sd2156885, 32'sd852180, 32'sd1968421, 32'sd370791, 32'sd358156, -32'sd1541916, 32'sd1581909, 32'sd572469, 32'sd1755160, 32'sd165670, 32'sd800033, 32'sd1484529, 32'sd192509, -32'sd624253, -32'sd687414, 32'sd0, 32'sd62206, 32'sd85512, -32'sd125988, -32'sd1241041, 32'sd1155472, -32'sd1552336, 32'sd518909, 32'sd1811043, 32'sd1361859, 32'sd415546, 32'sd3194022, 32'sd185760, 32'sd1242383, -32'sd307445, 32'sd2599581, 32'sd1863833, 32'sd50536, 32'sd290254, -32'sd1666646, 32'sd1797519, 32'sd431646, 32'sd541484, -32'sd278763, -32'sd328653, 32'sd733364, -32'sd2036494, 32'sd0, 32'sd0, 32'sd0, 32'sd203036, -32'sd292211, -32'sd1883086, 32'sd1259992, 32'sd1264383, 32'sd195564, 32'sd81221, 32'sd2139250, 32'sd2807837, 32'sd2434643, 32'sd2055783, 32'sd650338, 32'sd757596, 32'sd1108526, 32'sd87390, 32'sd2619577, 32'sd184240, -32'sd109903, 32'sd1218607, 32'sd504254, -32'sd3152377, -32'sd1907146, 32'sd754323, 32'sd1058785, -32'sd1386836, 32'sd0, 32'sd0, 32'sd0, 32'sd1104144, -32'sd597682, 32'sd232578, 32'sd12378, 32'sd2187258, 32'sd1924541, 32'sd1248876, 32'sd361196, 32'sd1903157, -32'sd601443, 32'sd1212538, 32'sd1113600, 32'sd195686, -32'sd1797924, 32'sd919429, 32'sd139569, 32'sd1301334, -32'sd217000, 32'sd645166, 32'sd293124, 32'sd927071, -32'sd689951, -32'sd399390, -32'sd1215172, -32'sd1223621, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd512649, 32'sd595655, 32'sd538159, -32'sd2139762, -32'sd1833275, -32'sd1484505, -32'sd2511954, -32'sd762529, -32'sd2310251, -32'sd639662, -32'sd1162475, -32'sd2842172, -32'sd2043691, -32'sd1059464, -32'sd657566, -32'sd634962, -32'sd381293, -32'sd1571758, -32'sd2247666, -32'sd1454831, -32'sd1502953, -32'sd321283, 32'sd549114, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1570300, -32'sd1850069, -32'sd1111543, -32'sd707387, -32'sd1666960, -32'sd646813, 32'sd289233, 32'sd427897, -32'sd1431494, -32'sd1557427, -32'sd435546, -32'sd1913255, -32'sd665815, 32'sd91252, 32'sd8861, -32'sd295723, -32'sd1880733, -32'sd534062, -32'sd918237, -32'sd1272466, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd705694, 32'sd144601, -32'sd432328, -32'sd13324, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd423586, -32'sd248896, 32'sd1246126, 32'sd289244, -32'sd286687, 32'sd410498, -32'sd225603, 32'sd1354015, -32'sd1213557, -32'sd488532, -32'sd193600, -32'sd839666, 32'sd58471, 32'sd200400, -32'sd522909, 32'sd1038688, 32'sd702770, 32'sd598412, 32'sd63083, 32'sd453782, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd451438, -32'sd270010, 32'sd505109, -32'sd606756, 32'sd137066, 32'sd424330, -32'sd1341719, 32'sd91763, 32'sd578137, 32'sd761338, 32'sd232549, 32'sd582706, -32'sd120895, 32'sd587796, -32'sd576554, 32'sd873362, 32'sd1787187, 32'sd1520881, 32'sd1786402, 32'sd1969343, -32'sd838618, -32'sd133093, 32'sd459790, 32'sd2185841, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1859259, 32'sd434484, 32'sd262573, 32'sd571162, -32'sd659066, -32'sd672648, -32'sd1543285, 32'sd811688, 32'sd726997, 32'sd474790, -32'sd205415, 32'sd799935, -32'sd947335, 32'sd640734, 32'sd569325, -32'sd1511621, -32'sd224389, 32'sd220287, 32'sd733213, -32'sd333159, 32'sd1648436, 32'sd1064618, 32'sd884899, 32'sd686196, 32'sd952122, 32'sd0, 32'sd0, 32'sd426617, 32'sd1166747, 32'sd535050, -32'sd1137963, 32'sd1412354, 32'sd80759, 32'sd152318, -32'sd879915, -32'sd2408257, -32'sd2944, -32'sd2558612, -32'sd74610, -32'sd1224232, -32'sd154167, -32'sd1637827, 32'sd694669, 32'sd1926902, 32'sd1307411, 32'sd901533, 32'sd799061, -32'sd1209475, 32'sd2287394, -32'sd75827, -32'sd933262, -32'sd2536531, 32'sd183827, 32'sd912975, 32'sd0, 32'sd983218, 32'sd400188, -32'sd877601, 32'sd709092, -32'sd59472, -32'sd606852, 32'sd990908, -32'sd383315, -32'sd1428490, -32'sd3069180, -32'sd3115556, -32'sd1671814, 32'sd799847, 32'sd469171, 32'sd1688572, -32'sd830255, 32'sd1582244, -32'sd268880, 32'sd177315, 32'sd260934, 32'sd441015, 32'sd1063741, -32'sd186327, 32'sd453110, -32'sd639611, -32'sd97487, -32'sd1170919, 32'sd0, 32'sd880456, 32'sd850536, -32'sd323892, 32'sd1256189, 32'sd1245010, -32'sd2078528, -32'sd876222, -32'sd801386, -32'sd2215320, -32'sd984675, -32'sd552691, -32'sd171256, -32'sd1626807, -32'sd1177681, -32'sd1442079, 32'sd547447, -32'sd764179, 32'sd1498487, 32'sd1309632, -32'sd1094707, 32'sd1179580, 32'sd322645, 32'sd1145666, -32'sd1396076, 32'sd691548, -32'sd1020094, 32'sd1421707, 32'sd1471552, -32'sd136462, -32'sd31458, -32'sd419011, 32'sd840419, 32'sd754967, -32'sd180282, -32'sd189949, -32'sd359548, -32'sd1049052, -32'sd1596435, -32'sd668235, 32'sd620133, -32'sd1281207, 32'sd214601, 32'sd796187, 32'sd825744, 32'sd975799, 32'sd432462, 32'sd172733, -32'sd183660, -32'sd584291, 32'sd1518249, -32'sd1219445, -32'sd276081, 32'sd1009493, 32'sd657292, -32'sd409538, 32'sd345636, 32'sd173446, 32'sd1315014, 32'sd298566, 32'sd996707, 32'sd480996, 32'sd1859859, 32'sd362046, -32'sd269680, -32'sd2458297, -32'sd295103, -32'sd2311489, -32'sd307267, 32'sd1398390, -32'sd1698278, -32'sd736771, 32'sd1828669, 32'sd54639, -32'sd1232408, 32'sd1165175, -32'sd340521, -32'sd1908815, 32'sd965978, 32'sd1425320, -32'sd919663, -32'sd197693, -32'sd598106, 32'sd2719, 32'sd262588, 32'sd379054, -32'sd783930, 32'sd1127255, 32'sd324370, 32'sd2094210, 32'sd140886, 32'sd1669751, -32'sd684428, -32'sd1714749, -32'sd39397, -32'sd809219, -32'sd1921732, -32'sd1527073, -32'sd2470751, -32'sd936442, 32'sd62375, -32'sd2442043, -32'sd1302399, 32'sd1240438, -32'sd332018, -32'sd488509, 32'sd201072, 32'sd799523, 32'sd717031, 32'sd1039802, -32'sd325866, -32'sd438762, -32'sd508824, -32'sd678483, 32'sd1341747, 32'sd339214, -32'sd558223, 32'sd2357189, 32'sd3396673, 32'sd2082085, -32'sd115876, 32'sd1957742, 32'sd1146303, 32'sd865327, -32'sd1174017, -32'sd1129109, -32'sd1341070, -32'sd1872588, -32'sd761239, -32'sd1548073, -32'sd1175779, -32'sd373230, 32'sd720903, 32'sd482654, 32'sd1763493, 32'sd511548, -32'sd364570, -32'sd1322258, -32'sd1347280, 32'sd1368348, -32'sd582479, -32'sd921905, 32'sd862283, 32'sd62133, 32'sd1876644, 32'sd1189510, 32'sd3857515, 32'sd1229138, -32'sd75816, 32'sd2210971, 32'sd1374613, 32'sd1867849, -32'sd1030413, -32'sd1335280, -32'sd2581762, -32'sd1073354, 32'sd579227, 32'sd440346, -32'sd691655, 32'sd1437309, 32'sd2348701, 32'sd234518, 32'sd1410181, 32'sd241384, -32'sd147423, -32'sd1200487, -32'sd1665385, -32'sd776183, 32'sd786853, 32'sd149930, -32'sd1050402, -32'sd1461788, 32'sd1014050, 32'sd1399096, 32'sd1939193, 32'sd3352934, 32'sd1444428, 32'sd788661, -32'sd199515, 32'sd568288, 32'sd800516, -32'sd149912, -32'sd1365263, -32'sd2279964, 32'sd778296, 32'sd798196, 32'sd1160400, 32'sd136446, -32'sd646052, 32'sd777954, 32'sd217787, -32'sd1217394, -32'sd1219773, -32'sd585044, -32'sd1913630, 32'sd183289, 32'sd205764, -32'sd97981, 32'sd31724, -32'sd969028, -32'sd1015209, -32'sd2782704, -32'sd296362, 32'sd87042, 32'sd2604571, 32'sd2673253, -32'sd611061, -32'sd472446, -32'sd2943707, -32'sd2246016, -32'sd670455, -32'sd38015, -32'sd496032, -32'sd1154601, 32'sd1879522, -32'sd585858, -32'sd1441545, 32'sd563590, 32'sd103220, -32'sd502952, -32'sd502671, -32'sd1189696, -32'sd429573, 32'sd1666381, 32'sd470148, 32'sd771451, 32'sd945941, 32'sd179790, -32'sd1246837, -32'sd865736, 32'sd414236, -32'sd909625, -32'sd1228703, -32'sd2521300, -32'sd2664658, -32'sd2110318, -32'sd3632664, 32'sd204851, 32'sd2365380, -32'sd1378066, 32'sd281173, -32'sd388314, -32'sd2121163, -32'sd707488, -32'sd242620, -32'sd2716149, -32'sd2264782, 32'sd758572, -32'sd472029, 32'sd575096, 32'sd2600487, 32'sd1186171, 32'sd723692, -32'sd1257116, 32'sd70817, 32'sd1127995, 32'sd802465, -32'sd1513679, -32'sd676102, -32'sd1918745, -32'sd3738668, -32'sd3633054, -32'sd4426837, -32'sd4044321, -32'sd1748528, 32'sd1122065, 32'sd2943951, -32'sd716065, -32'sd501764, -32'sd298068, -32'sd75597, -32'sd488249, -32'sd2160924, -32'sd667494, -32'sd28224, 32'sd891179, 32'sd666096, 32'sd1998109, 32'sd227531, 32'sd475310, 32'sd826465, -32'sd1041164, -32'sd504678, -32'sd377243, 32'sd1690438, -32'sd39606, -32'sd833109, -32'sd998691, -32'sd4182661, -32'sd5057989, -32'sd3982312, -32'sd1673190, 32'sd83660, 32'sd2490783, 32'sd2493386, 32'sd510937, 32'sd1970465, -32'sd351496, -32'sd579849, -32'sd483716, -32'sd1377445, -32'sd994277, 32'sd2400, 32'sd1883728, 32'sd286680, -32'sd497026, -32'sd1731256, -32'sd727553, 32'sd0, 32'sd765704, 32'sd244311, -32'sd838004, -32'sd1217940, -32'sd1958127, -32'sd2104581, -32'sd4305550, -32'sd2938629, -32'sd3614801, -32'sd1856476, 32'sd1404312, 32'sd4483042, 32'sd975407, 32'sd1652202, -32'sd761931, 32'sd1097266, 32'sd1914879, 32'sd1276020, -32'sd557177, 32'sd592350, -32'sd2632216, -32'sd174380, 32'sd375183, -32'sd234915, -32'sd1708365, -32'sd1832354, 32'sd518832, -32'sd386120, 32'sd1157441, -32'sd1701468, -32'sd600137, 32'sd726230, -32'sd1370655, -32'sd1284271, -32'sd5121529, -32'sd4304533, -32'sd1731618, 32'sd2028843, 32'sd2000083, 32'sd4520506, 32'sd3402863, -32'sd1448824, -32'sd1565063, -32'sd2328814, -32'sd210492, 32'sd167521, 32'sd1127009, -32'sd1872642, -32'sd2470184, -32'sd2080542, -32'sd1024944, 32'sd834521, -32'sd179212, -32'sd846830, -32'sd511168, 32'sd476497, -32'sd1409549, -32'sd881620, 32'sd1355214, -32'sd737832, -32'sd2593307, -32'sd2601662, -32'sd1727602, -32'sd1208386, 32'sd810080, 32'sd930388, 32'sd2421312, 32'sd2838129, 32'sd1587460, -32'sd1545814, -32'sd2069038, -32'sd471979, 32'sd623250, 32'sd495022, 32'sd570994, 32'sd311659, -32'sd219178, -32'sd1462079, -32'sd1288820, -32'sd221786, -32'sd1860299, -32'sd649582, 32'sd860607, 32'sd0, -32'sd528705, 32'sd282972, 32'sd207141, -32'sd1029473, -32'sd2384213, -32'sd2582339, -32'sd1045074, -32'sd485777, -32'sd266386, 32'sd1569572, 32'sd3352276, 32'sd4407853, -32'sd242977, 32'sd368479, 32'sd502964, 32'sd762278, 32'sd820279, 32'sd2177804, 32'sd324501, -32'sd1463449, 32'sd829564, -32'sd1672314, -32'sd1084761, -32'sd1216249, -32'sd792610, -32'sd844786, 32'sd727251, 32'sd1653223, 32'sd847494, 32'sd634077, -32'sd306612, -32'sd1539219, 32'sd38102, 32'sd627184, -32'sd659403, -32'sd2836033, -32'sd166266, 32'sd492027, 32'sd1216860, 32'sd2534350, 32'sd260817, 32'sd464364, 32'sd1023849, 32'sd937546, 32'sd1469121, 32'sd1235167, 32'sd1736958, -32'sd146055, 32'sd233880, 32'sd780333, 32'sd1602187, 32'sd2380317, 32'sd884391, 32'sd1342228, 32'sd422237, 32'sd917714, -32'sd509920, -32'sd426918, -32'sd999698, 32'sd440726, -32'sd185610, -32'sd260041, -32'sd736935, -32'sd2705404, 32'sd198620, -32'sd214255, 32'sd166367, 32'sd1255626, 32'sd267800, -32'sd871131, -32'sd650366, 32'sd1209550, 32'sd2206860, 32'sd2688718, 32'sd426708, -32'sd1242673, -32'sd1014948, 32'sd1943598, 32'sd669805, -32'sd19080, 32'sd903534, 32'sd1202718, 32'sd632178, 32'sd0, 32'sd834220, 32'sd640756, -32'sd1017068, -32'sd1835516, -32'sd499872, 32'sd562227, 32'sd381265, -32'sd1766205, 32'sd571085, -32'sd1140533, 32'sd899296, 32'sd524173, 32'sd2264072, 32'sd770718, 32'sd2770837, 32'sd1234413, 32'sd1464291, 32'sd66457, 32'sd1579713, 32'sd464650, -32'sd1991159, -32'sd31705, 32'sd1676950, 32'sd538476, 32'sd705058, -32'sd378533, 32'sd0, 32'sd0, 32'sd0, -32'sd35110, -32'sd1332986, -32'sd2626265, -32'sd845240, -32'sd48586, -32'sd1531309, -32'sd260398, -32'sd1371655, -32'sd1813715, 32'sd133404, 32'sd1818555, 32'sd771614, 32'sd1594667, 32'sd527503, 32'sd462082, -32'sd630097, 32'sd1199718, 32'sd1487808, 32'sd1386240, -32'sd919383, 32'sd77617, 32'sd856428, 32'sd1064762, 32'sd1247244, 32'sd588986, 32'sd0, 32'sd0, 32'sd0, -32'sd390872, 32'sd553341, 32'sd955377, 32'sd344874, 32'sd2122157, -32'sd874033, -32'sd751452, -32'sd291591, -32'sd1102676, 32'sd154274, 32'sd1277200, -32'sd41678, 32'sd1778438, 32'sd2214157, -32'sd857208, 32'sd53683, -32'sd1975423, -32'sd569420, -32'sd439771, 32'sd206746, -32'sd1539440, -32'sd815678, -32'sd2335, -32'sd10166, -32'sd37596, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd564589, -32'sd527557, -32'sd102377, 32'sd762610, -32'sd780930, 32'sd1491551, -32'sd150611, 32'sd14404, 32'sd1207867, -32'sd395071, -32'sd697298, -32'sd2354463, -32'sd1158206, -32'sd1568074, 32'sd640497, 32'sd881808, 32'sd621137, 32'sd711242, -32'sd1031629, 32'sd2065149, 32'sd611890, -32'sd602395, 32'sd701059, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1736979, 32'sd1017288, -32'sd174684, 32'sd1699447, -32'sd866978, -32'sd190349, -32'sd851515, 32'sd85394, 32'sd970195, 32'sd1869620, 32'sd2244950, 32'sd1088509, 32'sd2991891, 32'sd2009962, 32'sd843243, 32'sd1194753, 32'sd99244, 32'sd402354, 32'sd216439, 32'sd56233, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd283679, 32'sd754835, 32'sd2041494, 32'sd1490764, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd221925, 32'sd58053, 32'sd975736, -32'sd871052, 32'sd756060, 32'sd785149, 32'sd1176411, 32'sd1122391, -32'sd319383, -32'sd895046, 32'sd690014, -32'sd616917, 32'sd1433064, 32'sd919, 32'sd449979, 32'sd868137, -32'sd411890, 32'sd1399979, 32'sd1502027, 32'sd1247857, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd967815, 32'sd872189, -32'sd1927391, 32'sd1327659, 32'sd1283547, 32'sd1231718, 32'sd289700, 32'sd210145, 32'sd349639, -32'sd612756, -32'sd333506, -32'sd956647, -32'sd569017, -32'sd1908017, 32'sd384967, 32'sd2394142, 32'sd1785537, -32'sd2606514, -32'sd2050925, 32'sd1395234, 32'sd513857, 32'sd1131184, 32'sd1198792, 32'sd1424761, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1357792, -32'sd337960, -32'sd373180, 32'sd382959, 32'sd131038, -32'sd947155, 32'sd15680, -32'sd525746, 32'sd917767, 32'sd202268, 32'sd1133659, 32'sd1439094, 32'sd1064899, -32'sd1335059, 32'sd460653, 32'sd282825, 32'sd1349441, 32'sd752987, -32'sd951077, 32'sd788218, 32'sd669303, -32'sd987066, -32'sd484587, 32'sd442068, -32'sd1681376, 32'sd0, 32'sd0, -32'sd24294, 32'sd717541, 32'sd208556, 32'sd1363392, -32'sd279513, 32'sd1025537, -32'sd406651, 32'sd337467, -32'sd845366, 32'sd113046, 32'sd1487110, 32'sd1785180, 32'sd1805955, -32'sd301208, -32'sd514746, -32'sd21524, -32'sd2102738, -32'sd1116215, -32'sd2194165, -32'sd560659, 32'sd123241, -32'sd1056990, 32'sd102941, 32'sd1044493, -32'sd145448, -32'sd967415, 32'sd1299714, 32'sd0, 32'sd863953, -32'sd580386, -32'sd770189, 32'sd1443323, 32'sd970452, 32'sd587912, 32'sd764614, 32'sd2112846, 32'sd159516, 32'sd2622762, 32'sd3620018, 32'sd3782548, 32'sd962460, 32'sd2407832, -32'sd619090, 32'sd1020505, -32'sd350092, -32'sd3403528, -32'sd2681401, -32'sd1036519, 32'sd1016966, -32'sd223028, 32'sd1660566, 32'sd870151, 32'sd346262, -32'sd1259732, 32'sd602804, 32'sd0, 32'sd691914, 32'sd178385, 32'sd977767, -32'sd331282, 32'sd1057675, 32'sd1291896, 32'sd1242309, 32'sd2830588, 32'sd1846063, 32'sd3850560, 32'sd1691989, 32'sd3274709, 32'sd1298420, -32'sd1267416, 32'sd303097, -32'sd1162180, 32'sd774601, -32'sd475246, 32'sd430241, -32'sd677495, -32'sd1197712, 32'sd868384, -32'sd53023, 32'sd2223512, 32'sd974036, -32'sd886272, -32'sd43123, 32'sd2024271, 32'sd794938, 32'sd828, 32'sd919477, 32'sd1945624, 32'sd2106464, 32'sd410399, 32'sd488018, 32'sd683566, 32'sd3668624, 32'sd3544429, 32'sd2116300, 32'sd814489, 32'sd443145, -32'sd2413456, -32'sd2466494, -32'sd67235, 32'sd2022927, 32'sd800789, -32'sd690775, -32'sd75271, -32'sd980112, -32'sd522891, -32'sd686688, 32'sd3636577, 32'sd1586492, 32'sd154689, -32'sd165484, 32'sd1227103, 32'sd1511260, -32'sd105731, 32'sd2229857, 32'sd1852219, 32'sd1212424, 32'sd2278122, 32'sd1710820, 32'sd174573, 32'sd2521825, 32'sd2062210, 32'sd391147, 32'sd826280, 32'sd2350215, -32'sd1351596, -32'sd1984652, 32'sd145308, 32'sd1258896, 32'sd2568153, -32'sd115716, 32'sd457571, -32'sd2247156, -32'sd129228, 32'sd2127989, 32'sd3119535, 32'sd548337, 32'sd17362, 32'sd140051, 32'sd722266, 32'sd22393, 32'sd2541040, 32'sd2183814, -32'sd933365, -32'sd1067844, -32'sd2731186, -32'sd2351162, -32'sd1309790, -32'sd297199, 32'sd8724, 32'sd7136, 32'sd848370, -32'sd328208, 32'sd345745, -32'sd699561, -32'sd1319881, 32'sd3006522, -32'sd651188, -32'sd1769794, 32'sd290753, 32'sd1848449, -32'sd395668, 32'sd2313849, 32'sd980555, 32'sd548681, -32'sd382715, 32'sd1195906, 32'sd1347691, 32'sd635384, -32'sd295404, 32'sd1592669, -32'sd956207, -32'sd1692978, -32'sd992176, -32'sd3089584, -32'sd2917381, -32'sd1295477, 32'sd956964, -32'sd530094, -32'sd1951086, -32'sd1530818, -32'sd3192700, 32'sd925330, 32'sd390059, 32'sd2388595, 32'sd215425, -32'sd277168, -32'sd778024, -32'sd697708, 32'sd1241596, 32'sd934778, 32'sd227850, -32'sd560520, 32'sd256253, -32'sd118059, 32'sd1552637, -32'sd225536, 32'sd683905, -32'sd760508, -32'sd1634898, -32'sd1086894, -32'sd2776390, -32'sd2413979, -32'sd1352268, 32'sd249886, -32'sd308256, -32'sd1537592, 32'sd164287, -32'sd460196, -32'sd1850502, -32'sd1008829, -32'sd175823, 32'sd74668, 32'sd757254, -32'sd1499428, -32'sd1840258, 32'sd57678, 32'sd232739, -32'sd306649, 32'sd55845, 32'sd211834, 32'sd12747, 32'sd389078, 32'sd910024, 32'sd1216535, 32'sd1093120, -32'sd668770, -32'sd540711, -32'sd3322244, -32'sd3599508, -32'sd3723587, -32'sd2085229, -32'sd3737594, -32'sd2349237, -32'sd1884429, -32'sd436946, 32'sd470785, -32'sd1739510, 32'sd804310, 32'sd2598480, 32'sd828903, 32'sd1064699, 32'sd366352, 32'sd492655, -32'sd120972, -32'sd126836, 32'sd860373, 32'sd1735991, 32'sd79544, -32'sd317339, -32'sd81856, 32'sd1159953, 32'sd1463188, 32'sd1193073, 32'sd493974, -32'sd1813737, -32'sd2600435, -32'sd4292070, -32'sd2974780, -32'sd2488724, -32'sd2843523, 32'sd841933, 32'sd495102, 32'sd1364627, 32'sd1765779, -32'sd1943273, -32'sd660190, 32'sd1002649, -32'sd2180308, -32'sd402268, 32'sd402996, 32'sd746589, 32'sd1209207, 32'sd633170, -32'sd112286, 32'sd762520, -32'sd2276427, -32'sd1114525, 32'sd568223, -32'sd381147, -32'sd829617, 32'sd531313, -32'sd949774, 32'sd1427949, -32'sd821325, -32'sd654053, -32'sd3676869, -32'sd3804343, -32'sd2940701, 32'sd1726749, 32'sd1992169, 32'sd1821123, 32'sd346373, -32'sd530351, -32'sd104336, -32'sd2546376, -32'sd1030970, -32'sd100401, 32'sd75573, -32'sd1007780, 32'sd1186494, -32'sd1519629, -32'sd1614173, -32'sd1196010, 32'sd2304199, -32'sd810007, -32'sd721952, 32'sd1541104, 32'sd363558, 32'sd1251470, 32'sd1810400, 32'sd709060, -32'sd1058199, 32'sd704452, 32'sd233495, -32'sd2260268, -32'sd22672, 32'sd1588860, 32'sd2282203, -32'sd516322, 32'sd148903, -32'sd326819, 32'sd1150331, -32'sd664464, 32'sd69168, 32'sd1421047, 32'sd69315, 32'sd178510, 32'sd1186591, -32'sd126893, 32'sd1450070, 32'sd1170645, 32'sd2951798, 32'sd931038, -32'sd433127, 32'sd1186689, -32'sd1394530, 32'sd603666, 32'sd885926, -32'sd1432379, 32'sd1641159, -32'sd245506, 32'sd2214371, 32'sd435606, 32'sd1249715, 32'sd2018431, -32'sd667665, -32'sd533873, 32'sd676747, 32'sd343101, -32'sd731538, -32'sd629637, 32'sd2351626, 32'sd1239462, 32'sd1710983, -32'sd193346, 32'sd2091675, 32'sd704911, 32'sd305462, 32'sd676969, 32'sd1521867, 32'sd983095, 32'sd413271, 32'sd0, 32'sd135762, -32'sd336240, -32'sd364689, 32'sd650593, -32'sd451700, -32'sd106493, 32'sd992155, -32'sd399111, 32'sd2550367, 32'sd440496, 32'sd357965, 32'sd246138, -32'sd9279, -32'sd563513, -32'sd1176874, -32'sd82287, -32'sd2026908, -32'sd519532, 32'sd797579, 32'sd1073979, 32'sd993323, -32'sd104002, -32'sd366384, -32'sd570168, 32'sd812628, 32'sd33697, -32'sd276241, -32'sd242782, -32'sd197300, -32'sd433430, 32'sd149862, 32'sd1308776, 32'sd117122, -32'sd1024712, 32'sd301462, -32'sd70058, 32'sd1059815, 32'sd535317, 32'sd1212184, 32'sd743685, -32'sd346004, -32'sd2288859, -32'sd62896, -32'sd2380007, -32'sd972636, 32'sd167816, -32'sd721622, -32'sd1056557, -32'sd1753390, -32'sd267684, 32'sd637969, 32'sd900286, 32'sd375051, 32'sd741522, 32'sd445795, 32'sd910128, 32'sd236573, 32'sd1206054, 32'sd1658154, 32'sd346306, 32'sd260751, -32'sd2204017, -32'sd1271999, -32'sd905572, -32'sd10031, 32'sd578102, 32'sd3722578, 32'sd257579, 32'sd1163264, 32'sd770857, 32'sd1175470, -32'sd1569495, -32'sd619038, 32'sd578526, 32'sd540391, -32'sd14050, -32'sd789195, 32'sd1330828, 32'sd998206, 32'sd608839, -32'sd13043, 32'sd183215, -32'sd251757, 32'sd0, 32'sd966439, 32'sd256252, 32'sd828008, -32'sd1724052, -32'sd176216, -32'sd2199794, -32'sd2220921, 32'sd124298, -32'sd1354929, 32'sd1282438, 32'sd2102853, 32'sd304010, 32'sd735080, -32'sd897914, 32'sd279227, -32'sd1978467, -32'sd650827, -32'sd2007899, -32'sd1354441, -32'sd1555958, -32'sd679611, -32'sd1263937, 32'sd575507, 32'sd21426, 32'sd53368, -32'sd949657, 32'sd731977, 32'sd734811, -32'sd561288, 32'sd280452, 32'sd949478, -32'sd728196, -32'sd1121608, -32'sd2610180, -32'sd2297936, -32'sd1404034, -32'sd1249814, 32'sd595403, 32'sd1663932, 32'sd304441, 32'sd1860173, 32'sd2530870, 32'sd948831, -32'sd306887, -32'sd1405231, -32'sd1965657, 32'sd842779, -32'sd2630540, 32'sd345078, 32'sd1874327, 32'sd1256725, -32'sd244317, 32'sd1811127, 32'sd128482, 32'sd670015, -32'sd398975, -32'sd1834832, 32'sd2026629, 32'sd728607, 32'sd1381032, -32'sd794527, -32'sd2034842, 32'sd562150, -32'sd1045285, -32'sd1541336, 32'sd221187, 32'sd950352, 32'sd2360753, 32'sd1610336, -32'sd1256720, -32'sd915375, -32'sd777408, -32'sd1200942, -32'sd2576193, -32'sd2153121, 32'sd707164, 32'sd1556349, 32'sd575610, 32'sd516138, -32'sd711941, -32'sd492566, -32'sd1737440, -32'sd597083, 32'sd0, 32'sd1377148, 32'sd2573600, 32'sd856243, 32'sd1073299, -32'sd2173286, -32'sd3026494, -32'sd504419, -32'sd929491, -32'sd1225080, 32'sd731789, 32'sd469696, -32'sd610125, 32'sd455220, -32'sd455874, -32'sd297529, -32'sd221786, -32'sd848898, -32'sd1186438, 32'sd779360, -32'sd844245, -32'sd840228, -32'sd1417183, -32'sd1569186, -32'sd1679758, 32'sd489703, 32'sd146795, 32'sd0, 32'sd0, 32'sd0, 32'sd12488, 32'sd1066650, 32'sd102182, -32'sd1582984, -32'sd1338335, -32'sd141131, 32'sd2397915, 32'sd5222, -32'sd1151061, 32'sd294981, 32'sd350245, 32'sd1806301, 32'sd2478678, -32'sd31743, -32'sd1284003, 32'sd471897, -32'sd1009105, -32'sd651656, -32'sd529915, -32'sd2807467, 32'sd982489, -32'sd363926, -32'sd80280, 32'sd47629, 32'sd1047607, 32'sd0, 32'sd0, 32'sd0, 32'sd652998, 32'sd144176, -32'sd396162, 32'sd588594, -32'sd201382, 32'sd2228528, -32'sd406708, -32'sd836639, -32'sd888822, 32'sd693908, 32'sd152788, 32'sd407611, -32'sd307912, 32'sd3107562, 32'sd2822389, 32'sd2694489, 32'sd1298991, 32'sd1424596, 32'sd95463, -32'sd616470, -32'sd1191785, -32'sd1791392, 32'sd704907, 32'sd52625, 32'sd291099, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2042074, -32'sd330577, -32'sd211858, -32'sd2148325, -32'sd439916, 32'sd301625, 32'sd538848, 32'sd781602, -32'sd519871, 32'sd1051648, 32'sd2009827, 32'sd2106058, 32'sd2105776, 32'sd820849, 32'sd2160250, -32'sd105272, 32'sd485026, -32'sd188779, -32'sd430446, -32'sd912097, 32'sd876997, -32'sd53760, 32'sd2146326, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1803321, 32'sd974381, 32'sd326047, 32'sd1530324, 32'sd1633456, 32'sd220727, 32'sd1194248, 32'sd63652, 32'sd1550028, 32'sd86564, 32'sd1478013, 32'sd2063539, -32'sd385379, 32'sd787406, 32'sd452529, -32'sd749655, 32'sd315463, 32'sd454620, -32'sd1376086, 32'sd2050930, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd30341, -32'sd931067, 32'sd529609, -32'sd105964, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1292844, -32'sd674988, -32'sd694146, -32'sd891479, 32'sd356108, 32'sd501077, 32'sd989150, 32'sd1604034, -32'sd613292, -32'sd767542, -32'sd566733, 32'sd1296726, 32'sd325630, 32'sd627670, 32'sd696309, 32'sd1104259, 32'sd1178816, 32'sd1088592, 32'sd1384690, 32'sd482484, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd920014, 32'sd1202062, 32'sd495549, 32'sd48640, -32'sd14586, 32'sd742623, 32'sd893370, -32'sd1646541, 32'sd37319, -32'sd22821, -32'sd1852518, -32'sd1315348, -32'sd1703829, -32'sd3557754, -32'sd822933, -32'sd1976246, -32'sd2409915, -32'sd383993, 32'sd31668, -32'sd136892, 32'sd891440, -32'sd470814, 32'sd385861, 32'sd1024845, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd99593, 32'sd1006339, -32'sd780658, -32'sd1202856, 32'sd1263040, -32'sd692515, -32'sd349555, 32'sd1643169, -32'sd1502966, -32'sd865866, -32'sd3000953, -32'sd2024293, -32'sd2252804, -32'sd32379, 32'sd351693, 32'sd1183232, -32'sd213537, -32'sd3038960, -32'sd1381715, -32'sd2365195, -32'sd334694, 32'sd167077, -32'sd1403983, -32'sd1745236, 32'sd487167, 32'sd0, 32'sd0, 32'sd324604, -32'sd283010, 32'sd858778, 32'sd239785, 32'sd512756, 32'sd340287, -32'sd2632336, -32'sd2819284, -32'sd2288746, -32'sd4534306, -32'sd2628634, -32'sd3723537, -32'sd1940067, 32'sd385945, 32'sd237592, 32'sd1052833, -32'sd520976, -32'sd290938, -32'sd420205, -32'sd1840283, 32'sd188594, -32'sd468581, -32'sd95534, -32'sd1151264, -32'sd814027, -32'sd1623811, 32'sd594918, 32'sd0, 32'sd941158, 32'sd1353136, -32'sd907765, -32'sd1488101, -32'sd1557432, 32'sd507757, -32'sd1757748, -32'sd1320698, 32'sd1297612, -32'sd642459, -32'sd1651992, -32'sd2566067, 32'sd148469, 32'sd625893, -32'sd143402, -32'sd646, -32'sd1194771, -32'sd2413044, -32'sd4350475, -32'sd2583786, -32'sd21272, 32'sd667345, -32'sd2654043, -32'sd114679, -32'sd1750439, 32'sd1792773, 32'sd50975, 32'sd0, 32'sd880821, -32'sd337714, 32'sd478038, -32'sd586160, 32'sd697013, 32'sd164881, -32'sd882850, -32'sd2308128, -32'sd1178611, -32'sd206723, -32'sd2288713, -32'sd508233, -32'sd1065045, 32'sd543761, 32'sd393387, -32'sd1142349, -32'sd1238503, -32'sd1949245, -32'sd1116365, -32'sd1079259, 32'sd243914, 32'sd479708, -32'sd533482, -32'sd946623, 32'sd77441, 32'sd1170601, -32'sd80241, 32'sd488562, 32'sd62890, -32'sd1100997, -32'sd1176443, -32'sd453436, -32'sd1302046, 32'sd917560, -32'sd2872382, -32'sd868458, 32'sd2479064, -32'sd1240472, -32'sd1397602, -32'sd3043160, -32'sd1939522, -32'sd603721, 32'sd956079, -32'sd1200263, -32'sd1187870, -32'sd441734, -32'sd1073146, -32'sd751463, 32'sd233673, 32'sd818505, 32'sd443069, -32'sd184246, 32'sd852349, 32'sd1585688, 32'sd1686559, 32'sd143673, 32'sd838755, 32'sd834148, -32'sd789142, 32'sd202314, 32'sd508494, 32'sd1643438, -32'sd1738392, -32'sd1131251, 32'sd582846, -32'sd1167181, -32'sd1611141, -32'sd266684, 32'sd699804, 32'sd1714201, 32'sd572902, 32'sd1080940, -32'sd1275166, 32'sd1132289, 32'sd216919, 32'sd390701, 32'sd238919, 32'sd1457385, 32'sd440573, 32'sd1637702, 32'sd831158, 32'sd1631479, -32'sd708121, 32'sd190888, -32'sd253678, -32'sd521946, 32'sd1772514, -32'sd790842, -32'sd868779, 32'sd866119, 32'sd1535671, -32'sd108885, -32'sd1329950, 32'sd46587, 32'sd834354, 32'sd133128, -32'sd806150, 32'sd1559543, 32'sd1276369, 32'sd1571912, -32'sd2379979, -32'sd875037, 32'sd1867519, 32'sd1380170, 32'sd305676, -32'sd875508, 32'sd1275359, 32'sd2712781, -32'sd195995, 32'sd1914440, -32'sd147374, 32'sd230875, 32'sd639534, 32'sd76012, 32'sd2617141, 32'sd1849237, -32'sd163777, 32'sd1034732, 32'sd1703262, 32'sd1300308, 32'sd1844820, 32'sd1517314, -32'sd644601, 32'sd1981680, -32'sd508431, 32'sd1162044, 32'sd638267, 32'sd68322, 32'sd1398565, -32'sd295488, -32'sd39707, 32'sd1617025, 32'sd1145314, -32'sd194880, 32'sd1018849, 32'sd349599, 32'sd1656790, -32'sd594606, 32'sd839579, 32'sd43154, 32'sd2224643, 32'sd1168882, -32'sd1048669, -32'sd859718, 32'sd1751660, -32'sd129647, 32'sd125172, 32'sd329197, 32'sd2340309, 32'sd3073341, 32'sd2272135, 32'sd1501568, -32'sd1118124, -32'sd660085, 32'sd1571955, 32'sd1827962, 32'sd1436306, -32'sd1692542, -32'sd927763, -32'sd150678, -32'sd55984, -32'sd1595506, 32'sd354428, 32'sd116272, -32'sd371748, -32'sd1545322, -32'sd1152325, 32'sd680584, 32'sd443191, -32'sd49894, 32'sd325777, -32'sd3888057, -32'sd2623317, 32'sd724252, -32'sd118777, -32'sd1303759, 32'sd2327694, 32'sd613570, 32'sd640540, 32'sd1499956, 32'sd1602579, -32'sd322637, 32'sd708075, 32'sd1172134, 32'sd153143, 32'sd382057, -32'sd1037946, 32'sd422975, -32'sd99472, -32'sd1183220, 32'sd509418, 32'sd1015209, -32'sd1087063, -32'sd214776, -32'sd356762, 32'sd560057, 32'sd651462, 32'sd726899, -32'sd109179, -32'sd3783732, -32'sd198049, -32'sd1481246, -32'sd1288975, 32'sd1011513, 32'sd1965579, 32'sd137097, 32'sd2464237, 32'sd1822821, -32'sd704347, -32'sd1085219, 32'sd897599, 32'sd136650, -32'sd68685, -32'sd1462646, -32'sd503175, -32'sd416018, -32'sd766652, -32'sd568845, 32'sd429897, -32'sd245609, -32'sd566175, -32'sd2182906, 32'sd181974, 32'sd1848705, -32'sd739139, -32'sd84406, -32'sd1360875, -32'sd1646778, 32'sd564604, 32'sd910407, 32'sd1896844, 32'sd669274, 32'sd1517536, 32'sd2225451, 32'sd2774364, 32'sd1313243, 32'sd558348, -32'sd385516, -32'sd1523290, -32'sd1048161, 32'sd493373, -32'sd641949, 32'sd896188, -32'sd1923191, -32'sd1271427, 32'sd857191, 32'sd503547, 32'sd1685146, -32'sd3211583, -32'sd1497447, -32'sd1088064, 32'sd1385657, -32'sd1125994, -32'sd896112, -32'sd141259, -32'sd342964, 32'sd830096, 32'sd284370, 32'sd3650137, 32'sd1209540, 32'sd1294445, 32'sd1548907, 32'sd705576, 32'sd2139122, -32'sd2775085, -32'sd1574573, -32'sd584765, 32'sd260373, -32'sd1734067, -32'sd485660, -32'sd343459, -32'sd1369504, -32'sd596089, -32'sd376969, 32'sd2162299, 32'sd3791537, -32'sd1280455, -32'sd1736298, 32'sd141432, 32'sd272228, 32'sd81786, -32'sd141956, -32'sd956630, -32'sd1038563, 32'sd530143, 32'sd2159307, 32'sd1076370, 32'sd4641249, 32'sd2320055, 32'sd2845780, -32'sd178474, -32'sd620091, -32'sd2676377, -32'sd3600931, -32'sd702256, -32'sd1609383, -32'sd561314, -32'sd631934, 32'sd1516407, 32'sd138727, 32'sd259389, 32'sd343899, 32'sd2133361, 32'sd3022336, -32'sd1113184, -32'sd3607269, 32'sd1373251, 32'sd0, 32'sd538589, -32'sd198368, -32'sd1056611, 32'sd395394, 32'sd1532316, 32'sd1418709, -32'sd884228, 32'sd2806845, 32'sd3067446, 32'sd2219235, 32'sd1149202, -32'sd1993231, -32'sd1916180, -32'sd2139744, -32'sd40869, 32'sd1438490, 32'sd1220132, 32'sd172937, -32'sd122350, 32'sd2244025, 32'sd1474084, 32'sd932673, 32'sd1320137, 32'sd70464, -32'sd190439, -32'sd952999, -32'sd530124, -32'sd835896, 32'sd37053, 32'sd931621, -32'sd503085, 32'sd2203839, 32'sd718959, -32'sd1279446, 32'sd97451, 32'sd3336831, 32'sd2959619, 32'sd791523, -32'sd1775217, -32'sd1031507, -32'sd1375574, 32'sd479668, -32'sd840305, 32'sd849226, -32'sd608698, -32'sd1296411, -32'sd1558707, 32'sd1911165, 32'sd8661, -32'sd1290520, -32'sd874114, 32'sd1101179, 32'sd928209, -32'sd1181957, 32'sd900161, 32'sd772369, 32'sd309587, -32'sd933983, 32'sd1143852, 32'sd267676, 32'sd254526, -32'sd732053, -32'sd1784076, 32'sd2835669, 32'sd2656219, 32'sd921669, -32'sd3487268, -32'sd2581886, -32'sd760328, -32'sd681340, -32'sd1913871, 32'sd579816, -32'sd371561, -32'sd1299641, -32'sd1572261, -32'sd548611, -32'sd1318357, -32'sd3424720, -32'sd1508488, 32'sd1882782, -32'sd68427, -32'sd1440943, 32'sd1392712, 32'sd0, 32'sd226172, -32'sd901869, 32'sd198026, 32'sd110307, -32'sd419682, 32'sd237791, -32'sd1841045, -32'sd136184, -32'sd471590, -32'sd1256142, 32'sd473264, -32'sd1173760, -32'sd1261797, -32'sd1244412, -32'sd1195815, -32'sd1307835, -32'sd177454, -32'sd2067258, -32'sd1053506, -32'sd504197, -32'sd3021975, -32'sd2917700, -32'sd1493331, -32'sd1671270, 32'sd424762, -32'sd1172279, 32'sd543916, 32'sd780037, 32'sd1634539, -32'sd1637717, 32'sd1867667, -32'sd646307, 32'sd748195, -32'sd972430, -32'sd879949, -32'sd193300, -32'sd45622, 32'sd378099, 32'sd242282, -32'sd2585878, -32'sd3153810, -32'sd3768055, -32'sd1075143, -32'sd273233, -32'sd1093841, -32'sd1682017, -32'sd285939, 32'sd242721, 32'sd895052, -32'sd549127, -32'sd1383511, -32'sd1893383, -32'sd1632102, 32'sd530072, 32'sd79906, 32'sd814907, 32'sd1114884, 32'sd431083, -32'sd793425, -32'sd2229303, -32'sd199869, 32'sd258742, 32'sd1076836, 32'sd605011, 32'sd951431, 32'sd397540, -32'sd86071, -32'sd153187, -32'sd1179911, -32'sd417587, -32'sd1038004, 32'sd735104, -32'sd1380836, -32'sd1986101, -32'sd1032208, 32'sd261532, 32'sd465196, -32'sd292694, -32'sd596789, -32'sd405115, -32'sd2087591, 32'sd304391, 32'sd605871, 32'sd0, 32'sd377299, -32'sd130250, -32'sd1304301, -32'sd944078, 32'sd839675, 32'sd649523, -32'sd973048, -32'sd227979, -32'sd639809, 32'sd1506013, -32'sd932117, -32'sd54177, -32'sd1980803, -32'sd1227708, 32'sd711881, -32'sd395101, -32'sd1385614, -32'sd1137946, 32'sd739916, 32'sd1176530, 32'sd342215, -32'sd132561, -32'sd1072421, -32'sd35153, -32'sd976918, 32'sd403107, 32'sd0, 32'sd0, 32'sd0, -32'sd346314, 32'sd224180, 32'sd1246476, 32'sd640616, -32'sd1374482, -32'sd821102, 32'sd918639, 32'sd1488126, 32'sd1129016, 32'sd147363, -32'sd274679, 32'sd1274995, 32'sd176065, -32'sd1464538, -32'sd153721, -32'sd1503789, 32'sd857757, 32'sd827325, -32'sd713553, 32'sd360824, -32'sd1130524, -32'sd998278, 32'sd188502, 32'sd1389897, 32'sd73967, 32'sd0, 32'sd0, 32'sd0, 32'sd718727, -32'sd1011981, -32'sd1256529, -32'sd522284, -32'sd1781820, -32'sd1011130, -32'sd539553, 32'sd1781350, -32'sd2737950, -32'sd392966, 32'sd412127, -32'sd1917894, -32'sd945347, -32'sd447946, -32'sd2340240, -32'sd1955456, -32'sd347395, -32'sd1305036, 32'sd459577, -32'sd183612, -32'sd2270262, 32'sd720975, 32'sd1118893, 32'sd504288, 32'sd273637, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1074700, 32'sd95293, -32'sd1200287, -32'sd1789786, -32'sd1155671, -32'sd2536900, -32'sd1176278, -32'sd430295, -32'sd913751, 32'sd904701, -32'sd1060872, -32'sd2882574, -32'sd2469142, 32'sd218138, 32'sd131867, -32'sd235831, 32'sd272826, -32'sd1494246, -32'sd2247602, -32'sd423890, -32'sd1044754, -32'sd184439, 32'sd347121, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1334966, 32'sd76858, 32'sd57916, 32'sd1350575, -32'sd10316, -32'sd46641, -32'sd90594, -32'sd1188445, 32'sd1097484, 32'sd488802, -32'sd2429976, -32'sd2409197, -32'sd2276089, -32'sd405960, 32'sd14350, -32'sd293178, -32'sd627579, 32'sd771314, -32'sd146530, 32'sd115664, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2491894, 32'sd2529544, -32'sd256008, 32'sd694465, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2127609, 32'sd390924, 32'sd181904, 32'sd880974, -32'sd54219, 32'sd1638064, 32'sd1193079, -32'sd843071, -32'sd88167, 32'sd2894056, 32'sd30031, 32'sd2227288, 32'sd741254, 32'sd1161915, -32'sd451651, 32'sd1087642, 32'sd1060125, 32'sd556392, -32'sd666326, 32'sd710480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd870099, 32'sd1629224, 32'sd910437, -32'sd763474, -32'sd1345440, 32'sd715091, 32'sd2466946, 32'sd2460611, 32'sd268895, 32'sd2434415, 32'sd1496735, -32'sd489186, 32'sd896176, 32'sd2230428, 32'sd495475, 32'sd1666891, 32'sd1265300, -32'sd1127138, 32'sd54427, 32'sd838511, -32'sd1604207, -32'sd1501054, 32'sd648141, 32'sd2198081, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd224689, 32'sd413293, 32'sd80900, 32'sd1029787, -32'sd211831, 32'sd1837973, 32'sd2423526, 32'sd2017513, -32'sd975556, 32'sd2228181, 32'sd885238, 32'sd2368399, 32'sd1097583, 32'sd1667639, 32'sd718894, -32'sd1465713, 32'sd479257, 32'sd1707283, 32'sd549349, 32'sd940564, -32'sd94435, 32'sd493992, 32'sd587836, -32'sd144285, 32'sd1872388, 32'sd0, 32'sd0, 32'sd518314, 32'sd737474, 32'sd469692, 32'sd1136998, -32'sd379571, -32'sd351224, 32'sd467051, 32'sd1776281, 32'sd1221838, -32'sd294770, 32'sd43365, 32'sd2863049, 32'sd2806997, 32'sd909228, 32'sd1913889, -32'sd1810297, -32'sd725990, -32'sd1330230, -32'sd1665830, -32'sd591347, -32'sd71782, -32'sd1834458, 32'sd239955, -32'sd33648, 32'sd871590, 32'sd490000, 32'sd1477745, 32'sd0, 32'sd1289846, 32'sd847044, 32'sd663105, -32'sd96232, -32'sd710187, 32'sd2323696, -32'sd203227, -32'sd322727, -32'sd2500420, -32'sd2389100, -32'sd668093, 32'sd884827, 32'sd364615, 32'sd283633, 32'sd1119954, -32'sd1121311, -32'sd314414, -32'sd1633726, -32'sd536915, -32'sd1043637, -32'sd667231, -32'sd1753411, -32'sd1604955, -32'sd400779, 32'sd91644, 32'sd989019, 32'sd301419, 32'sd0, 32'sd696395, 32'sd494375, -32'sd847109, -32'sd1897154, -32'sd1611528, -32'sd346825, 32'sd284212, -32'sd389410, -32'sd696291, 32'sd29334, 32'sd262341, 32'sd1287386, 32'sd2116119, 32'sd2010960, 32'sd1088533, -32'sd1409761, -32'sd923485, -32'sd1867252, -32'sd2027500, -32'sd2893807, -32'sd655721, -32'sd3381826, -32'sd1329320, 32'sd125441, -32'sd162900, 32'sd2215412, -32'sd825268, 32'sd653784, -32'sd497238, 32'sd60739, -32'sd355611, -32'sd1094549, -32'sd2164055, -32'sd2333488, 32'sd837079, 32'sd966427, -32'sd1506708, -32'sd379816, 32'sd2093401, 32'sd2309481, 32'sd3402664, 32'sd1685142, 32'sd1154085, -32'sd2286646, -32'sd3937215, -32'sd506462, -32'sd2557668, -32'sd2411888, -32'sd3269170, 32'sd171390, -32'sd1125709, 32'sd463171, 32'sd1669197, 32'sd321106, 32'sd939094, 32'sd525662, 32'sd1212984, 32'sd534205, -32'sd1879633, -32'sd654152, -32'sd953377, -32'sd1111482, -32'sd565554, -32'sd317836, -32'sd86538, 32'sd1778919, 32'sd574626, 32'sd31408, 32'sd2925973, 32'sd42985, -32'sd2343525, -32'sd3180202, -32'sd656553, -32'sd321364, -32'sd2227753, -32'sd2056936, -32'sd2096837, -32'sd883470, -32'sd2520632, -32'sd1311655, 32'sd1219804, 32'sd2091766, 32'sd276528, 32'sd11451, 32'sd860188, 32'sd1001926, 32'sd1057114, 32'sd79868, 32'sd174699, -32'sd400764, 32'sd1826096, 32'sd1018789, 32'sd2223857, -32'sd13435, 32'sd668525, -32'sd1331045, 32'sd806154, 32'sd249269, -32'sd1975733, -32'sd601921, 32'sd387348, 32'sd489504, 32'sd455267, -32'sd489844, -32'sd1104367, -32'sd20847, -32'sd517374, 32'sd1313937, 32'sd254730, 32'sd1474256, -32'sd374161, -32'sd688376, -32'sd330777, 32'sd139768, -32'sd765889, 32'sd1266542, -32'sd398374, 32'sd399237, 32'sd607968, -32'sd255755, -32'sd1716062, -32'sd87620, -32'sd471170, -32'sd322015, 32'sd1296032, -32'sd771824, -32'sd2518101, 32'sd335558, 32'sd800700, -32'sd327417, 32'sd641328, -32'sd636638, -32'sd1677841, 32'sd1049960, 32'sd116176, -32'sd1710917, 32'sd542531, 32'sd2069658, 32'sd470500, 32'sd1245688, -32'sd335071, -32'sd4018, 32'sd1249673, -32'sd375671, 32'sd386722, 32'sd482486, 32'sd432040, -32'sd207753, -32'sd297229, -32'sd614034, 32'sd373254, -32'sd722960, 32'sd1356702, 32'sd810600, -32'sd1918616, 32'sd448597, 32'sd34967, 32'sd1301091, 32'sd1958880, 32'sd1529875, -32'sd43507, -32'sd856490, -32'sd1787800, -32'sd885239, 32'sd759937, 32'sd799515, 32'sd960439, 32'sd384825, 32'sd339837, -32'sd155397, -32'sd1673205, 32'sd1900849, 32'sd458230, -32'sd189764, 32'sd44118, -32'sd843074, -32'sd347632, -32'sd1476163, -32'sd974226, -32'sd1784969, -32'sd1442706, 32'sd964710, -32'sd991250, 32'sd1121744, 32'sd1571284, 32'sd2085115, 32'sd2019147, 32'sd976820, 32'sd139733, -32'sd1308911, 32'sd357705, 32'sd2764062, 32'sd1568822, -32'sd1477323, -32'sd94687, 32'sd143045, -32'sd318616, 32'sd689552, -32'sd1173977, -32'sd1322096, -32'sd39389, 32'sd183333, -32'sd608678, -32'sd1338547, -32'sd82527, -32'sd255763, -32'sd1486262, -32'sd3008741, -32'sd2863664, 32'sd373080, 32'sd1166573, 32'sd1922363, 32'sd1547656, -32'sd359590, 32'sd1181149, -32'sd172938, 32'sd964753, -32'sd734776, 32'sd481581, 32'sd970033, -32'sd107150, -32'sd156741, 32'sd798983, 32'sd286312, -32'sd731440, 32'sd742736, -32'sd1502669, -32'sd3184652, -32'sd393632, -32'sd1003875, 32'sd1148091, 32'sd543988, 32'sd152728, -32'sd1645906, -32'sd2024740, -32'sd1458811, -32'sd1241560, -32'sd349709, 32'sd1533007, 32'sd2131611, 32'sd170789, -32'sd167309, -32'sd1927645, -32'sd810512, -32'sd1124835, 32'sd1523871, 32'sd618524, -32'sd634767, -32'sd594194, -32'sd93774, 32'sd1391800, 32'sd352162, 32'sd60830, -32'sd537081, -32'sd1079671, -32'sd1971182, -32'sd300325, 32'sd637470, 32'sd836496, 32'sd288193, -32'sd2011941, -32'sd2427513, -32'sd431257, -32'sd947335, -32'sd493798, 32'sd2213973, 32'sd1227584, 32'sd327984, 32'sd295003, 32'sd474369, -32'sd106022, 32'sd414738, 32'sd238430, 32'sd397120, 32'sd916873, 32'sd600751, -32'sd1181842, 32'sd944762, 32'sd211992, 32'sd557818, 32'sd551134, 32'sd506706, -32'sd155477, -32'sd365537, -32'sd863071, -32'sd1264355, 32'sd634365, -32'sd258551, -32'sd2543659, -32'sd3154574, -32'sd1150212, -32'sd1084737, 32'sd1594777, 32'sd1918926, 32'sd1264163, 32'sd79468, 32'sd1169725, -32'sd935991, -32'sd2406346, -32'sd339562, -32'sd875507, -32'sd411647, -32'sd241871, 32'sd1347577, 32'sd1060092, 32'sd362219, 32'sd890545, 32'sd0, 32'sd486950, -32'sd976267, 32'sd1137382, 32'sd1801465, -32'sd36982, -32'sd210005, -32'sd931228, -32'sd2356219, -32'sd2641338, -32'sd1504669, -32'sd89694, -32'sd72819, 32'sd2507403, 32'sd369843, 32'sd1449632, -32'sd1019595, -32'sd87680, -32'sd1067591, -32'sd185189, -32'sd586974, -32'sd225539, 32'sd55903, 32'sd1770290, 32'sd1183865, 32'sd2220862, 32'sd957086, -32'sd1138480, 32'sd1574692, 32'sd1067192, -32'sd363748, -32'sd636276, -32'sd3851, -32'sd1624425, 32'sd53344, -32'sd1198059, -32'sd2217090, -32'sd1714886, -32'sd1798816, -32'sd1077213, 32'sd1237178, 32'sd566837, 32'sd836416, 32'sd1485042, -32'sd711365, -32'sd313608, 32'sd451816, -32'sd278261, -32'sd1358593, -32'sd708937, 32'sd242001, -32'sd1773418, 32'sd1682290, 32'sd1989099, -32'sd1495392, 32'sd220005, 32'sd707149, 32'sd1072416, -32'sd521526, -32'sd2846974, 32'sd1567341, -32'sd644877, -32'sd664092, 32'sd124751, -32'sd4665, -32'sd1271862, -32'sd120277, -32'sd83038, 32'sd2169663, -32'sd1682966, -32'sd35222, 32'sd120914, 32'sd574909, 32'sd542825, 32'sd329439, -32'sd42297, 32'sd1297327, 32'sd1440815, -32'sd1245624, -32'sd1498617, 32'sd44734, -32'sd189058, 32'sd438984, -32'sd713365, 32'sd0, 32'sd747301, -32'sd1434033, 32'sd349160, -32'sd511522, -32'sd2229128, -32'sd129000, -32'sd1626729, -32'sd1021679, -32'sd442688, 32'sd2610078, 32'sd1141376, 32'sd1938325, 32'sd251323, 32'sd3664872, 32'sd2539635, 32'sd2084469, 32'sd835461, 32'sd2515088, -32'sd251729, 32'sd1946138, 32'sd1121928, -32'sd895758, -32'sd615212, 32'sd1651484, 32'sd169773, -32'sd479163, 32'sd755611, 32'sd632332, -32'sd450724, -32'sd20326, 32'sd142013, 32'sd1688701, 32'sd1034771, -32'sd1197888, -32'sd1621119, -32'sd636873, -32'sd627957, 32'sd727742, 32'sd576764, -32'sd595523, 32'sd1303323, 32'sd1619401, 32'sd3402025, 32'sd1728097, 32'sd2494464, 32'sd2174625, 32'sd994685, 32'sd423772, -32'sd681827, -32'sd2761815, 32'sd1308750, 32'sd2656651, -32'sd426892, 32'sd1355990, -32'sd54290, 32'sd1489796, 32'sd400919, -32'sd734618, 32'sd491084, 32'sd1847495, 32'sd1230606, 32'sd593385, -32'sd592053, -32'sd1929498, 32'sd404430, -32'sd1919152, -32'sd844108, -32'sd71672, -32'sd426118, -32'sd675437, 32'sd822364, -32'sd255314, -32'sd324248, 32'sd976089, -32'sd613967, 32'sd346426, 32'sd12931, -32'sd1080090, -32'sd1285900, -32'sd1011939, 32'sd657499, 32'sd806350, 32'sd765581, 32'sd0, -32'sd286472, 32'sd13296, -32'sd911932, 32'sd1095706, 32'sd829801, 32'sd1108180, 32'sd394573, -32'sd57987, -32'sd1690100, -32'sd791560, -32'sd507869, -32'sd1389875, -32'sd487459, -32'sd1190365, 32'sd1302012, 32'sd1548797, 32'sd1650188, 32'sd563896, -32'sd482363, 32'sd1266327, 32'sd473110, -32'sd429724, 32'sd680500, 32'sd523607, -32'sd1022026, -32'sd291547, 32'sd0, 32'sd0, 32'sd0, 32'sd569091, -32'sd114868, -32'sd908812, -32'sd641765, 32'sd472080, 32'sd87072, -32'sd201946, 32'sd534312, 32'sd788698, 32'sd845832, -32'sd461848, -32'sd265611, 32'sd1073102, -32'sd4137, 32'sd1627190, 32'sd633333, 32'sd542534, 32'sd1306802, 32'sd499098, 32'sd1101823, 32'sd869371, 32'sd1779292, -32'sd45324, 32'sd116304, 32'sd238215, 32'sd0, 32'sd0, 32'sd0, -32'sd1379018, 32'sd1522292, -32'sd883086, -32'sd869258, -32'sd336056, 32'sd634426, -32'sd185979, -32'sd436332, -32'sd979236, -32'sd774775, 32'sd164538, -32'sd662517, -32'sd246098, 32'sd545368, -32'sd1478309, -32'sd75429, -32'sd682273, 32'sd162512, -32'sd1073192, 32'sd798131, 32'sd1473816, 32'sd537444, -32'sd801447, 32'sd332545, 32'sd1671776, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd204205, 32'sd229332, 32'sd744263, -32'sd2119281, -32'sd393272, 32'sd241687, -32'sd2521157, -32'sd477346, -32'sd11910, -32'sd736905, -32'sd3133770, 32'sd241376, -32'sd181952, 32'sd1354891, 32'sd1982022, 32'sd2352944, -32'sd951382, -32'sd713007, -32'sd32646, 32'sd1329894, 32'sd1346918, 32'sd36254, 32'sd170964, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd743870, 32'sd182918, 32'sd154338, 32'sd212758, -32'sd748952, -32'sd261443, -32'sd1032485, -32'sd393321, -32'sd1301807, 32'sd985663, 32'sd2021184, 32'sd268986, 32'sd1277516, -32'sd1235059, -32'sd1013172, -32'sd204042, -32'sd1157505, 32'sd294886, -32'sd1508416, 32'sd1058716, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd181347, -32'sd494376, 32'sd1407663, 32'sd1878049, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd473803, 32'sd302194, -32'sd1608793, 32'sd561262, -32'sd1599312, -32'sd86091, -32'sd204784, -32'sd236457, -32'sd525992, 32'sd1723779, 32'sd1164078, 32'sd967808, -32'sd525662, 32'sd190152, -32'sd571272, -32'sd879478, 32'sd410563, -32'sd126694, 32'sd710492, 32'sd932267, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1746754, 32'sd235448, -32'sd379622, -32'sd749653, 32'sd897679, 32'sd61788, 32'sd296284, 32'sd96658, 32'sd2129261, 32'sd673815, 32'sd1957984, 32'sd2965215, 32'sd1442071, 32'sd1327454, -32'sd975993, 32'sd606670, -32'sd966747, -32'sd409080, -32'sd96573, 32'sd939097, -32'sd369776, 32'sd2493631, 32'sd974838, 32'sd1587741, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1045757, -32'sd150556, -32'sd163999, 32'sd1415052, 32'sd9999, 32'sd1437088, -32'sd420507, 32'sd1412279, 32'sd2429985, 32'sd2955936, 32'sd4650186, 32'sd3396427, 32'sd3004346, 32'sd1063281, 32'sd3214884, 32'sd2009204, 32'sd3320625, 32'sd1368180, -32'sd444636, -32'sd1862386, 32'sd354307, -32'sd2045574, 32'sd1108893, 32'sd133350, -32'sd1500189, 32'sd0, 32'sd0, 32'sd655249, 32'sd760765, 32'sd304605, -32'sd432884, 32'sd590082, -32'sd459832, -32'sd451986, -32'sd813980, -32'sd1036439, 32'sd3928467, 32'sd2462286, 32'sd1319703, 32'sd2017242, 32'sd3457344, 32'sd2297255, 32'sd3084144, 32'sd1637465, 32'sd1261539, 32'sd1258936, -32'sd239625, -32'sd1025820, -32'sd1635013, -32'sd2203574, 32'sd327600, 32'sd554164, -32'sd813718, 32'sd243835, 32'sd0, 32'sd2099946, -32'sd1045409, 32'sd204153, -32'sd1012945, 32'sd315524, -32'sd723309, -32'sd161731, -32'sd2414000, -32'sd2052342, 32'sd885016, -32'sd1290104, 32'sd888239, 32'sd765503, 32'sd968949, 32'sd2600975, 32'sd1525833, 32'sd565248, 32'sd2776031, 32'sd1836301, 32'sd816068, -32'sd239271, 32'sd1418346, 32'sd855500, 32'sd646954, 32'sd577158, -32'sd1570601, -32'sd548642, 32'sd0, 32'sd1384322, -32'sd558969, 32'sd1334527, -32'sd2267170, -32'sd12726, -32'sd648859, 32'sd150404, -32'sd1074288, -32'sd323691, -32'sd201229, -32'sd1487075, -32'sd1718377, 32'sd2176921, 32'sd517224, -32'sd123309, 32'sd1532121, 32'sd643565, 32'sd1220890, 32'sd788431, -32'sd229543, -32'sd586043, 32'sd116542, -32'sd360961, 32'sd996334, -32'sd1686091, 32'sd292165, 32'sd822818, 32'sd1487776, 32'sd1288178, 32'sd807926, 32'sd1419425, -32'sd396886, -32'sd1104913, 32'sd408673, -32'sd2142724, -32'sd2044274, -32'sd938489, -32'sd2146199, -32'sd562396, -32'sd1597895, -32'sd1093253, 32'sd521092, 32'sd1599645, 32'sd785684, 32'sd1937838, 32'sd2335917, 32'sd699432, 32'sd575789, 32'sd741630, 32'sd1475209, 32'sd1140395, 32'sd535440, -32'sd904551, 32'sd176113, 32'sd856757, 32'sd573125, 32'sd604484, -32'sd148052, -32'sd1068578, -32'sd465339, -32'sd2173165, -32'sd1342365, -32'sd1377332, -32'sd495358, 32'sd1696623, -32'sd80543, -32'sd2750540, -32'sd2024769, -32'sd2714550, -32'sd1375327, -32'sd1536709, 32'sd775249, 32'sd2125679, 32'sd783018, 32'sd1549170, 32'sd776346, 32'sd674950, -32'sd93786, 32'sd282216, -32'sd2521516, 32'sd441738, 32'sd133224, 32'sd1039329, 32'sd250890, -32'sd699694, -32'sd721501, 32'sd1473513, -32'sd401410, -32'sd1746761, -32'sd1618954, -32'sd1472687, -32'sd2735904, -32'sd697979, -32'sd3270717, -32'sd5451040, -32'sd5395157, -32'sd4807829, -32'sd1498539, -32'sd1391432, 32'sd443789, 32'sd2007413, 32'sd882512, 32'sd1294275, 32'sd1276147, 32'sd1941884, -32'sd911845, 32'sd101462, -32'sd1082739, -32'sd498418, -32'sd197542, 32'sd93599, 32'sd908919, -32'sd1081498, 32'sd965147, 32'sd1059666, 32'sd541345, -32'sd24678, -32'sd1821839, -32'sd3732081, -32'sd4385595, -32'sd2783022, -32'sd3892306, -32'sd6705160, -32'sd3673083, -32'sd2976042, 32'sd953825, -32'sd843077, 32'sd631504, -32'sd371611, -32'sd61671, -32'sd291119, -32'sd104139, 32'sd880849, -32'sd662192, -32'sd612245, -32'sd1099342, 32'sd413913, -32'sd388568, -32'sd807834, -32'sd358112, 32'sd856288, 32'sd631803, -32'sd778416, -32'sd1193113, -32'sd3388046, -32'sd3176321, -32'sd3971356, -32'sd4346134, -32'sd2527580, -32'sd2725926, -32'sd4563636, -32'sd2789504, 32'sd814061, 32'sd2406937, 32'sd1571138, -32'sd3301118, -32'sd323148, -32'sd1399597, 32'sd461699, -32'sd245565, 32'sd75877, 32'sd1519427, -32'sd309019, -32'sd2880829, -32'sd340265, -32'sd1457537, 32'sd123119, 32'sd1237533, -32'sd1224808, -32'sd1635541, -32'sd1226395, -32'sd2949631, -32'sd1344229, -32'sd1900944, -32'sd2369263, -32'sd675306, -32'sd478609, -32'sd530210, 32'sd202201, 32'sd1846757, 32'sd1880298, 32'sd3001163, 32'sd1198510, -32'sd1716448, -32'sd1830827, -32'sd131083, -32'sd2656592, -32'sd2912818, 32'sd489462, -32'sd836185, -32'sd315159, -32'sd2602462, -32'sd1723272, -32'sd501555, 32'sd677774, 32'sd1077405, -32'sd714467, 32'sd309309, -32'sd411457, -32'sd445268, -32'sd1852654, -32'sd1597082, 32'sd600193, -32'sd37169, 32'sd2238301, 32'sd1991250, 32'sd3151845, 32'sd2273320, 32'sd2575795, 32'sd3441110, -32'sd232684, -32'sd1039208, -32'sd2403678, -32'sd172740, -32'sd2663735, -32'sd52785, 32'sd354000, 32'sd617586, 32'sd1849647, -32'sd679640, 32'sd58990, 32'sd258724, 32'sd1224052, 32'sd966373, -32'sd309488, 32'sd578114, 32'sd117051, 32'sd2684033, 32'sd2108433, 32'sd1385478, 32'sd1577133, 32'sd3261301, 32'sd2611403, 32'sd2577689, 32'sd672000, 32'sd1639756, -32'sd783123, 32'sd360201, -32'sd673562, -32'sd446343, 32'sd546118, 32'sd1913772, -32'sd213508, -32'sd1280820, -32'sd82293, -32'sd173090, 32'sd863983, 32'sd662938, 32'sd243054, -32'sd1402426, 32'sd1412806, -32'sd1153971, -32'sd2401, -32'sd733589, 32'sd1256954, 32'sd2262119, 32'sd1193268, 32'sd260104, 32'sd1712384, 32'sd1468267, 32'sd100967, 32'sd108482, 32'sd819791, -32'sd1965153, -32'sd3038193, -32'sd1703763, -32'sd1170797, -32'sd275790, 32'sd1258481, 32'sd472566, -32'sd693059, -32'sd2193183, 32'sd880267, 32'sd385647, -32'sd1312683, -32'sd1134423, -32'sd829000, 32'sd667585, 32'sd897529, 32'sd1270337, 32'sd1289764, 32'sd278663, -32'sd554647, 32'sd1221830, 32'sd1622282, -32'sd430682, 32'sd1383590, -32'sd343638, 32'sd731437, -32'sd331889, 32'sd261050, -32'sd482929, -32'sd2289632, -32'sd2846230, 32'sd844820, 32'sd539163, 32'sd3744700, 32'sd1234241, 32'sd1114441, -32'sd41615, 32'sd484819, 32'sd304763, -32'sd207209, -32'sd65742, 32'sd386924, 32'sd1502509, 32'sd1161046, 32'sd0, 32'sd53245, 32'sd1249101, 32'sd645365, 32'sd126038, -32'sd280409, 32'sd695268, 32'sd1137545, -32'sd430886, 32'sd560606, -32'sd783074, 32'sd467762, -32'sd3109425, -32'sd3638267, -32'sd1717469, 32'sd461476, 32'sd3982848, 32'sd2441728, 32'sd2618989, 32'sd1540819, 32'sd576083, 32'sd2267280, 32'sd319482, 32'sd369808, 32'sd1016738, 32'sd761763, 32'sd184230, 32'sd657630, 32'sd418016, 32'sd1313416, 32'sd1683748, 32'sd2094809, 32'sd601143, 32'sd1306045, 32'sd471686, 32'sd502754, 32'sd165152, 32'sd372523, -32'sd1022105, 32'sd508375, -32'sd3227104, -32'sd2031600, 32'sd259248, 32'sd1342414, 32'sd1780287, 32'sd2078226, 32'sd1373184, -32'sd830383, 32'sd284015, 32'sd675944, -32'sd108095, 32'sd386651, -32'sd932322, 32'sd1081064, -32'sd1253444, 32'sd188329, 32'sd1198383, -32'sd407316, -32'sd419946, -32'sd562161, -32'sd237858, 32'sd469339, 32'sd684048, 32'sd885583, 32'sd446771, -32'sd564401, -32'sd277320, -32'sd1907689, -32'sd313901, 32'sd771038, 32'sd375730, 32'sd3817663, 32'sd1624407, -32'sd368512, -32'sd298432, -32'sd1543267, -32'sd1489427, -32'sd439582, -32'sd328152, -32'sd1383192, -32'sd834135, -32'sd1888332, 32'sd1312649, 32'sd24850, 32'sd0, 32'sd896345, 32'sd1415579, 32'sd1195688, -32'sd967963, 32'sd282906, 32'sd2115864, 32'sd1206979, 32'sd651948, 32'sd796495, 32'sd1384176, 32'sd1177912, 32'sd2351097, 32'sd1006242, -32'sd297667, -32'sd1940381, 32'sd1566463, 32'sd761308, -32'sd1333839, -32'sd2430740, -32'sd1535108, -32'sd2030767, -32'sd568600, -32'sd1356003, -32'sd23947, -32'sd1279958, -32'sd609376, 32'sd747391, -32'sd264651, -32'sd582776, 32'sd168882, 32'sd1782961, 32'sd714799, -32'sd1295814, 32'sd1312951, 32'sd284677, 32'sd2253724, -32'sd963534, 32'sd214002, 32'sd900959, 32'sd1304014, -32'sd1065043, -32'sd1818058, -32'sd2281381, -32'sd1514861, -32'sd1025099, -32'sd1639785, -32'sd873455, -32'sd317398, -32'sd324757, 32'sd369110, 32'sd1715969, -32'sd2216212, 32'sd98377, 32'sd493215, 32'sd170982, -32'sd196754, 32'sd1058901, 32'sd1243140, -32'sd812104, -32'sd455301, -32'sd1434731, 32'sd1931927, 32'sd1954052, 32'sd26653, -32'sd1244354, -32'sd359621, 32'sd665, 32'sd647562, 32'sd1053447, -32'sd770168, -32'sd471736, -32'sd1235341, -32'sd906247, -32'sd519857, -32'sd196604, -32'sd634325, 32'sd1243031, 32'sd1356157, -32'sd1094666, 32'sd476569, -32'sd289734, -32'sd728398, 32'sd1196520, 32'sd0, 32'sd1103058, -32'sd985058, -32'sd387733, 32'sd882997, -32'sd609784, -32'sd680760, -32'sd408147, -32'sd1339550, 32'sd1025978, 32'sd1152649, 32'sd1963765, 32'sd2652435, 32'sd430436, 32'sd888816, -32'sd1327035, -32'sd1278522, -32'sd2530550, -32'sd3134790, -32'sd255041, 32'sd576367, -32'sd181477, 32'sd293214, -32'sd2031964, 32'sd931714, 32'sd1064558, 32'sd1043495, 32'sd0, 32'sd0, 32'sd0, -32'sd124934, 32'sd664894, 32'sd1453527, -32'sd452158, 32'sd246906, -32'sd106982, 32'sd2180937, 32'sd1046201, -32'sd1812506, -32'sd12733, -32'sd569870, -32'sd485107, 32'sd779394, 32'sd1169634, -32'sd2363804, -32'sd2739063, -32'sd1478188, -32'sd1010812, 32'sd1341762, -32'sd958745, 32'sd515461, 32'sd633158, 32'sd777473, -32'sd113014, 32'sd1298667, 32'sd0, 32'sd0, 32'sd0, 32'sd1519177, -32'sd1055051, 32'sd344427, 32'sd147351, -32'sd405160, -32'sd2418988, -32'sd646221, -32'sd1360997, -32'sd2293603, -32'sd559335, -32'sd1748938, -32'sd207097, 32'sd365597, -32'sd1078587, -32'sd196556, 32'sd312525, 32'sd217344, 32'sd1399960, 32'sd909502, -32'sd638097, -32'sd795059, -32'sd1879030, 32'sd160672, 32'sd613530, -32'sd903371, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1634328, 32'sd463606, 32'sd1155484, 32'sd469568, 32'sd18084, -32'sd996508, 32'sd187799, 32'sd1544874, -32'sd56158, 32'sd579965, 32'sd1388775, 32'sd2146649, 32'sd1538368, 32'sd526391, -32'sd447126, 32'sd1029036, -32'sd73609, 32'sd204617, -32'sd847266, -32'sd462292, -32'sd204707, 32'sd347864, 32'sd527045, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1210884, -32'sd361440, 32'sd1219613, -32'sd867777, 32'sd795888, -32'sd62166, 32'sd945714, 32'sd1204319, 32'sd916133, 32'sd1224638, 32'sd1471568, 32'sd1259709, 32'sd1441549, 32'sd2386233, 32'sd846986, 32'sd1208380, 32'sd479814, -32'sd218597, 32'sd1601323, 32'sd903377, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd69376, -32'sd5432, 32'sd24274, -32'sd571407, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd19348, -32'sd814302, -32'sd162259, 32'sd74001, 32'sd161348, -32'sd191819, -32'sd575520, 32'sd749102, -32'sd807787, 32'sd540588, -32'sd94539, 32'sd421614, 32'sd723444, 32'sd696186, -32'sd165641, 32'sd758011, -32'sd1251994, 32'sd503014, -32'sd135464, -32'sd440583, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd433715, -32'sd798218, -32'sd649010, -32'sd189214, -32'sd1286261, 32'sd749974, 32'sd1251770, -32'sd1354807, 32'sd79966, -32'sd69284, -32'sd149234, 32'sd1154763, -32'sd18590, -32'sd1689490, -32'sd1737453, -32'sd1049318, 32'sd290174, -32'sd293444, 32'sd390527, -32'sd1512723, 32'sd834137, -32'sd1256094, 32'sd386203, 32'sd356686, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd715547, -32'sd822801, 32'sd537298, -32'sd1375283, -32'sd1262572, -32'sd972227, 32'sd685816, -32'sd1020226, -32'sd1312958, -32'sd1304626, -32'sd897594, -32'sd621287, -32'sd1919228, -32'sd897254, -32'sd1175054, 32'sd334126, 32'sd747630, 32'sd390309, 32'sd460656, 32'sd1431018, -32'sd303855, -32'sd427468, 32'sd1444538, -32'sd268940, 32'sd902130, 32'sd0, 32'sd0, 32'sd294514, 32'sd114815, 32'sd65064, -32'sd1505178, -32'sd1346829, -32'sd1336497, -32'sd1766321, -32'sd2005055, -32'sd2562760, -32'sd2992856, -32'sd978701, -32'sd1365131, -32'sd1466562, -32'sd2697420, -32'sd1722352, -32'sd555379, 32'sd1177691, 32'sd3273372, 32'sd2837732, 32'sd548262, -32'sd204175, 32'sd936727, -32'sd1465515, 32'sd185009, -32'sd1632293, 32'sd1671972, 32'sd890281, 32'sd0, -32'sd548900, 32'sd1334277, -32'sd39247, -32'sd947295, -32'sd628184, -32'sd835580, -32'sd2102274, -32'sd1549901, -32'sd1418647, -32'sd1874186, -32'sd1111306, -32'sd1182614, -32'sd988647, -32'sd353163, -32'sd1131759, -32'sd1212368, -32'sd1596332, 32'sd1890092, 32'sd2470382, 32'sd1765882, -32'sd163280, 32'sd1330764, -32'sd472987, -32'sd190142, 32'sd1831940, 32'sd1099344, 32'sd459175, 32'sd0, -32'sd82026, -32'sd376725, -32'sd377699, 32'sd1070680, -32'sd944014, 32'sd846586, -32'sd893080, -32'sd2400834, -32'sd126929, -32'sd1557651, -32'sd396059, -32'sd1955385, -32'sd250755, 32'sd1676403, 32'sd182595, 32'sd308354, 32'sd372522, 32'sd330457, -32'sd1523733, -32'sd2356402, -32'sd1193822, -32'sd1521785, -32'sd87554, 32'sd63695, 32'sd469536, 32'sd684814, 32'sd719908, 32'sd332553, -32'sd1078235, 32'sd140151, -32'sd774580, -32'sd87016, -32'sd102505, -32'sd724291, -32'sd2099848, -32'sd1378688, -32'sd3331561, -32'sd1923467, -32'sd854839, 32'sd431785, 32'sd939877, 32'sd106586, 32'sd1731519, 32'sd51165, 32'sd678532, 32'sd672337, 32'sd78112, 32'sd1232610, -32'sd1188195, 32'sd1168587, 32'sd753032, -32'sd826305, 32'sd207131, 32'sd846473, 32'sd136024, -32'sd666695, 32'sd1038037, -32'sd422896, -32'sd1340387, -32'sd103605, -32'sd1196175, -32'sd1919415, -32'sd2061396, -32'sd1469041, -32'sd1185228, -32'sd1126508, -32'sd401846, 32'sd1769543, 32'sd269372, 32'sd209755, 32'sd12570, -32'sd278724, 32'sd723875, -32'sd202005, 32'sd2649975, 32'sd1200172, -32'sd258711, 32'sd991202, -32'sd2090246, 32'sd253438, -32'sd161283, 32'sd836844, 32'sd971548, -32'sd713518, -32'sd231224, -32'sd912954, -32'sd1420562, 32'sd1425216, -32'sd1408488, -32'sd535178, -32'sd2027432, -32'sd1036791, 32'sd1933558, 32'sd3351749, 32'sd291372, -32'sd297700, 32'sd751508, -32'sd3433242, -32'sd2256440, -32'sd301270, 32'sd3067831, 32'sd3013930, 32'sd2012489, 32'sd1208195, 32'sd2341087, -32'sd1182177, -32'sd1646460, -32'sd1446579, 32'sd531019, 32'sd310300, -32'sd235, -32'sd1034851, -32'sd149889, -32'sd2729829, -32'sd1108067, -32'sd7637, -32'sd1271360, -32'sd1734172, 32'sd595449, 32'sd2269486, 32'sd3087761, 32'sd859816, 32'sd600976, -32'sd300651, -32'sd2723697, -32'sd850312, -32'sd717321, 32'sd1280171, 32'sd1551790, 32'sd3132885, 32'sd2140005, 32'sd939034, -32'sd842983, -32'sd276858, -32'sd116664, -32'sd2555112, 32'sd634287, 32'sd1020919, 32'sd1459854, -32'sd113482, -32'sd1046568, -32'sd1967145, -32'sd1345269, -32'sd205914, -32'sd161330, 32'sd1194138, 32'sd805856, 32'sd1649486, 32'sd969745, -32'sd1268488, -32'sd3127483, -32'sd3272077, -32'sd2536828, -32'sd854799, 32'sd592460, 32'sd2564580, 32'sd2515381, 32'sd1879168, 32'sd2401064, 32'sd3080257, 32'sd1051681, -32'sd452254, -32'sd1810821, -32'sd1579521, 32'sd1063098, -32'sd201290, -32'sd10567, -32'sd593500, -32'sd7557, -32'sd877954, -32'sd837686, 32'sd1267379, 32'sd1367672, 32'sd1245282, 32'sd1103688, -32'sd161007, -32'sd875205, -32'sd3170856, -32'sd2090553, -32'sd1253908, 32'sd243425, 32'sd1935780, 32'sd3778716, 32'sd3284418, 32'sd3668564, 32'sd3268736, 32'sd3038831, 32'sd2706813, 32'sd371268, 32'sd436193, 32'sd205613, -32'sd2096769, 32'sd586637, 32'sd629559, -32'sd699752, 32'sd866812, -32'sd745542, 32'sd882671, -32'sd2116623, 32'sd198514, 32'sd404983, 32'sd1883250, -32'sd1279231, -32'sd526875, -32'sd3179227, -32'sd2329728, -32'sd1372626, -32'sd1159253, 32'sd1967214, 32'sd4905230, 32'sd3429067, 32'sd2346880, 32'sd2320461, 32'sd2838827, 32'sd1015008, -32'sd1125832, -32'sd55003, -32'sd668858, -32'sd2623679, -32'sd2529699, -32'sd1086636, 32'sd642982, -32'sd1050558, -32'sd674943, -32'sd450277, -32'sd1780882, -32'sd1843076, 32'sd603131, -32'sd1047875, -32'sd466836, -32'sd1797696, -32'sd746715, -32'sd1517354, -32'sd401367, 32'sd1324738, 32'sd2458494, 32'sd1919010, 32'sd3916833, 32'sd2715186, 32'sd1525459, 32'sd28120, 32'sd1379967, -32'sd804822, -32'sd2002934, -32'sd2654261, 32'sd308402, 32'sd1146412, -32'sd164058, 32'sd1322891, 32'sd91248, -32'sd427889, 32'sd893739, -32'sd685277, -32'sd1332953, -32'sd1466434, 32'sd766016, 32'sd127638, -32'sd405215, -32'sd165121, -32'sd343557, -32'sd1827327, -32'sd2154940, -32'sd618007, 32'sd1886003, 32'sd2353068, 32'sd1246434, 32'sd386168, 32'sd2004255, -32'sd529166, -32'sd2885514, -32'sd1347100, -32'sd1094931, -32'sd1674112, -32'sd512270, 32'sd188210, -32'sd145587, -32'sd1471875, -32'sd453569, 32'sd379578, 32'sd1142427, -32'sd1035744, 32'sd809380, 32'sd65330, -32'sd879951, -32'sd2364238, -32'sd524392, 32'sd1618513, 32'sd1418670, 32'sd1506166, 32'sd1179371, 32'sd3201825, 32'sd1392043, 32'sd3624141, 32'sd1828339, -32'sd907628, -32'sd762052, -32'sd1221821, -32'sd2832872, -32'sd1318069, -32'sd1901070, -32'sd817264, -32'sd1879997, 32'sd310446, 32'sd2026103, -32'sd276155, -32'sd1473907, -32'sd722296, 32'sd0, -32'sd1001046, 32'sd851258, -32'sd1672982, -32'sd2885750, -32'sd2686599, -32'sd1687333, 32'sd922593, 32'sd2214214, -32'sd7166, 32'sd1348992, 32'sd3539458, 32'sd2561767, 32'sd4469774, 32'sd276626, -32'sd3323634, -32'sd1258359, -32'sd1931753, -32'sd1720738, -32'sd817521, -32'sd467330, -32'sd2479779, -32'sd1439809, -32'sd9211, 32'sd581335, -32'sd933546, -32'sd855181, -32'sd787051, 32'sd100650, 32'sd534929, -32'sd416062, 32'sd1151682, -32'sd23562, -32'sd1324436, -32'sd1508038, 32'sd1271048, 32'sd581418, 32'sd79468, 32'sd1061278, 32'sd967565, -32'sd608663, -32'sd21384, 32'sd560258, -32'sd700386, -32'sd2270960, -32'sd357526, -32'sd1318243, -32'sd2081218, -32'sd565675, -32'sd1355833, -32'sd741360, 32'sd68150, -32'sd340992, 32'sd411348, -32'sd560852, -32'sd387023, 32'sd662760, -32'sd859318, -32'sd777922, 32'sd2053069, 32'sd112666, -32'sd82103, -32'sd98664, 32'sd1835274, 32'sd314842, -32'sd1733983, -32'sd3321529, -32'sd2425496, -32'sd2754568, -32'sd1218184, -32'sd284041, -32'sd556146, 32'sd2058274, 32'sd7661, 32'sd690105, -32'sd1714904, -32'sd1194369, -32'sd898149, 32'sd547927, -32'sd634407, -32'sd2196439, 32'sd144546, -32'sd1730561, 32'sd1848609, 32'sd0, -32'sd739144, 32'sd1107098, 32'sd615085, 32'sd1392158, -32'sd738144, -32'sd519726, 32'sd1004305, 32'sd235623, -32'sd1145403, -32'sd2699865, -32'sd1701749, -32'sd765913, -32'sd2030258, -32'sd1005672, 32'sd1789013, 32'sd560725, 32'sd405949, 32'sd882900, -32'sd1840436, -32'sd765791, -32'sd720768, 32'sd207402, -32'sd1369967, 32'sd1176642, -32'sd986930, -32'sd1641879, 32'sd82535, -32'sd71807, -32'sd1028790, 32'sd1648873, 32'sd899856, 32'sd619835, 32'sd1414184, 32'sd668016, 32'sd1115034, 32'sd1302775, 32'sd179508, 32'sd1093030, -32'sd2122589, -32'sd2165749, -32'sd1678558, -32'sd16034, -32'sd461239, 32'sd1709729, -32'sd770280, 32'sd293438, 32'sd65277, -32'sd74385, -32'sd1678090, 32'sd124417, 32'sd739902, -32'sd260335, -32'sd267772, -32'sd958215, -32'sd539638, -32'sd245802, -32'sd834292, -32'sd925163, -32'sd995578, 32'sd35516, 32'sd2267037, 32'sd1086643, 32'sd108054, 32'sd347004, 32'sd564640, -32'sd290073, -32'sd985418, -32'sd2216736, -32'sd1059486, -32'sd2660535, -32'sd1047710, -32'sd815130, -32'sd817374, -32'sd1083009, -32'sd2077312, -32'sd873416, -32'sd1542493, -32'sd1156146, 32'sd514883, -32'sd1846149, -32'sd973741, -32'sd238651, -32'sd271953, 32'sd0, -32'sd258988, -32'sd771371, -32'sd1571576, -32'sd289603, 32'sd1205430, -32'sd1214959, 32'sd749889, 32'sd1435395, 32'sd1065568, 32'sd156370, 32'sd1614621, -32'sd413989, -32'sd167625, -32'sd1708372, -32'sd1006586, -32'sd666390, -32'sd1536551, 32'sd1443813, -32'sd673, -32'sd1137199, -32'sd1533547, -32'sd189321, -32'sd214193, 32'sd1130819, -32'sd560283, 32'sd1539881, 32'sd0, 32'sd0, 32'sd0, 32'sd812532, -32'sd2307400, 32'sd1748665, -32'sd506243, -32'sd318612, 32'sd958604, -32'sd938150, -32'sd207405, -32'sd169410, -32'sd671330, -32'sd15440, -32'sd859220, 32'sd356558, -32'sd1218573, 32'sd414550, -32'sd497059, -32'sd70097, -32'sd1349336, -32'sd1455095, 32'sd200999, -32'sd236916, -32'sd406054, 32'sd1756204, -32'sd1019736, -32'sd689169, 32'sd0, 32'sd0, 32'sd0, -32'sd652905, -32'sd256410, 32'sd477399, 32'sd1952692, 32'sd492477, 32'sd1624603, 32'sd2545513, 32'sd624120, 32'sd1062110, 32'sd690623, 32'sd94643, 32'sd1529836, -32'sd441683, 32'sd1828185, 32'sd673281, -32'sd1217992, -32'sd90311, -32'sd1911996, -32'sd1418502, -32'sd1178367, 32'sd654021, 32'sd173748, -32'sd2027930, -32'sd150310, -32'sd375990, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd583417, -32'sd34010, 32'sd666112, 32'sd1362183, 32'sd1701465, 32'sd3309303, 32'sd1843562, 32'sd1355254, 32'sd1491820, 32'sd129681, 32'sd1157703, 32'sd1500300, 32'sd276985, -32'sd1275260, 32'sd284920, -32'sd125041, 32'sd1575774, 32'sd1474420, 32'sd1296135, -32'sd511885, -32'sd1227395, 32'sd1061477, -32'sd555229, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd674301, 32'sd1099846, 32'sd864384, -32'sd678127, 32'sd720759, 32'sd148175, -32'sd1977519, -32'sd225727, 32'sd650961, 32'sd134927, -32'sd302713, 32'sd1453695, 32'sd439969, 32'sd692787, -32'sd338167, 32'sd1127917, -32'sd386022, -32'sd766172, -32'sd367024, -32'sd339032, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd788482, -32'sd998117, 32'sd552965, -32'sd714939, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd854178, 32'sd570370, -32'sd805330, -32'sd799985, 32'sd887375, -32'sd2258918, -32'sd1246924, 32'sd832165, 32'sd1235695, 32'sd148976, 32'sd19052, 32'sd316065, 32'sd936013, -32'sd196709, 32'sd1123727, 32'sd1718171, -32'sd155088, 32'sd1267967, 32'sd1322090, 32'sd91410, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd80807, 32'sd1429146, 32'sd531287, 32'sd64264, -32'sd990198, -32'sd596450, 32'sd402529, -32'sd361603, -32'sd2017585, 32'sd487904, 32'sd1023627, -32'sd401974, 32'sd1429193, 32'sd2030618, 32'sd107068, 32'sd119478, -32'sd664927, 32'sd380329, 32'sd1086293, -32'sd377628, 32'sd1641031, 32'sd963134, 32'sd838105, 32'sd1742735, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd438413, -32'sd248556, 32'sd532018, -32'sd837690, -32'sd1220429, -32'sd1501635, -32'sd678042, -32'sd514645, 32'sd2081269, 32'sd1263553, 32'sd1029471, 32'sd486588, 32'sd2625142, 32'sd485396, 32'sd1375124, -32'sd751794, 32'sd610248, -32'sd302208, 32'sd1189729, 32'sd834594, -32'sd90479, 32'sd126243, -32'sd443648, 32'sd807890, -32'sd70998, 32'sd0, 32'sd0, 32'sd797750, 32'sd958733, -32'sd1519496, 32'sd242601, 32'sd29388, -32'sd1448909, -32'sd717977, -32'sd578344, 32'sd1639967, 32'sd759730, 32'sd998800, 32'sd354515, -32'sd242078, 32'sd2344031, 32'sd2495945, 32'sd905604, 32'sd508289, -32'sd622021, 32'sd395727, 32'sd1224275, 32'sd554678, -32'sd28484, -32'sd1400594, -32'sd700062, -32'sd900401, -32'sd176471, 32'sd1503447, 32'sd0, 32'sd540372, -32'sd157881, -32'sd1188944, -32'sd670819, -32'sd1608140, -32'sd1057710, 32'sd46251, -32'sd537064, 32'sd283960, 32'sd1193043, 32'sd1223204, 32'sd1617296, 32'sd235682, 32'sd2759054, 32'sd837250, -32'sd614197, 32'sd1257488, 32'sd701528, -32'sd839258, -32'sd1305965, 32'sd51480, 32'sd694513, -32'sd642655, 32'sd1039000, 32'sd1113993, 32'sd521742, 32'sd534160, 32'sd0, 32'sd526759, 32'sd605733, -32'sd569957, -32'sd366306, -32'sd2624973, -32'sd825455, 32'sd543155, 32'sd105248, -32'sd869864, 32'sd907889, 32'sd1017464, 32'sd1295062, 32'sd2115192, 32'sd847331, -32'sd996803, -32'sd2441294, 32'sd981906, -32'sd492631, 32'sd161286, 32'sd187619, -32'sd842123, 32'sd2164716, -32'sd452420, 32'sd154407, 32'sd706985, -32'sd117357, 32'sd593438, 32'sd133377, 32'sd710397, -32'sd589031, -32'sd274027, -32'sd2176940, -32'sd3346932, -32'sd1022989, -32'sd636956, -32'sd1186504, 32'sd1164211, 32'sd1136022, 32'sd2040214, 32'sd433405, 32'sd869643, -32'sd823654, -32'sd539198, -32'sd2198331, -32'sd1245996, -32'sd687469, -32'sd1606068, 32'sd576936, 32'sd1884171, 32'sd3906486, 32'sd136940, 32'sd100281, 32'sd703170, -32'sd1139125, 32'sd625611, 32'sd305425, 32'sd1316347, -32'sd1653764, -32'sd297034, -32'sd2902608, -32'sd2277378, -32'sd412689, -32'sd877016, 32'sd876977, 32'sd1023735, 32'sd1782534, 32'sd1488529, 32'sd618599, 32'sd608531, -32'sd1230099, -32'sd1100827, -32'sd1297256, -32'sd2308993, -32'sd1219143, -32'sd1966930, 32'sd83505, -32'sd244662, 32'sd147466, -32'sd369045, -32'sd1226382, -32'sd1606642, -32'sd143533, 32'sd242234, -32'sd490021, 32'sd34526, 32'sd267820, 32'sd1738001, -32'sd691238, -32'sd2604127, 32'sd1256941, 32'sd183814, 32'sd1343093, 32'sd1677410, 32'sd233200, -32'sd545889, -32'sd315072, -32'sd2820598, -32'sd3756686, -32'sd1491382, -32'sd745012, -32'sd2268553, -32'sd1642810, -32'sd2665745, -32'sd561694, -32'sd590402, 32'sd217229, -32'sd1113835, -32'sd367176, -32'sd159741, -32'sd807235, -32'sd182823, 32'sd88842, 32'sd977296, -32'sd382913, -32'sd1188840, -32'sd2939049, -32'sd1315953, 32'sd616649, 32'sd1834146, 32'sd2106969, 32'sd2685110, 32'sd563845, -32'sd2650978, -32'sd414019, -32'sd2447287, -32'sd3327152, -32'sd2155697, 32'sd182183, 32'sd1088247, -32'sd1457392, -32'sd2698284, -32'sd306157, -32'sd631485, -32'sd1155721, -32'sd208217, 32'sd2452134, 32'sd1069876, -32'sd659601, 32'sd166830, 32'sd208619, -32'sd196298, 32'sd549677, -32'sd507679, -32'sd1640528, -32'sd1036063, -32'sd552367, 32'sd2171387, 32'sd3236693, 32'sd1244969, -32'sd1452201, 32'sd38955, 32'sd2331249, 32'sd858238, -32'sd1656756, -32'sd2045363, -32'sd228436, 32'sd3570225, 32'sd684982, -32'sd1608142, -32'sd2523339, -32'sd2123600, -32'sd1246517, 32'sd2057661, 32'sd1610681, -32'sd196330, -32'sd688391, -32'sd532297, 32'sd315223, -32'sd560813, 32'sd138831, -32'sd810912, -32'sd2094324, -32'sd1577869, 32'sd316779, 32'sd113375, 32'sd1769350, 32'sd1976681, 32'sd68388, 32'sd730280, 32'sd822210, 32'sd2188457, -32'sd538585, -32'sd1506962, -32'sd642031, 32'sd2136122, 32'sd2407314, 32'sd571110, -32'sd1559551, -32'sd1582115, -32'sd2888072, -32'sd1012103, 32'sd1963867, -32'sd2211641, -32'sd110442, 32'sd1176111, 32'sd102066, -32'sd470540, -32'sd391131, -32'sd1232909, -32'sd4543729, -32'sd3201238, 32'sd254253, 32'sd2278031, 32'sd1465918, 32'sd878914, 32'sd533861, 32'sd1045379, 32'sd2155287, 32'sd1138747, 32'sd2341969, 32'sd1560226, 32'sd836678, -32'sd1933863, 32'sd980134, 32'sd1095616, 32'sd1245491, -32'sd1061386, -32'sd881202, 32'sd773443, -32'sd45196, -32'sd1910457, -32'sd24649, 32'sd663638, 32'sd1573619, -32'sd282485, 32'sd193264, -32'sd57087, -32'sd2682709, -32'sd1510758, -32'sd1775024, -32'sd857005, 32'sd1995687, -32'sd744923, 32'sd173781, 32'sd141850, -32'sd271888, -32'sd192028, 32'sd1602750, 32'sd818019, 32'sd442279, 32'sd1249016, 32'sd325829, -32'sd542709, 32'sd897777, -32'sd655845, 32'sd1340956, 32'sd527196, 32'sd1273902, -32'sd203192, 32'sd605359, -32'sd404919, 32'sd83279, 32'sd889092, 32'sd1785463, 32'sd157479, -32'sd347709, -32'sd1570243, 32'sd25747, -32'sd95093, 32'sd1190136, 32'sd137853, -32'sd292869, 32'sd89220, -32'sd120207, 32'sd380236, 32'sd1262566, 32'sd615555, 32'sd637437, 32'sd448582, 32'sd1181803, -32'sd1556733, -32'sd52600, -32'sd582143, -32'sd916597, -32'sd154808, -32'sd496431, -32'sd1784677, 32'sd924128, 32'sd1009039, 32'sd628928, -32'sd724058, -32'sd18595, -32'sd424205, 32'sd1050564, 32'sd160772, -32'sd1006720, 32'sd477918, 32'sd2030177, 32'sd1202680, -32'sd1031358, 32'sd1162019, 32'sd637174, 32'sd2322157, 32'sd964202, -32'sd64455, 32'sd2318789, 32'sd1202793, 32'sd1576000, -32'sd885731, -32'sd2241404, -32'sd1427367, -32'sd1629305, 32'sd1257240, -32'sd1482909, 32'sd913919, -32'sd370504, 32'sd1258407, 32'sd0, 32'sd628230, 32'sd1417144, -32'sd1814896, -32'sd5225, -32'sd1510732, -32'sd308500, 32'sd72265, -32'sd1567591, -32'sd884840, 32'sd1077425, 32'sd1712483, 32'sd2905360, 32'sd2226046, -32'sd2032396, 32'sd329835, 32'sd2906270, 32'sd262817, 32'sd700702, -32'sd582202, 32'sd687225, 32'sd188713, 32'sd2457396, 32'sd778953, -32'sd346860, 32'sd141600, -32'sd1174427, 32'sd662617, 32'sd138671, -32'sd401862, -32'sd254393, -32'sd17309, -32'sd2206969, -32'sd2154062, -32'sd1235383, -32'sd1536752, -32'sd13786, -32'sd966217, -32'sd1390023, -32'sd1130565, 32'sd217617, 32'sd1396720, -32'sd2219939, -32'sd1256392, -32'sd944759, 32'sd22769, 32'sd1454283, -32'sd928094, 32'sd394119, 32'sd119330, 32'sd844479, -32'sd307040, -32'sd95001, 32'sd1637022, -32'sd423892, 32'sd6905, 32'sd257289, -32'sd145907, -32'sd315713, -32'sd313480, -32'sd2123200, -32'sd2412156, -32'sd832112, -32'sd1975045, 32'sd1457409, 32'sd1569368, -32'sd1630095, -32'sd2202395, 32'sd3378759, 32'sd478673, -32'sd293241, -32'sd1072216, -32'sd2901905, -32'sd673099, 32'sd1718821, 32'sd592724, -32'sd486827, 32'sd2131302, -32'sd193744, -32'sd731663, -32'sd1001771, 32'sd848121, -32'sd2367978, -32'sd2125249, 32'sd0, -32'sd67992, -32'sd1993757, 32'sd74965, -32'sd1763274, -32'sd1040848, -32'sd61663, -32'sd521948, -32'sd1364665, 32'sd1489844, -32'sd1408350, -32'sd26689, -32'sd244903, 32'sd1606803, -32'sd136233, -32'sd388626, -32'sd1862663, -32'sd1190620, 32'sd820267, 32'sd674225, 32'sd1243319, 32'sd1718196, 32'sd1579343, -32'sd1549975, -32'sd2192203, 32'sd125954, -32'sd239076, 32'sd900071, 32'sd549360, -32'sd703109, -32'sd314002, -32'sd107375, 32'sd967862, 32'sd1060442, 32'sd489752, -32'sd536560, 32'sd1528721, 32'sd484912, 32'sd414111, -32'sd375068, 32'sd960492, -32'sd311451, 32'sd963693, -32'sd277013, -32'sd551487, 32'sd1919729, 32'sd1891482, 32'sd2139427, 32'sd823596, 32'sd1366389, 32'sd317011, 32'sd181908, -32'sd119099, -32'sd1159403, -32'sd951078, 32'sd546167, 32'sd1133269, 32'sd1618832, 32'sd458355, -32'sd2023490, -32'sd723133, 32'sd10058, -32'sd562973, -32'sd1169038, -32'sd567015, 32'sd323835, 32'sd263593, 32'sd439721, -32'sd1995588, -32'sd1321914, -32'sd585273, 32'sd927665, 32'sd441314, 32'sd1760269, 32'sd1468454, 32'sd1367864, -32'sd814963, -32'sd1954309, -32'sd961496, -32'sd196033, -32'sd946298, 32'sd516084, -32'sd1801204, 32'sd729624, 32'sd0, 32'sd792102, -32'sd1345372, 32'sd654797, 32'sd1234001, 32'sd1319922, -32'sd590129, -32'sd1438385, 32'sd1865647, -32'sd852514, 32'sd219406, 32'sd84362, 32'sd250889, -32'sd1212282, 32'sd1218536, 32'sd1229852, 32'sd1042449, 32'sd2776901, -32'sd481096, 32'sd305382, -32'sd96177, -32'sd2834944, 32'sd32381, -32'sd247402, 32'sd796224, -32'sd1127123, -32'sd20199, 32'sd0, 32'sd0, 32'sd0, 32'sd718365, -32'sd1429319, -32'sd659219, 32'sd327727, -32'sd1099207, 32'sd298184, 32'sd72770, 32'sd881696, -32'sd1576339, -32'sd1151313, 32'sd1164863, 32'sd1954863, -32'sd37588, 32'sd1550427, 32'sd3027707, -32'sd926740, -32'sd1543413, -32'sd27452, 32'sd817331, -32'sd1228508, -32'sd720099, 32'sd467199, 32'sd887358, 32'sd675946, 32'sd1302306, 32'sd0, 32'sd0, 32'sd0, -32'sd28272, -32'sd115715, 32'sd904989, -32'sd107813, 32'sd5988, -32'sd229105, 32'sd160272, -32'sd508054, 32'sd1209976, 32'sd1627639, 32'sd2680702, 32'sd770296, 32'sd771352, 32'sd1698636, 32'sd741215, 32'sd1490519, 32'sd2755517, 32'sd829741, 32'sd1470848, 32'sd1612889, 32'sd170448, 32'sd1398304, 32'sd1508137, 32'sd972986, -32'sd1135928, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1212656, 32'sd532814, -32'sd1387247, -32'sd1233802, 32'sd511720, 32'sd364969, -32'sd472643, -32'sd336688, 32'sd399153, 32'sd758170, 32'sd226709, 32'sd182763, 32'sd616729, -32'sd513003, 32'sd1597308, 32'sd290576, 32'sd571595, 32'sd518757, 32'sd80640, 32'sd1017063, 32'sd2046996, 32'sd396691, 32'sd571853, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd227296, 32'sd252465, 32'sd1136461, 32'sd200039, -32'sd184682, -32'sd297944, -32'sd184165, -32'sd185610, 32'sd168155, 32'sd741933, 32'sd1057706, 32'sd1230918, 32'sd201870, -32'sd1343987, 32'sd1113825, 32'sd550667, 32'sd498872, -32'sd1909168, -32'sd150888, -32'sd15959, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd123063, -32'sd492704, 32'sd182318, 32'sd414393, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1040915, 32'sd1506552, -32'sd1004137, -32'sd795254, -32'sd557840, -32'sd1398832, 32'sd540176, -32'sd874479, 32'sd259255, 32'sd41533, 32'sd843664, -32'sd730883, 32'sd663805, 32'sd1938658, 32'sd458031, 32'sd1557282, 32'sd49904, 32'sd1407574, 32'sd1565561, 32'sd1032781, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd693294, 32'sd1205751, 32'sd894353, -32'sd323769, -32'sd553403, -32'sd116798, -32'sd415711, -32'sd1177371, 32'sd367868, -32'sd1026878, -32'sd214347, 32'sd2294580, 32'sd774859, 32'sd266986, 32'sd597401, 32'sd1553426, 32'sd1656640, 32'sd2320153, 32'sd746743, 32'sd234443, 32'sd1516635, 32'sd198008, 32'sd413765, 32'sd1774738, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1937601, 32'sd839974, 32'sd107147, -32'sd1268339, 32'sd120633, -32'sd851641, -32'sd2235579, 32'sd572194, 32'sd1633856, -32'sd3373778, -32'sd925323, 32'sd276924, 32'sd330256, -32'sd624223, 32'sd1752011, 32'sd2335777, 32'sd3603472, 32'sd1004388, 32'sd2156597, 32'sd1251888, -32'sd335620, -32'sd20998, -32'sd11116, -32'sd334419, -32'sd547250, 32'sd0, 32'sd0, 32'sd682579, 32'sd602045, -32'sd918339, -32'sd649495, -32'sd530455, -32'sd1260913, 32'sd405851, -32'sd1604425, 32'sd1313281, -32'sd1078993, -32'sd2802694, 32'sd375873, 32'sd342097, 32'sd207979, 32'sd1507643, 32'sd81791, 32'sd759105, 32'sd809150, -32'sd441507, 32'sd406124, 32'sd2813006, 32'sd499233, 32'sd888934, -32'sd601085, -32'sd359784, 32'sd896010, 32'sd936076, 32'sd0, 32'sd1005061, -32'sd1303556, 32'sd197282, 32'sd154303, -32'sd109018, -32'sd68247, 32'sd821875, 32'sd1698402, -32'sd989937, -32'sd1320616, -32'sd348850, -32'sd2240429, -32'sd1459773, -32'sd762346, 32'sd1004850, 32'sd629846, 32'sd1423563, 32'sd2706154, 32'sd74153, 32'sd1583340, -32'sd129322, 32'sd1149304, 32'sd1448624, -32'sd1106617, 32'sd718112, -32'sd519431, 32'sd57282, 32'sd0, 32'sd207910, 32'sd797425, -32'sd253880, -32'sd1246539, -32'sd174177, 32'sd987640, 32'sd1511719, 32'sd846678, -32'sd14814, 32'sd264476, 32'sd1505704, 32'sd2230956, 32'sd1659141, 32'sd1966824, 32'sd1313843, 32'sd2824382, 32'sd3246960, 32'sd2160133, 32'sd3402516, 32'sd1158144, 32'sd1222899, -32'sd682008, 32'sd1034776, 32'sd1309236, 32'sd2177726, 32'sd575320, 32'sd512789, 32'sd1799687, 32'sd683653, 32'sd619765, 32'sd153478, 32'sd448002, 32'sd424261, 32'sd189581, 32'sd1819101, 32'sd449784, 32'sd644972, 32'sd1061082, 32'sd68077, 32'sd253830, 32'sd1374505, 32'sd895914, 32'sd801018, 32'sd2326872, 32'sd2799202, 32'sd3629447, 32'sd1445587, 32'sd2844574, 32'sd182048, 32'sd926438, 32'sd2184673, 32'sd1018443, 32'sd1557665, 32'sd821841, 32'sd406440, 32'sd745387, 32'sd1742935, 32'sd1343136, -32'sd1341818, -32'sd1295989, -32'sd465388, 32'sd260986, 32'sd2632368, -32'sd1133100, 32'sd2027232, 32'sd1566709, 32'sd465465, -32'sd650034, -32'sd5496, 32'sd48685, 32'sd1175580, 32'sd870386, 32'sd655087, 32'sd248422, -32'sd2489761, 32'sd62504, -32'sd1411829, -32'sd1664348, 32'sd1132527, 32'sd71400, -32'sd1843116, 32'sd173503, -32'sd165191, 32'sd471037, 32'sd1062267, -32'sd1662922, -32'sd360427, 32'sd865153, -32'sd1122067, 32'sd2220845, 32'sd495761, -32'sd708234, 32'sd155456, 32'sd2392129, 32'sd1538412, 32'sd840700, 32'sd1109349, 32'sd685345, -32'sd389921, -32'sd4896234, -32'sd3154988, -32'sd3540304, -32'sd3622142, -32'sd3217029, -32'sd2441001, -32'sd2156072, -32'sd1685921, 32'sd1282505, -32'sd767607, 32'sd648690, -32'sd120202, 32'sd1813801, 32'sd974771, 32'sd371881, -32'sd1227909, 32'sd806421, 32'sd772455, 32'sd2004780, -32'sd651757, 32'sd1419141, -32'sd279414, 32'sd3028531, 32'sd1216444, 32'sd1215682, 32'sd737221, -32'sd2000198, -32'sd2175986, -32'sd1965297, -32'sd3619430, -32'sd1929710, -32'sd3658472, -32'sd4937845, -32'sd3900794, -32'sd2157517, -32'sd1531827, -32'sd2058710, -32'sd1717608, 32'sd216522, 32'sd206502, 32'sd1319429, -32'sd114247, -32'sd556372, 32'sd760661, 32'sd211689, 32'sd1538056, 32'sd1470390, 32'sd49006, -32'sd1226615, -32'sd919135, -32'sd643953, -32'sd247156, -32'sd2063308, -32'sd3298066, -32'sd2340808, 32'sd930160, 32'sd781662, 32'sd128412, -32'sd681935, -32'sd3044951, -32'sd3585531, -32'sd3329608, -32'sd639379, -32'sd1216878, -32'sd2064800, -32'sd624742, 32'sd689880, -32'sd1196219, 32'sd330239, -32'sd1078717, -32'sd115644, 32'sd1569288, 32'sd1574029, 32'sd690397, 32'sd355617, 32'sd269507, 32'sd1110647, 32'sd939515, 32'sd525451, -32'sd587457, -32'sd1596023, -32'sd1102214, -32'sd148516, 32'sd1236788, 32'sd1201704, 32'sd1294005, 32'sd1430714, -32'sd758536, -32'sd1407320, -32'sd2837967, -32'sd108965, -32'sd2499431, -32'sd178368, -32'sd1384885, 32'sd960110, -32'sd665806, 32'sd725330, 32'sd1333280, -32'sd243701, 32'sd917485, 32'sd1736887, 32'sd1074831, -32'sd373558, -32'sd423531, 32'sd429046, -32'sd2604497, -32'sd2444910, -32'sd829621, -32'sd2198408, -32'sd2053750, -32'sd910950, -32'sd217763, 32'sd975839, 32'sd1391478, 32'sd34948, 32'sd1189796, -32'sd1581639, -32'sd733276, 32'sd392951, -32'sd826342, -32'sd1488306, -32'sd991748, 32'sd1042806, 32'sd481716, 32'sd869680, -32'sd730962, 32'sd197921, 32'sd435201, -32'sd127510, 32'sd685175, -32'sd808761, -32'sd1657976, -32'sd986551, -32'sd2402753, -32'sd1188517, -32'sd1726822, -32'sd2061490, -32'sd1102683, -32'sd1337816, 32'sd2476713, 32'sd3975121, -32'sd153744, -32'sd769509, 32'sd1017216, 32'sd1042858, 32'sd599746, 32'sd143373, 32'sd134214, -32'sd107622, -32'sd794884, -32'sd296704, 32'sd36666, 32'sd1836147, 32'sd514958, -32'sd377866, -32'sd227953, -32'sd569933, 32'sd1183783, -32'sd618883, -32'sd2563364, -32'sd664780, -32'sd542099, 32'sd545588, -32'sd2527847, -32'sd2080420, -32'sd2003798, 32'sd767054, 32'sd3125352, 32'sd2976644, 32'sd1373015, 32'sd650107, 32'sd1159050, -32'sd198584, 32'sd194909, -32'sd180405, -32'sd1386948, -32'sd922463, -32'sd1495366, 32'sd162458, 32'sd1046568, 32'sd1175320, 32'sd671995, 32'sd377197, 32'sd762540, -32'sd1178981, -32'sd1083033, 32'sd295681, -32'sd438658, -32'sd1071472, -32'sd258220, 32'sd510402, 32'sd330436, -32'sd630958, -32'sd421340, 32'sd2566648, 32'sd5376877, 32'sd2761407, 32'sd1457379, -32'sd157170, 32'sd2135738, 32'sd814713, 32'sd2216305, -32'sd579501, 32'sd345116, 32'sd1575743, 32'sd703660, -32'sd189452, 32'sd1111734, 32'sd0, -32'sd84990, 32'sd1388552, 32'sd1420236, -32'sd467661, -32'sd1425308, 32'sd1230189, -32'sd66228, 32'sd2637092, 32'sd1348678, -32'sd471570, -32'sd1088608, -32'sd979078, -32'sd1082146, 32'sd2606103, 32'sd4029122, 32'sd2641680, 32'sd1688130, 32'sd765040, 32'sd254978, 32'sd2555368, 32'sd604851, -32'sd715480, 32'sd649680, 32'sd1678985, 32'sd240644, 32'sd1709474, 32'sd587891, -32'sd111012, 32'sd538469, 32'sd1432816, 32'sd409120, 32'sd221471, -32'sd1121259, 32'sd1074644, 32'sd137051, 32'sd1075492, -32'sd132148, -32'sd1673046, -32'sd2053641, -32'sd4851776, -32'sd2148659, 32'sd1954103, 32'sd3452940, 32'sd3153794, -32'sd329454, -32'sd1427856, 32'sd1095261, 32'sd64430, 32'sd167139, 32'sd1136257, 32'sd851006, 32'sd530477, 32'sd530743, -32'sd846930, -32'sd493203, 32'sd1463756, -32'sd114608, 32'sd730623, 32'sd535335, 32'sd1249128, -32'sd4327, -32'sd2019838, -32'sd811503, -32'sd759355, 32'sd127638, -32'sd2666733, -32'sd1735156, -32'sd2496045, -32'sd1673325, 32'sd2529676, 32'sd2336477, 32'sd2305886, -32'sd541924, 32'sd1066863, -32'sd469822, 32'sd1224473, 32'sd1095302, 32'sd1062120, -32'sd380331, 32'sd1931475, 32'sd548925, 32'sd20531, -32'sd2065430, 32'sd0, 32'sd848545, 32'sd1459087, -32'sd102845, 32'sd1357614, 32'sd993007, 32'sd342904, -32'sd1103303, -32'sd1268369, -32'sd937336, -32'sd1625557, -32'sd1869161, -32'sd1632858, 32'sd787530, 32'sd1428835, 32'sd1636622, 32'sd3316276, 32'sd2209020, 32'sd3825628, 32'sd361411, 32'sd645306, 32'sd1242978, 32'sd1357405, 32'sd563917, 32'sd1298696, -32'sd1597637, -32'sd1551262, 32'sd1299254, 32'sd1220199, -32'sd603013, 32'sd450239, 32'sd1322359, 32'sd2006304, 32'sd1341303, 32'sd456660, -32'sd235832, 32'sd441652, 32'sd1107364, -32'sd558574, 32'sd155056, 32'sd1283394, 32'sd1019952, 32'sd2023470, 32'sd1522808, 32'sd2437104, 32'sd1834902, 32'sd2156077, 32'sd292344, -32'sd454393, 32'sd1094134, 32'sd1276231, -32'sd542561, 32'sd1037780, 32'sd520142, 32'sd668953, -32'sd59623, 32'sd758048, -32'sd6859, -32'sd636180, -32'sd703827, 32'sd2218014, -32'sd528368, -32'sd1955314, 32'sd908904, -32'sd239920, 32'sd938843, 32'sd669572, 32'sd500674, 32'sd38147, 32'sd362899, 32'sd3302730, 32'sd3236785, 32'sd594991, -32'sd252391, 32'sd473347, 32'sd183810, 32'sd56432, -32'sd1542738, -32'sd3147412, 32'sd402403, -32'sd84713, 32'sd646226, -32'sd1801310, 32'sd401047, 32'sd0, 32'sd1066018, -32'sd947536, 32'sd446724, -32'sd567286, -32'sd1065784, -32'sd1215889, 32'sd835679, -32'sd1057162, 32'sd454842, 32'sd1182900, -32'sd1981862, 32'sd442315, 32'sd1408834, 32'sd2083261, 32'sd1970272, -32'sd1028196, -32'sd215490, -32'sd2819895, 32'sd597267, -32'sd1443574, -32'sd3628374, -32'sd3347989, -32'sd1418941, -32'sd3178981, -32'sd1729350, -32'sd337703, 32'sd0, 32'sd0, 32'sd0, -32'sd406544, 32'sd32034, -32'sd52412, 32'sd161526, 32'sd600671, 32'sd128539, 32'sd341170, 32'sd620516, -32'sd1131567, 32'sd142833, 32'sd931349, -32'sd876885, 32'sd1293354, 32'sd78531, -32'sd1513993, 32'sd456512, -32'sd1343883, -32'sd387453, -32'sd992155, -32'sd823390, -32'sd10358, 32'sd43594, 32'sd1393227, 32'sd1731184, 32'sd745660, 32'sd0, 32'sd0, 32'sd0, -32'sd42174, 32'sd364339, -32'sd737325, 32'sd536895, 32'sd354140, -32'sd1417116, -32'sd1633884, 32'sd901480, -32'sd819609, -32'sd183296, 32'sd1391654, 32'sd2630972, 32'sd2436699, 32'sd1303727, -32'sd1119277, -32'sd1544516, 32'sd80476, 32'sd373728, 32'sd74027, 32'sd1398166, -32'sd955847, -32'sd724676, 32'sd981827, 32'sd1143855, 32'sd566529, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd662693, 32'sd969006, -32'sd706075, 32'sd2878672, -32'sd536150, -32'sd640318, -32'sd666520, -32'sd178466, 32'sd261530, -32'sd1989085, 32'sd201671, -32'sd191018, -32'sd427086, 32'sd1596063, -32'sd755421, 32'sd892168, 32'sd738837, 32'sd1119046, -32'sd1505711, -32'sd387621, -32'sd935629, 32'sd1429533, 32'sd1416770, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1998055, 32'sd702861, 32'sd1033136, 32'sd1479178, 32'sd617874, 32'sd1122509, -32'sd120397, 32'sd1082026, 32'sd2110308, 32'sd1059577, 32'sd1404723, 32'sd1166535, 32'sd17415, 32'sd1454110, 32'sd1509552, -32'sd416873, -32'sd974038, 32'sd494939, -32'sd556065, 32'sd695719, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd985613, -32'sd771515, -32'sd340603, 32'sd478049, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd824933, 32'sd1728647, -32'sd1737699, -32'sd441798, 32'sd257682, -32'sd1918159, 32'sd132113, 32'sd631138, -32'sd336338, 32'sd1125400, 32'sd998212, -32'sd628387, 32'sd865329, 32'sd2147065, 32'sd915450, 32'sd923327, 32'sd849847, 32'sd1484801, 32'sd436639, 32'sd854047, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd813107, 32'sd1684877, 32'sd411543, 32'sd1182208, 32'sd694917, 32'sd39683, -32'sd1172080, -32'sd607387, -32'sd445097, -32'sd491759, 32'sd1325572, -32'sd451246, 32'sd215030, -32'sd1825113, 32'sd540072, -32'sd17384, 32'sd543434, 32'sd1111994, -32'sd111888, -32'sd295761, 32'sd1000635, 32'sd804456, -32'sd290171, 32'sd818578, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd422416, 32'sd129046, -32'sd411148, -32'sd149227, 32'sd1650025, 32'sd1610905, 32'sd2354364, -32'sd801417, 32'sd662198, -32'sd331695, -32'sd744520, -32'sd995794, 32'sd2156625, 32'sd491285, -32'sd593167, 32'sd187288, -32'sd1237740, -32'sd2307451, -32'sd1138733, -32'sd783880, 32'sd1432076, -32'sd69885, 32'sd1183617, 32'sd615648, 32'sd1666307, 32'sd0, 32'sd0, 32'sd878549, 32'sd864934, 32'sd606132, 32'sd23436, 32'sd813609, 32'sd481695, -32'sd175974, 32'sd47571, -32'sd50241, -32'sd87359, 32'sd1169707, 32'sd1655074, 32'sd628659, 32'sd136803, -32'sd133021, 32'sd1209784, -32'sd1453210, 32'sd1304376, 32'sd259616, -32'sd2233046, 32'sd190717, -32'sd2413205, 32'sd891195, 32'sd1030259, 32'sd392900, 32'sd1193920, 32'sd1384178, 32'sd0, 32'sd728281, -32'sd400540, -32'sd945936, -32'sd948695, 32'sd902720, -32'sd1197209, 32'sd772884, -32'sd1056475, -32'sd1091047, 32'sd1509044, -32'sd148813, -32'sd590305, 32'sd207744, 32'sd1791186, 32'sd1548461, -32'sd529304, -32'sd2706177, -32'sd1886547, -32'sd351933, -32'sd466618, -32'sd809850, -32'sd701776, 32'sd527912, 32'sd550623, 32'sd240899, -32'sd848203, 32'sd230390, 32'sd0, 32'sd1007103, 32'sd845274, -32'sd393829, -32'sd326718, -32'sd767736, -32'sd2582354, -32'sd2456194, -32'sd1431100, 32'sd858443, -32'sd943738, -32'sd1848761, -32'sd862504, -32'sd699040, -32'sd352478, 32'sd162277, 32'sd243450, -32'sd1210677, -32'sd1575722, -32'sd3716893, -32'sd702689, -32'sd1014508, -32'sd828221, 32'sd48959, 32'sd179897, -32'sd1720980, -32'sd2005838, -32'sd718788, 32'sd641038, 32'sd307535, 32'sd1426407, -32'sd265616, -32'sd146994, 32'sd1607014, -32'sd164566, 32'sd1943, 32'sd901337, -32'sd909202, -32'sd524147, -32'sd1895144, -32'sd623477, 32'sd1536450, 32'sd237237, 32'sd1115422, 32'sd3324671, 32'sd544108, -32'sd1547170, -32'sd280933, -32'sd71061, 32'sd231063, -32'sd1385839, 32'sd398744, 32'sd511099, 32'sd388721, 32'sd723221, 32'sd334646, 32'sd945279, 32'sd778697, -32'sd428418, 32'sd1746032, 32'sd1056232, -32'sd377891, -32'sd917310, 32'sd1335267, 32'sd1685095, 32'sd481793, -32'sd2099520, -32'sd2502088, -32'sd2091499, -32'sd1722072, 32'sd675703, 32'sd1489357, 32'sd2621412, 32'sd1574851, 32'sd53831, 32'sd529498, 32'sd1034896, -32'sd641423, -32'sd2074582, -32'sd2057442, 32'sd8280, 32'sd1660558, 32'sd1268814, 32'sd674471, -32'sd114441, -32'sd247115, 32'sd2365981, -32'sd201326, -32'sd645301, 32'sd116704, 32'sd3717, -32'sd361793, 32'sd2049637, -32'sd825588, -32'sd736131, -32'sd198344, -32'sd2258688, -32'sd1187241, 32'sd1775737, 32'sd214777, 32'sd547003, 32'sd1300349, -32'sd817971, 32'sd1842040, -32'sd1538404, 32'sd578715, -32'sd100937, -32'sd742351, -32'sd353319, -32'sd455529, 32'sd1172645, -32'sd144375, -32'sd470329, 32'sd1640935, 32'sd315310, 32'sd954435, -32'sd868068, 32'sd983454, -32'sd1075453, 32'sd1042543, 32'sd48927, -32'sd1525170, -32'sd844670, -32'sd1733958, -32'sd1701147, 32'sd1392425, 32'sd1147340, -32'sd726709, -32'sd1443322, 32'sd933050, -32'sd695644, 32'sd1502934, -32'sd439833, -32'sd241176, 32'sd69023, 32'sd580935, 32'sd187768, 32'sd865028, 32'sd261155, 32'sd1374074, -32'sd476755, -32'sd473438, 32'sd917816, -32'sd1934735, -32'sd1595784, -32'sd344170, -32'sd734192, 32'sd921250, 32'sd1118640, -32'sd1051077, -32'sd624009, -32'sd1797935, 32'sd56752, 32'sd2009214, 32'sd997539, 32'sd1296870, -32'sd78970, 32'sd19743, -32'sd893281, 32'sd1362368, 32'sd1434221, 32'sd1270263, 32'sd1141250, 32'sd1533818, -32'sd205479, -32'sd1979854, 32'sd665635, 32'sd364602, 32'sd1713126, 32'sd1097884, 32'sd870861, -32'sd2532757, 32'sd17370, -32'sd1334232, 32'sd443270, 32'sd1524850, 32'sd1417807, -32'sd538357, -32'sd109248, -32'sd1070088, 32'sd2315899, 32'sd3341277, 32'sd3114755, 32'sd687702, 32'sd1725147, -32'sd66921, 32'sd1061127, 32'sd41464, 32'sd117717, 32'sd143018, 32'sd2097458, 32'sd1860725, 32'sd3388287, 32'sd2336493, 32'sd76216, -32'sd1146604, 32'sd845515, -32'sd1353105, 32'sd437139, -32'sd995355, -32'sd1916408, 32'sd1078840, 32'sd2095537, 32'sd1956685, 32'sd1216659, -32'sd952884, -32'sd465163, 32'sd2395188, 32'sd2965441, 32'sd1758408, 32'sd1663278, 32'sd1435210, 32'sd2562397, 32'sd1352502, 32'sd1315891, -32'sd1889221, 32'sd244409, -32'sd1153327, -32'sd909018, 32'sd1613518, 32'sd1789603, -32'sd1473093, 32'sd462991, 32'sd133660, 32'sd2139501, -32'sd377233, -32'sd371621, -32'sd1160677, -32'sd2492056, 32'sd846584, -32'sd845668, 32'sd763648, 32'sd642388, 32'sd649488, -32'sd129484, 32'sd1250046, 32'sd3343487, 32'sd3476304, 32'sd2180633, -32'sd130562, 32'sd603339, 32'sd809404, -32'sd1670285, -32'sd2971796, -32'sd756866, -32'sd1733812, 32'sd626692, 32'sd1725894, 32'sd2181594, -32'sd1053541, 32'sd588771, 32'sd863078, 32'sd1861490, 32'sd1235560, 32'sd562776, 32'sd209884, -32'sd798747, 32'sd328348, -32'sd397518, -32'sd1224473, -32'sd479016, -32'sd2376009, -32'sd942246, 32'sd2021184, 32'sd2387263, -32'sd357901, -32'sd306660, 32'sd44198, 32'sd300313, -32'sd437475, 32'sd1067574, -32'sd2033698, 32'sd701662, -32'sd617160, -32'sd783774, 32'sd870965, 32'sd683716, -32'sd568968, 32'sd1746752, 32'sd212605, 32'sd744835, 32'sd1034804, 32'sd1430335, -32'sd1199597, -32'sd1636480, -32'sd1709699, -32'sd3542880, -32'sd3954101, -32'sd3349167, -32'sd4593871, -32'sd943891, 32'sd409090, -32'sd254536, -32'sd846459, -32'sd1592052, -32'sd3077161, 32'sd94111, 32'sd494596, 32'sd1639048, -32'sd878319, 32'sd1645495, -32'sd41957, 32'sd478740, 32'sd1311764, -32'sd254984, -32'sd752656, 32'sd318731, -32'sd375868, 32'sd0, -32'sd276446, -32'sd841035, -32'sd183164, 32'sd922483, 32'sd95206, -32'sd1934404, -32'sd3107034, -32'sd2806835, -32'sd3106373, -32'sd3130587, -32'sd1262678, -32'sd1344780, -32'sd1693326, -32'sd743085, -32'sd1097008, -32'sd275151, -32'sd1851453, -32'sd1422743, 32'sd306005, -32'sd432225, 32'sd838880, 32'sd155433, -32'sd1216332, 32'sd797871, -32'sd540708, 32'sd510948, 32'sd398146, -32'sd125004, 32'sd543597, -32'sd968955, 32'sd1572359, -32'sd463970, 32'sd1147040, 32'sd1408262, -32'sd1292998, -32'sd2529729, -32'sd996014, -32'sd1188236, -32'sd1427945, -32'sd1420815, -32'sd723896, -32'sd1666219, 32'sd57347, -32'sd434340, 32'sd256380, -32'sd154210, 32'sd1155802, -32'sd501259, 32'sd418471, -32'sd1480072, -32'sd1986624, -32'sd491576, -32'sd456925, -32'sd757477, 32'sd456697, 32'sd602810, 32'sd386963, 32'sd754951, 32'sd2143398, 32'sd1071893, 32'sd860075, 32'sd1474157, 32'sd1201748, 32'sd728263, 32'sd1572930, -32'sd674095, -32'sd1398978, -32'sd1046586, -32'sd487919, -32'sd1068349, -32'sd1733919, -32'sd407164, -32'sd345259, 32'sd2005439, 32'sd483321, -32'sd431628, 32'sd893420, -32'sd2469032, -32'sd2437255, -32'sd1618336, -32'sd1699911, 32'sd1158136, -32'sd142004, 32'sd0, -32'sd1162677, 32'sd295337, 32'sd316764, 32'sd913110, -32'sd537195, 32'sd765881, 32'sd2350491, 32'sd224570, 32'sd465479, 32'sd593803, -32'sd278292, -32'sd517394, -32'sd1831204, 32'sd1057367, 32'sd980090, 32'sd2061067, 32'sd1674881, 32'sd1879347, -32'sd1514191, -32'sd85365, -32'sd342907, -32'sd2808258, -32'sd1237801, -32'sd2171162, -32'sd1645643, 32'sd1717645, 32'sd544200, 32'sd2171144, 32'sd569211, 32'sd384146, -32'sd532038, 32'sd142511, -32'sd1000968, -32'sd609215, 32'sd103624, -32'sd931823, 32'sd605766, 32'sd1153715, 32'sd1625907, -32'sd71003, 32'sd148351, 32'sd1795968, -32'sd190248, 32'sd1253780, 32'sd584077, 32'sd930548, -32'sd284157, 32'sd1385794, -32'sd2515230, -32'sd416122, -32'sd1189519, -32'sd1698410, -32'sd416153, -32'sd269310, -32'sd509337, 32'sd1337038, 32'sd1091037, 32'sd622633, -32'sd422294, 32'sd1452424, -32'sd528279, -32'sd1463467, 32'sd292520, 32'sd390038, -32'sd759927, 32'sd1474747, -32'sd242266, -32'sd268030, -32'sd249300, 32'sd269468, -32'sd930101, 32'sd902213, -32'sd42108, -32'sd1225662, -32'sd940965, -32'sd1942498, -32'sd1569256, -32'sd1559177, 32'sd619582, -32'sd1687673, -32'sd364960, 32'sd1736675, 32'sd410860, 32'sd0, 32'sd733282, 32'sd254272, 32'sd2111484, 32'sd148144, 32'sd57851, -32'sd1279501, -32'sd517331, 32'sd712389, 32'sd208579, 32'sd3338233, 32'sd3146014, -32'sd70800, 32'sd71165, 32'sd395898, -32'sd1575531, -32'sd463673, 32'sd1016501, -32'sd678401, -32'sd1389291, 32'sd935756, -32'sd307942, -32'sd939834, 32'sd43804, 32'sd687141, 32'sd192088, 32'sd540051, 32'sd0, 32'sd0, 32'sd0, 32'sd424999, 32'sd1716957, 32'sd336751, 32'sd345589, -32'sd272633, 32'sd478397, -32'sd46192, 32'sd3434033, 32'sd2104152, -32'sd464690, -32'sd1229404, 32'sd1260821, 32'sd1952280, -32'sd363268, 32'sd1518381, 32'sd618111, 32'sd346651, 32'sd1622229, 32'sd112253, -32'sd1322164, -32'sd33127, -32'sd772429, 32'sd37784, 32'sd1068440, 32'sd185998, 32'sd0, 32'sd0, 32'sd0, 32'sd1251012, 32'sd1030701, 32'sd481211, -32'sd574126, 32'sd626635, -32'sd517584, -32'sd798159, 32'sd2034796, 32'sd491924, -32'sd1045166, -32'sd459267, -32'sd971517, 32'sd566941, -32'sd1065626, -32'sd821872, -32'sd1451502, -32'sd177255, 32'sd121895, 32'sd569597, -32'sd455335, -32'sd648136, 32'sd734463, 32'sd830479, -32'sd563342, -32'sd178919, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd562955, -32'sd776456, 32'sd198162, -32'sd1041753, 32'sd558163, -32'sd1385735, 32'sd247021, -32'sd464817, -32'sd1447001, -32'sd817562, 32'sd511695, -32'sd273136, -32'sd1114982, -32'sd541565, 32'sd690671, -32'sd45321, -32'sd2158763, 32'sd395821, -32'sd1631822, -32'sd523805, -32'sd400221, 32'sd831868, -32'sd177611, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd655171, 32'sd644117, 32'sd323788, 32'sd481183, -32'sd168190, -32'sd273952, 32'sd1136804, -32'sd38568, 32'sd316881, -32'sd788342, -32'sd314682, 32'sd1604295, -32'sd316755, 32'sd737389, -32'sd744119, -32'sd585978, 32'sd133296, -32'sd47057, -32'sd1160444, 32'sd611390, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd280330, -32'sd399496, -32'sd148443, -32'sd400397, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1009748, -32'sd1516603, -32'sd1318807, -32'sd1052894, -32'sd882321, 32'sd102605, -32'sd164699, -32'sd1889924, -32'sd571631, -32'sd1773801, -32'sd616582, -32'sd1669521, -32'sd263203, -32'sd969662, 32'sd835379, -32'sd545521, -32'sd1473072, -32'sd1051690, -32'sd500721, -32'sd889966, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd396982, -32'sd1378527, -32'sd628709, -32'sd845248, -32'sd329136, 32'sd836441, 32'sd183696, 32'sd387464, 32'sd349029, -32'sd353035, -32'sd1361347, -32'sd2195336, -32'sd3275566, -32'sd408235, -32'sd496343, -32'sd1385691, 32'sd774145, 32'sd2396313, 32'sd165584, -32'sd827979, -32'sd550376, -32'sd1886171, -32'sd1172313, 32'sd34518, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1312981, 32'sd729462, -32'sd1682956, 32'sd975372, 32'sd1005310, -32'sd1043392, -32'sd1442218, 32'sd100926, 32'sd370082, -32'sd1239614, -32'sd1552657, -32'sd1879689, 32'sd866626, 32'sd168917, -32'sd331269, 32'sd2390975, 32'sd1053053, 32'sd696534, 32'sd1856548, -32'sd424610, -32'sd891435, -32'sd604496, 32'sd1346092, 32'sd1359387, 32'sd1041844, 32'sd0, 32'sd0, -32'sd880561, 32'sd665694, -32'sd900367, -32'sd2005751, -32'sd405306, -32'sd372813, -32'sd2331003, -32'sd920524, -32'sd1606134, 32'sd485613, -32'sd2388452, -32'sd1371415, -32'sd956308, 32'sd582895, -32'sd959548, 32'sd795128, -32'sd821612, -32'sd238000, 32'sd578518, -32'sd358081, -32'sd595108, 32'sd1014910, 32'sd427158, 32'sd1230542, -32'sd279434, -32'sd278595, 32'sd804547, 32'sd0, -32'sd82645, -32'sd22700, 32'sd1351573, -32'sd2361325, 32'sd131111, -32'sd178981, -32'sd917960, -32'sd3148617, 32'sd684691, 32'sd57449, -32'sd924307, 32'sd106691, -32'sd2024849, -32'sd108028, 32'sd1385582, 32'sd2052679, 32'sd2413686, 32'sd641649, 32'sd903622, 32'sd470317, 32'sd2379481, 32'sd1938941, -32'sd56865, 32'sd422685, -32'sd681527, 32'sd6358, 32'sd625389, 32'sd0, 32'sd736447, 32'sd565315, 32'sd1187349, -32'sd2068324, 32'sd589124, -32'sd1323054, -32'sd1981561, 32'sd412111, -32'sd592737, -32'sd1823019, -32'sd1701978, -32'sd1210337, -32'sd1000108, -32'sd237271, 32'sd1887938, -32'sd172698, 32'sd189631, -32'sd408299, 32'sd421308, 32'sd1396499, 32'sd839864, 32'sd979354, 32'sd1552210, 32'sd661325, 32'sd755009, -32'sd298287, -32'sd1088759, 32'sd290008, -32'sd273386, -32'sd706086, -32'sd461259, -32'sd1503587, -32'sd929335, -32'sd3179511, -32'sd274004, -32'sd1999334, -32'sd1015044, -32'sd1501976, -32'sd172232, -32'sd837561, -32'sd345694, 32'sd1197816, 32'sd1433394, 32'sd1027513, 32'sd771615, -32'sd2069233, 32'sd1011755, 32'sd1571164, -32'sd1146487, -32'sd1220454, -32'sd940772, 32'sd100492, -32'sd581310, -32'sd458187, 32'sd897668, -32'sd386105, -32'sd477658, -32'sd2429480, 32'sd236958, -32'sd2507480, -32'sd1808965, -32'sd2736395, -32'sd1526745, -32'sd402974, -32'sd1773034, 32'sd156737, 32'sd158630, -32'sd515890, 32'sd874039, 32'sd156289, -32'sd412110, -32'sd1649173, -32'sd1285967, -32'sd1161633, -32'sd644496, 32'sd273648, -32'sd262867, -32'sd1730638, -32'sd1908653, -32'sd2684400, -32'sd1776322, -32'sd1415508, 32'sd4881, -32'sd1039684, -32'sd2063485, 32'sd57935, 32'sd483681, -32'sd1569257, -32'sd679268, 32'sd114525, -32'sd85116, -32'sd2363950, -32'sd540760, -32'sd882944, 32'sd2073890, -32'sd1695584, -32'sd1810092, -32'sd1012192, 32'sd146429, -32'sd549974, 32'sd690938, -32'sd647664, -32'sd727415, -32'sd2792884, 32'sd711159, -32'sd2294489, -32'sd991179, -32'sd1173468, -32'sd1294647, -32'sd607319, -32'sd912861, -32'sd1148116, -32'sd1076560, -32'sd2028869, -32'sd426007, 32'sd1456583, 32'sd709094, -32'sd2803174, -32'sd440593, -32'sd2377424, -32'sd1758128, -32'sd648749, 32'sd1030130, 32'sd2141322, -32'sd849669, 32'sd2240976, 32'sd1427501, -32'sd1074801, 32'sd938481, 32'sd1033886, -32'sd1595107, -32'sd2151896, -32'sd2706014, -32'sd164577, -32'sd2540377, -32'sd1487864, 32'sd970222, -32'sd606842, -32'sd1041268, 32'sd384919, 32'sd276986, -32'sd528709, 32'sd669735, 32'sd1388143, -32'sd836710, -32'sd472719, -32'sd1343203, -32'sd3110532, -32'sd2281923, 32'sd589911, -32'sd614646, 32'sd1637800, 32'sd1579860, 32'sd3466438, 32'sd702440, 32'sd1388953, 32'sd572117, -32'sd1092332, -32'sd1182208, -32'sd3041939, -32'sd2118784, -32'sd2853542, -32'sd889113, -32'sd1222304, -32'sd1562812, 32'sd1065278, 32'sd1187838, 32'sd455674, 32'sd69319, -32'sd2801855, -32'sd1109418, -32'sd2780029, 32'sd469535, 32'sd1299648, -32'sd2596046, -32'sd2105882, -32'sd1210056, 32'sd1440179, 32'sd1249641, 32'sd2128247, 32'sd2668095, 32'sd2400840, 32'sd956037, 32'sd2389632, 32'sd533663, -32'sd561974, -32'sd443505, 32'sd1108052, -32'sd2939559, -32'sd962321, 32'sd873039, 32'sd331598, 32'sd702317, -32'sd24614, -32'sd612202, -32'sd455248, -32'sd542193, -32'sd2023774, -32'sd360355, -32'sd3346008, -32'sd753746, 32'sd657897, 32'sd481672, -32'sd2696007, 32'sd1548495, -32'sd25593, -32'sd21520, 32'sd2551963, 32'sd2089660, 32'sd2275558, 32'sd1429737, 32'sd2138227, 32'sd2190395, -32'sd134766, -32'sd20768, -32'sd293707, -32'sd2296051, -32'sd2431059, -32'sd1747503, -32'sd791089, -32'sd456100, 32'sd62585, -32'sd1026728, -32'sd1129226, -32'sd1484623, -32'sd268471, -32'sd1469682, -32'sd2538435, -32'sd2208956, -32'sd842323, -32'sd1761268, 32'sd1080953, 32'sd1938989, 32'sd175660, 32'sd344314, 32'sd1634672, 32'sd2148953, 32'sd1753294, -32'sd519455, 32'sd1618997, 32'sd2274233, -32'sd1273127, -32'sd605645, -32'sd443712, -32'sd768599, -32'sd297788, -32'sd2768346, -32'sd1806751, -32'sd328276, -32'sd293125, 32'sd175639, -32'sd862056, -32'sd1052321, -32'sd389987, -32'sd622612, -32'sd880429, -32'sd100661, -32'sd1087443, 32'sd96004, 32'sd109446, -32'sd776902, -32'sd2991246, -32'sd2505288, 32'sd966407, 32'sd143812, 32'sd638766, 32'sd181, 32'sd1249087, 32'sd1671027, -32'sd317152, 32'sd1562591, 32'sd1504608, 32'sd1313468, 32'sd436136, -32'sd1274042, -32'sd1212161, -32'sd1610569, -32'sd1616519, -32'sd824600, 32'sd194375, -32'sd1361930, -32'sd732162, 32'sd1385273, -32'sd411158, 32'sd871822, -32'sd2234303, -32'sd1949133, 32'sd271312, -32'sd993695, -32'sd303620, -32'sd823734, 32'sd145903, 32'sd19651, 32'sd1008315, 32'sd3022539, 32'sd1640401, -32'sd804550, 32'sd45322, 32'sd1856486, 32'sd374724, -32'sd821515, -32'sd177570, 32'sd1171817, -32'sd751492, -32'sd1643882, -32'sd171945, -32'sd1490340, 32'sd0, -32'sd452110, -32'sd937760, -32'sd113122, 32'sd919528, 32'sd153231, -32'sd569473, 32'sd963096, -32'sd798205, -32'sd756515, -32'sd1022315, -32'sd575357, -32'sd392569, -32'sd798446, -32'sd117978, 32'sd1400648, 32'sd1147, 32'sd2808722, 32'sd1546578, -32'sd357779, 32'sd708906, 32'sd304345, 32'sd354565, 32'sd234135, 32'sd201266, -32'sd1233324, 32'sd1040172, 32'sd290657, -32'sd465433, -32'sd1187271, 32'sd1121712, 32'sd399528, -32'sd998567, 32'sd320591, -32'sd1093699, 32'sd130127, 32'sd1643451, -32'sd464791, -32'sd828961, 32'sd630048, -32'sd856890, -32'sd663151, -32'sd1108430, 32'sd185439, 32'sd629908, 32'sd2391368, 32'sd1746027, 32'sd1893615, -32'sd763920, -32'sd1440496, -32'sd1914439, -32'sd1157872, -32'sd962307, -32'sd2188382, 32'sd90330, 32'sd880977, -32'sd668650, -32'sd1177624, 32'sd363700, -32'sd380137, 32'sd405355, -32'sd49059, -32'sd1037495, 32'sd1916884, 32'sd905191, -32'sd278978, 32'sd149167, 32'sd688892, -32'sd836364, -32'sd832598, -32'sd1429553, -32'sd2025802, 32'sd2306046, 32'sd610366, 32'sd498018, 32'sd1863982, -32'sd1307900, -32'sd1370986, -32'sd757514, -32'sd841350, -32'sd1241463, -32'sd2128947, 32'sd1201525, -32'sd700403, 32'sd0, -32'sd360393, -32'sd477325, 32'sd1068298, -32'sd1056475, -32'sd886169, 32'sd1952394, 32'sd704194, -32'sd1307998, 32'sd96365, -32'sd832635, -32'sd214512, -32'sd1146017, 32'sd303236, -32'sd1554524, 32'sd1754422, 32'sd1960050, 32'sd628872, 32'sd2047152, 32'sd1634460, -32'sd647160, -32'sd575609, -32'sd422923, -32'sd1440478, 32'sd428724, -32'sd405691, 32'sd634921, -32'sd703297, -32'sd703674, -32'sd1103843, 32'sd213509, 32'sd813257, 32'sd506865, 32'sd1540535, 32'sd1955224, 32'sd578478, -32'sd1702841, 32'sd1205102, -32'sd938624, -32'sd1039889, -32'sd193251, -32'sd1117738, 32'sd445193, -32'sd243867, 32'sd1737272, 32'sd201774, -32'sd926696, -32'sd1209177, -32'sd1513527, -32'sd3476911, -32'sd2661393, 32'sd482967, -32'sd1126466, -32'sd854854, 32'sd519842, 32'sd18102, -32'sd951543, -32'sd1520330, 32'sd835603, -32'sd1334111, -32'sd877191, -32'sd1001409, -32'sd1034022, 32'sd998566, 32'sd440371, -32'sd936551, -32'sd241322, -32'sd73296, 32'sd773247, 32'sd1407725, 32'sd1831382, 32'sd1756629, 32'sd1355640, -32'sd2580694, -32'sd208436, -32'sd1477531, -32'sd2784268, -32'sd3266748, -32'sd1430237, 32'sd707144, 32'sd164454, -32'sd438850, -32'sd49572, -32'sd1255607, 32'sd0, 32'sd61796, -32'sd690819, -32'sd562999, -32'sd473441, 32'sd13354, -32'sd48918, 32'sd263320, -32'sd125155, -32'sd958067, 32'sd518823, -32'sd200377, 32'sd79028, 32'sd1410624, 32'sd1552577, 32'sd2489255, 32'sd112730, -32'sd2078026, 32'sd1392239, -32'sd130403, -32'sd3024547, -32'sd2142421, -32'sd1087659, -32'sd102871, -32'sd918699, -32'sd311367, 32'sd229821, 32'sd0, 32'sd0, 32'sd0, 32'sd52289, -32'sd990992, -32'sd1525416, 32'sd2268468, 32'sd1199606, -32'sd389697, -32'sd918383, 32'sd790862, 32'sd243239, 32'sd524629, 32'sd558532, -32'sd87284, 32'sd37546, 32'sd475722, 32'sd2347111, -32'sd594128, -32'sd540855, -32'sd4092176, -32'sd1168378, 32'sd259207, 32'sd2123265, 32'sd1866460, 32'sd1188169, -32'sd2720423, -32'sd948694, 32'sd0, 32'sd0, 32'sd0, 32'sd672126, -32'sd1040156, -32'sd943846, -32'sd529314, -32'sd157079, 32'sd49007, 32'sd71370, -32'sd189557, -32'sd1068209, -32'sd101920, -32'sd1545754, -32'sd3069546, -32'sd1198560, -32'sd578229, -32'sd1103570, -32'sd2893512, -32'sd1965863, -32'sd2806680, -32'sd1194385, 32'sd656375, 32'sd1107216, 32'sd131288, 32'sd821549, 32'sd241890, -32'sd1291775, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd80747, -32'sd1763801, -32'sd1223741, 32'sd657042, 32'sd1506177, 32'sd897335, -32'sd1750586, -32'sd262567, 32'sd965983, -32'sd2113760, -32'sd1922813, -32'sd1972361, -32'sd618257, 32'sd1697765, 32'sd208970, -32'sd1753722, -32'sd1534703, -32'sd1417500, 32'sd680442, -32'sd1524362, -32'sd449246, -32'sd500440, -32'sd1165094, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd465584, -32'sd442579, -32'sd1822824, -32'sd128165, 32'sd967990, -32'sd225089, -32'sd1264459, -32'sd2117048, 32'sd988388, -32'sd1589949, 32'sd295389, 32'sd1231955, 32'sd1327012, 32'sd331945, -32'sd1236683, -32'sd1648810, -32'sd1547457, -32'sd663415, 32'sd102576, -32'sd983791, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1634844, 32'sd995884, 32'sd2013243, 32'sd1658204, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2203483, 32'sd2026066, -32'sd49484, 32'sd1572806, 32'sd1719945, 32'sd1062137, 32'sd1816671, 32'sd469889, 32'sd2009560, 32'sd1415040, 32'sd597125, 32'sd325201, 32'sd580457, 32'sd892735, 32'sd1954663, -32'sd588811, 32'sd1315348, 32'sd550690, 32'sd2698617, 32'sd2006860, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2450659, -32'sd162751, 32'sd401002, -32'sd290756, -32'sd1791297, -32'sd801025, 32'sd137061, -32'sd2144180, 32'sd168132, 32'sd166322, -32'sd37668, -32'sd942580, -32'sd11787, 32'sd1263675, -32'sd281214, 32'sd904117, -32'sd559317, 32'sd359402, -32'sd60568, -32'sd858509, -32'sd57870, 32'sd879875, -32'sd734521, 32'sd2635371, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1494420, 32'sd432679, -32'sd1098248, 32'sd1019169, -32'sd98698, -32'sd1115380, 32'sd1421998, -32'sd1567882, 32'sd446887, 32'sd447315, 32'sd755000, 32'sd772632, 32'sd935860, 32'sd2063023, 32'sd476985, -32'sd45310, 32'sd913249, 32'sd545414, 32'sd1638897, -32'sd221920, 32'sd763811, -32'sd1175026, 32'sd395795, 32'sd1625292, -32'sd160957, 32'sd0, 32'sd0, 32'sd2083449, -32'sd922514, 32'sd255967, 32'sd667175, 32'sd728798, -32'sd473058, -32'sd726525, 32'sd1634146, 32'sd315042, 32'sd1218017, 32'sd894314, 32'sd77250, 32'sd692069, 32'sd938354, 32'sd1069903, 32'sd359269, 32'sd127282, 32'sd1039508, 32'sd183351, 32'sd1495504, 32'sd365982, 32'sd981259, 32'sd1129698, 32'sd1240190, -32'sd1063536, -32'sd1075943, 32'sd1065881, 32'sd0, 32'sd1737304, 32'sd1082327, -32'sd190781, -32'sd1176584, -32'sd75525, 32'sd226482, -32'sd455845, 32'sd1591210, 32'sd1470271, -32'sd1381147, -32'sd1699076, -32'sd280547, -32'sd956735, -32'sd134555, -32'sd1405287, -32'sd532091, 32'sd758559, -32'sd1290797, -32'sd292611, -32'sd453410, 32'sd105905, -32'sd838235, -32'sd1314021, -32'sd534786, 32'sd229386, -32'sd1530353, 32'sd634937, 32'sd0, -32'sd269241, 32'sd150604, -32'sd1093089, -32'sd1467466, 32'sd844922, -32'sd32943, -32'sd1882104, -32'sd2192474, -32'sd924303, -32'sd1549193, -32'sd213115, -32'sd1615952, -32'sd1559234, -32'sd1082929, -32'sd2708077, -32'sd2014431, -32'sd2439452, -32'sd565312, -32'sd993048, 32'sd427140, 32'sd1270217, 32'sd1065391, -32'sd335258, -32'sd899293, 32'sd133647, -32'sd317456, -32'sd204792, 32'sd2284064, 32'sd1358467, -32'sd2040285, 32'sd671359, -32'sd1567641, -32'sd696207, 32'sd182417, 32'sd977383, -32'sd383294, -32'sd1155514, 32'sd56295, -32'sd2367370, -32'sd424320, -32'sd1606670, -32'sd2865468, -32'sd3533323, -32'sd1837493, -32'sd2358114, -32'sd2264687, -32'sd492947, -32'sd2838063, -32'sd1348067, -32'sd192697, 32'sd77328, -32'sd858111, 32'sd248562, -32'sd1584300, 32'sd340436, -32'sd288365, 32'sd354887, -32'sd1710645, 32'sd39657, -32'sd184594, 32'sd570993, 32'sd617271, -32'sd263260, 32'sd561277, 32'sd504928, 32'sd1584021, -32'sd1159036, 32'sd1092345, 32'sd774042, -32'sd1871000, 32'sd806092, 32'sd68381, -32'sd327257, -32'sd1027440, -32'sd391813, 32'sd807032, 32'sd500012, 32'sd534460, 32'sd69759, 32'sd1014720, 32'sd996049, 32'sd730253, 32'sd947603, 32'sd1528285, 32'sd70243, 32'sd248983, 32'sd844871, 32'sd1799873, 32'sd1989254, 32'sd1115445, 32'sd1120835, 32'sd2210794, 32'sd284860, 32'sd1719813, 32'sd1359890, 32'sd3135449, 32'sd1897778, 32'sd2520566, 32'sd2692533, 32'sd3302260, 32'sd2713309, 32'sd686861, 32'sd58650, 32'sd2222003, 32'sd2949592, 32'sd2174783, -32'sd24309, 32'sd1195173, 32'sd81320, 32'sd48900, -32'sd2151477, 32'sd1477916, 32'sd1547293, 32'sd2361069, -32'sd1236164, 32'sd983709, 32'sd205797, 32'sd93286, -32'sd415349, -32'sd1551203, 32'sd1388472, 32'sd1851351, 32'sd4670087, 32'sd2362098, 32'sd4286205, 32'sd2886922, 32'sd2690989, 32'sd2618886, 32'sd448804, 32'sd2895903, 32'sd2771993, 32'sd2973547, 32'sd4149009, 32'sd1867639, 32'sd1392130, 32'sd2622520, 32'sd331053, 32'sd116087, 32'sd1022937, 32'sd699690, 32'sd842093, 32'sd273760, 32'sd2581809, 32'sd768478, -32'sd1197038, -32'sd630755, 32'sd135163, 32'sd327214, 32'sd440544, 32'sd1368878, 32'sd3463802, 32'sd2789772, 32'sd1386936, 32'sd2975225, 32'sd2764090, -32'sd261466, 32'sd1473505, 32'sd2805329, 32'sd2750107, 32'sd1735806, -32'sd425486, 32'sd1374652, 32'sd1472592, 32'sd2192278, 32'sd1468186, -32'sd103301, -32'sd1548312, 32'sd2239707, -32'sd1007930, 32'sd1009260, -32'sd1291265, -32'sd1781727, -32'sd2119171, -32'sd1464628, -32'sd425520, 32'sd1116858, 32'sd667581, 32'sd1892968, 32'sd278620, -32'sd675637, -32'sd994077, -32'sd910483, -32'sd990823, 32'sd907839, -32'sd896881, -32'sd862116, 32'sd1107384, 32'sd184874, -32'sd903718, -32'sd137819, -32'sd1727052, -32'sd1834564, 32'sd277985, 32'sd1454702, 32'sd935761, 32'sd1871955, -32'sd20428, -32'sd450309, -32'sd1059000, -32'sd2809905, 32'sd259891, -32'sd989657, -32'sd123416, -32'sd654394, -32'sd973125, 32'sd191979, 32'sd422488, -32'sd1483492, -32'sd4139103, -32'sd1661559, -32'sd3552330, 32'sd527319, -32'sd255424, -32'sd2104773, -32'sd2325221, -32'sd2022732, -32'sd1894759, -32'sd3466569, -32'sd2194810, -32'sd2619084, -32'sd3483276, -32'sd1660967, 32'sd1732172, 32'sd2171906, 32'sd161793, 32'sd887745, -32'sd1559299, 32'sd127270, -32'sd1009574, -32'sd290360, -32'sd1863962, -32'sd1015252, -32'sd1468668, -32'sd620692, -32'sd1030562, -32'sd1054874, -32'sd3354740, -32'sd3805244, -32'sd872472, -32'sd679702, -32'sd2395948, -32'sd1012760, 32'sd360973, -32'sd406947, -32'sd1363229, -32'sd2505304, -32'sd2042270, -32'sd1180106, 32'sd2177044, -32'sd2723016, 32'sd1340268, 32'sd297158, -32'sd636493, -32'sd616029, -32'sd1126193, 32'sd890834, 32'sd1079555, 32'sd228699, -32'sd394248, -32'sd1517391, -32'sd1848951, 32'sd223897, -32'sd2566885, -32'sd1611427, -32'sd2211919, -32'sd1284601, -32'sd816079, -32'sd1607345, -32'sd1810731, -32'sd2453382, -32'sd319856, 32'sd417903, 32'sd998502, 32'sd1276316, 32'sd1019469, 32'sd1076994, 32'sd199971, 32'sd1274665, 32'sd286754, 32'sd1454517, -32'sd1082820, -32'sd455763, 32'sd1991842, 32'sd1403540, 32'sd1339335, 32'sd1350110, -32'sd123269, -32'sd1781739, -32'sd1220555, -32'sd2480048, -32'sd3061119, -32'sd1502358, -32'sd1252136, -32'sd2693340, -32'sd201305, -32'sd1682733, -32'sd788427, 32'sd509342, -32'sd68524, 32'sd2544837, 32'sd1998003, -32'sd1443277, -32'sd642953, 32'sd1136797, -32'sd844380, 32'sd565825, 32'sd368654, 32'sd0, 32'sd464732, -32'sd1600074, 32'sd93817, 32'sd1944697, 32'sd1906329, 32'sd1595161, -32'sd1124399, -32'sd1053193, 32'sd297966, -32'sd271977, 32'sd432121, -32'sd304777, -32'sd1864479, 32'sd107217, 32'sd137498, -32'sd178381, -32'sd718314, -32'sd123545, -32'sd2236840, 32'sd1539085, 32'sd1737344, -32'sd2922265, -32'sd1063901, 32'sd1024303, -32'sd229272, 32'sd669026, -32'sd36406, 32'sd360709, 32'sd676316, -32'sd349063, 32'sd173310, 32'sd969505, 32'sd2079272, 32'sd51569, -32'sd75404, 32'sd1087725, 32'sd76378, 32'sd1941786, 32'sd984939, 32'sd1712842, 32'sd1089541, -32'sd850610, -32'sd794808, 32'sd221849, 32'sd1208391, 32'sd636011, -32'sd1060287, 32'sd330652, 32'sd423495, -32'sd1656449, -32'sd1064242, 32'sd517478, -32'sd760011, 32'sd804349, -32'sd262394, 32'sd2147608, 32'sd772784, 32'sd1334179, 32'sd1895818, 32'sd1187697, 32'sd1209335, 32'sd1751438, 32'sd1502870, 32'sd2323610, 32'sd1220442, -32'sd335934, 32'sd1009157, 32'sd1110903, 32'sd1135757, -32'sd51451, 32'sd389707, 32'sd338551, 32'sd43772, -32'sd1568141, 32'sd956452, -32'sd723752, -32'sd1727524, -32'sd4023549, -32'sd1181436, 32'sd433006, 32'sd1138597, -32'sd1006267, -32'sd226539, 32'sd0, -32'sd7642, -32'sd182610, -32'sd136077, -32'sd713799, -32'sd191424, 32'sd279233, -32'sd642892, -32'sd380227, 32'sd1445504, 32'sd1961619, 32'sd527382, 32'sd79671, 32'sd1001089, 32'sd1643475, -32'sd1116566, 32'sd1063589, -32'sd850482, -32'sd849020, -32'sd1330453, -32'sd433725, -32'sd2781748, -32'sd3094765, -32'sd1313488, -32'sd1050081, -32'sd338959, -32'sd892869, 32'sd909855, 32'sd1479758, 32'sd1295413, -32'sd2321086, -32'sd1039774, -32'sd938866, -32'sd498, -32'sd268885, -32'sd856651, 32'sd500076, 32'sd1122769, 32'sd488471, -32'sd159626, 32'sd929755, -32'sd377360, -32'sd1036188, 32'sd282690, -32'sd105473, 32'sd844645, 32'sd1747159, 32'sd356034, -32'sd2561215, -32'sd2630715, -32'sd1993811, 32'sd212007, -32'sd803282, -32'sd227951, -32'sd2294616, 32'sd591812, 32'sd1272307, 32'sd2083781, -32'sd1049197, -32'sd1466913, -32'sd275041, 32'sd1248784, -32'sd793792, -32'sd384171, -32'sd1909790, 32'sd524216, 32'sd152625, -32'sd22870, 32'sd828758, -32'sd510864, -32'sd242567, 32'sd43777, 32'sd696066, 32'sd191774, 32'sd574773, -32'sd684292, -32'sd2745542, -32'sd690331, -32'sd1749493, 32'sd19075, -32'sd1031596, -32'sd601598, 32'sd1002337, 32'sd1325406, 32'sd0, 32'sd2362795, 32'sd822232, -32'sd99673, 32'sd1561791, 32'sd288468, -32'sd664362, -32'sd695870, -32'sd249698, 32'sd271843, 32'sd647616, -32'sd377834, 32'sd1119477, 32'sd351407, 32'sd1944594, 32'sd1500164, -32'sd446189, -32'sd1557707, -32'sd218998, 32'sd383171, -32'sd428808, 32'sd1349, 32'sd378317, 32'sd844291, 32'sd215664, 32'sd826849, -32'sd672404, 32'sd0, 32'sd0, 32'sd0, 32'sd926954, 32'sd86689, -32'sd213334, 32'sd632130, -32'sd451400, 32'sd564196, -32'sd76982, -32'sd43416, -32'sd555960, -32'sd510831, -32'sd597057, 32'sd828864, 32'sd749300, 32'sd606874, -32'sd700909, 32'sd1253018, -32'sd520172, -32'sd656473, -32'sd1356395, 32'sd361603, -32'sd341329, -32'sd1299801, 32'sd810617, 32'sd828327, -32'sd1559543, 32'sd0, 32'sd0, 32'sd0, 32'sd2267896, 32'sd1464348, 32'sd647822, -32'sd1382843, 32'sd278024, -32'sd341304, -32'sd717537, -32'sd57058, 32'sd1184364, -32'sd1779073, -32'sd147833, 32'sd1031184, -32'sd131138, -32'sd1111810, 32'sd1400580, 32'sd1046407, 32'sd1290231, 32'sd1108773, -32'sd184405, -32'sd1004607, -32'sd341041, -32'sd1555358, 32'sd915610, 32'sd2432266, 32'sd1390248, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2394790, 32'sd701661, 32'sd789931, 32'sd995878, 32'sd405093, -32'sd666885, -32'sd399769, 32'sd209548, -32'sd520340, 32'sd905393, 32'sd85457, 32'sd2319925, 32'sd713176, 32'sd402490, 32'sd359586, 32'sd660522, 32'sd427519, 32'sd648486, 32'sd483593, 32'sd92116, 32'sd551364, -32'sd145891, 32'sd2562671, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2434426, 32'sd1270704, 32'sd737537, 32'sd1163527, 32'sd1142303, 32'sd583304, 32'sd340395, 32'sd499781, 32'sd198882, 32'sd800383, 32'sd478298, 32'sd480351, 32'sd1445596, 32'sd154457, 32'sd276683, -32'sd727849, 32'sd699134, -32'sd173639, -32'sd1149049, 32'sd2029152, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1678550, 32'sd603117, 32'sd1485006, 32'sd485609, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd601806, 32'sd1344885, -32'sd1114090, 32'sd1450873, 32'sd648261, 32'sd21034, 32'sd1635417, -32'sd640267, 32'sd1210869, 32'sd863443, 32'sd2033609, 32'sd1339543, 32'sd1327605, 32'sd898004, 32'sd1494061, 32'sd117688, 32'sd943894, -32'sd178043, 32'sd605808, 32'sd358348, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd363026, 32'sd469931, 32'sd1922337, -32'sd105191, -32'sd582798, -32'sd136903, 32'sd999796, 32'sd994677, 32'sd1634772, 32'sd1020356, 32'sd374743, 32'sd2328930, 32'sd888607, 32'sd747647, 32'sd1036654, 32'sd595031, 32'sd249944, -32'sd982326, 32'sd1923252, 32'sd1570484, 32'sd1382718, -32'sd1504010, 32'sd1068946, 32'sd1592351, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1107992, 32'sd1879787, 32'sd68328, 32'sd1433774, 32'sd1221571, -32'sd618990, 32'sd1874706, 32'sd447108, -32'sd765039, 32'sd2839203, 32'sd2719982, 32'sd1914981, -32'sd1947646, -32'sd1933768, 32'sd725380, 32'sd1295196, -32'sd309179, -32'sd238267, -32'sd822991, -32'sd399650, 32'sd672809, -32'sd1448870, 32'sd3328, -32'sd631167, 32'sd151985, 32'sd0, 32'sd0, -32'sd86286, -32'sd487614, -32'sd1153692, 32'sd1006120, -32'sd188952, -32'sd159056, -32'sd66078, 32'sd893661, -32'sd1419221, -32'sd365757, 32'sd295107, 32'sd1415922, 32'sd81478, -32'sd248676, 32'sd496360, -32'sd664635, -32'sd930987, -32'sd677939, 32'sd898542, 32'sd617828, -32'sd1743973, -32'sd1194590, 32'sd901976, 32'sd972563, 32'sd888557, -32'sd2294795, 32'sd446276, 32'sd0, 32'sd130317, 32'sd1028380, 32'sd784352, 32'sd371835, -32'sd457402, -32'sd8938, -32'sd53792, 32'sd561751, -32'sd522231, 32'sd576806, -32'sd659270, 32'sd1021136, 32'sd3143, -32'sd848830, 32'sd77354, -32'sd67432, -32'sd562129, -32'sd2597187, -32'sd2730182, -32'sd1861082, 32'sd29217, -32'sd2533507, 32'sd895523, 32'sd1603374, 32'sd1418522, -32'sd431555, 32'sd793707, 32'sd0, -32'sd531380, 32'sd751020, 32'sd1414057, 32'sd942198, -32'sd993915, -32'sd333038, 32'sd1724315, 32'sd1151411, 32'sd780443, 32'sd378795, 32'sd783238, 32'sd1487481, -32'sd933868, -32'sd1382654, -32'sd3815041, -32'sd1655228, 32'sd199936, -32'sd1312507, -32'sd290612, -32'sd1990825, -32'sd1448800, -32'sd1810962, -32'sd222940, 32'sd702185, 32'sd537763, 32'sd96595, -32'sd455812, 32'sd723751, 32'sd1376874, 32'sd828263, -32'sd678628, 32'sd1459115, 32'sd523921, -32'sd451773, 32'sd768391, 32'sd164571, 32'sd1184697, 32'sd1674966, 32'sd57582, -32'sd666940, -32'sd1636234, -32'sd2130102, 32'sd86844, -32'sd356788, -32'sd1661794, 32'sd1568976, 32'sd1741938, 32'sd157798, 32'sd296705, 32'sd654803, -32'sd1606374, -32'sd1317153, -32'sd1845442, 32'sd90928, 32'sd455783, 32'sd416100, 32'sd1025518, 32'sd710961, 32'sd292854, 32'sd1524495, -32'sd1494671, 32'sd1117708, 32'sd2342880, 32'sd656146, 32'sd2464670, 32'sd2388637, 32'sd3182077, 32'sd180896, -32'sd3596901, -32'sd2347749, 32'sd276029, 32'sd1620606, -32'sd1390110, 32'sd1305982, -32'sd925830, 32'sd1263487, 32'sd1060640, 32'sd1957927, -32'sd413429, 32'sd562778, -32'sd243593, -32'sd1347413, 32'sd161734, 32'sd262703, -32'sd956313, -32'sd1214792, 32'sd824393, 32'sd1401869, 32'sd205137, 32'sd1187960, 32'sd1442282, 32'sd2165777, 32'sd801351, 32'sd365375, 32'sd575631, -32'sd2176053, -32'sd3224978, -32'sd1611353, -32'sd1246537, 32'sd650702, 32'sd1020119, 32'sd2732898, 32'sd159044, 32'sd2428238, 32'sd1976483, 32'sd675063, -32'sd87280, 32'sd1402677, 32'sd1734656, -32'sd588295, -32'sd1616836, 32'sd1654848, -32'sd840145, -32'sd45301, -32'sd706545, 32'sd2784159, 32'sd2027772, -32'sd4804, 32'sd274252, 32'sd1453288, -32'sd592930, 32'sd1138688, 32'sd896268, -32'sd1045680, -32'sd1087386, -32'sd2113282, -32'sd863974, 32'sd1730904, 32'sd563, 32'sd3980735, 32'sd2021190, 32'sd709914, -32'sd530991, 32'sd852040, 32'sd1483149, 32'sd2702530, 32'sd1474667, -32'sd406543, 32'sd134644, -32'sd68196, -32'sd575002, 32'sd1546317, 32'sd1572221, -32'sd331302, 32'sd1657413, 32'sd1475050, 32'sd859824, 32'sd2039808, 32'sd3629518, 32'sd705250, -32'sd10151, -32'sd1653616, -32'sd2852608, -32'sd2545442, 32'sd413643, 32'sd1420637, 32'sd1580708, 32'sd2397073, -32'sd75616, 32'sd325894, -32'sd1250952, 32'sd1793665, 32'sd1051529, 32'sd2300429, 32'sd568558, -32'sd1577861, -32'sd1060272, 32'sd1229934, 32'sd636188, 32'sd1089170, -32'sd1373690, -32'sd398437, 32'sd1357817, -32'sd1458003, 32'sd1519566, 32'sd3896087, 32'sd2266684, 32'sd510127, -32'sd956228, -32'sd2390320, -32'sd1515163, -32'sd2233928, -32'sd2060499, -32'sd1264909, 32'sd1519744, 32'sd22193, -32'sd436759, 32'sd329729, 32'sd262980, 32'sd258839, 32'sd633357, 32'sd2721821, 32'sd29540, -32'sd1348685, -32'sd55762, 32'sd489058, -32'sd556644, -32'sd1317949, -32'sd172849, -32'sd245571, 32'sd1790565, 32'sd1862449, 32'sd2677593, 32'sd1722300, 32'sd2453563, 32'sd1949932, -32'sd1620161, -32'sd3151742, -32'sd2559989, -32'sd3111653, -32'sd2048708, -32'sd1256523, 32'sd1522425, 32'sd681556, 32'sd73271, 32'sd796017, 32'sd1395185, -32'sd51484, 32'sd1377813, 32'sd668313, 32'sd349525, 32'sd473590, 32'sd889104, -32'sd350970, -32'sd122410, 32'sd276869, 32'sd763834, -32'sd215755, -32'sd304666, 32'sd1079499, 32'sd1999134, 32'sd656001, 32'sd701712, -32'sd48147, 32'sd591551, -32'sd1761220, -32'sd2795120, -32'sd3076586, -32'sd3270420, 32'sd2773884, 32'sd2391549, 32'sd2908633, 32'sd636094, 32'sd1222929, 32'sd1886134, 32'sd1633612, 32'sd1130346, -32'sd866785, 32'sd844653, 32'sd102586, 32'sd674850, 32'sd475702, -32'sd870412, -32'sd2616095, 32'sd1124921, -32'sd353961, -32'sd394917, 32'sd40284, 32'sd2553750, 32'sd1686537, -32'sd222364, -32'sd1247276, -32'sd581863, -32'sd2192457, -32'sd1428224, -32'sd3364207, -32'sd198058, 32'sd590229, 32'sd1762341, 32'sd1028939, 32'sd825139, 32'sd1018602, -32'sd442161, 32'sd1349101, 32'sd1740036, -32'sd1589971, 32'sd1645499, -32'sd943052, 32'sd121299, 32'sd576922, 32'sd614266, -32'sd1179384, 32'sd921430, 32'sd535524, 32'sd1675291, 32'sd989482, 32'sd1579571, 32'sd1705651, -32'sd1925274, 32'sd34465, -32'sd646418, -32'sd565053, -32'sd2430562, -32'sd1959557, -32'sd81536, 32'sd1142254, 32'sd4458338, 32'sd2128781, 32'sd503796, 32'sd1331503, 32'sd1001949, -32'sd920950, 32'sd837060, -32'sd495805, 32'sd639267, 32'sd418240, -32'sd432931, 32'sd0, 32'sd83335, 32'sd1200509, -32'sd105393, 32'sd460022, 32'sd533595, 32'sd282892, 32'sd1107314, 32'sd531068, 32'sd1066620, -32'sd775622, -32'sd1131768, -32'sd2553046, -32'sd3495027, 32'sd745460, 32'sd163470, 32'sd4021104, 32'sd3083716, 32'sd1712938, -32'sd339298, -32'sd2178379, -32'sd193744, 32'sd1776581, 32'sd301779, -32'sd171588, -32'sd469404, -32'sd647278, -32'sd94677, 32'sd114689, -32'sd1339350, 32'sd1586107, -32'sd2197767, -32'sd225810, 32'sd139275, -32'sd764406, -32'sd163257, -32'sd142231, 32'sd1665303, -32'sd285283, -32'sd2283427, -32'sd4514728, -32'sd792877, 32'sd391942, 32'sd2234846, 32'sd3525286, 32'sd2306816, 32'sd1408957, -32'sd1717120, -32'sd1985418, -32'sd1264995, 32'sd696060, -32'sd959149, 32'sd1378421, 32'sd1433813, 32'sd462944, 32'sd573161, 32'sd716189, 32'sd1461385, -32'sd401200, -32'sd1512057, -32'sd1371407, -32'sd450663, 32'sd88980, 32'sd1464421, 32'sd900759, 32'sd1100406, 32'sd570814, -32'sd1535459, -32'sd4838505, -32'sd3467582, 32'sd345898, 32'sd2542347, 32'sd3609120, 32'sd1395492, 32'sd1238183, 32'sd1331395, 32'sd554778, -32'sd2262545, 32'sd625274, 32'sd670378, 32'sd833713, 32'sd601079, -32'sd216663, -32'sd1505694, 32'sd0, -32'sd125828, 32'sd1856138, -32'sd340324, -32'sd1174012, 32'sd1688330, -32'sd609391, -32'sd126600, 32'sd1842347, 32'sd966002, -32'sd906949, -32'sd2077514, -32'sd1907129, -32'sd2390236, 32'sd638728, 32'sd3457270, 32'sd3643903, -32'sd818876, 32'sd1170186, 32'sd509146, -32'sd1249239, -32'sd1878630, -32'sd528415, -32'sd1535198, 32'sd1171518, 32'sd1193348, -32'sd2089151, -32'sd305794, 32'sd588120, 32'sd330488, -32'sd638633, -32'sd1599606, -32'sd2123864, 32'sd1552362, -32'sd1070038, -32'sd953942, 32'sd1050353, 32'sd737210, 32'sd1933385, 32'sd149378, -32'sd1796643, -32'sd983601, 32'sd922948, 32'sd2843287, 32'sd2286764, 32'sd2137214, -32'sd476096, -32'sd700012, -32'sd1179204, -32'sd1193337, 32'sd117300, -32'sd134020, 32'sd608371, -32'sd643005, -32'sd101595, 32'sd1402924, 32'sd160381, -32'sd241391, -32'sd603246, 32'sd341708, -32'sd1206761, 32'sd1475242, 32'sd668398, 32'sd422387, -32'sd236814, 32'sd1497990, -32'sd1344350, -32'sd1019087, -32'sd2768275, -32'sd961679, 32'sd623929, 32'sd3557890, 32'sd2489081, 32'sd1626050, -32'sd1941848, 32'sd302047, 32'sd521565, 32'sd161148, 32'sd66204, -32'sd3359882, -32'sd1053326, -32'sd920676, -32'sd1574773, -32'sd451347, 32'sd0, 32'sd1113610, -32'sd1127658, 32'sd188039, -32'sd952402, 32'sd63153, 32'sd1306372, 32'sd959000, 32'sd2514540, 32'sd295172, -32'sd586270, -32'sd3641760, -32'sd2374029, -32'sd465916, 32'sd3029744, 32'sd2145369, 32'sd2674303, 32'sd2181115, -32'sd2285769, -32'sd1595745, -32'sd365255, 32'sd509095, -32'sd1765669, 32'sd350182, -32'sd280064, 32'sd600842, -32'sd65687, 32'sd0, 32'sd0, 32'sd0, 32'sd562329, -32'sd96769, 32'sd151867, -32'sd767774, -32'sd525281, 32'sd415133, 32'sd869799, 32'sd1559173, -32'sd1510473, -32'sd3274805, -32'sd3056725, -32'sd1574350, -32'sd535702, 32'sd310145, 32'sd365833, 32'sd786152, -32'sd343873, -32'sd18994, 32'sd1957582, -32'sd542940, -32'sd767705, -32'sd95353, -32'sd1793773, 32'sd27618, 32'sd683266, 32'sd0, 32'sd0, 32'sd0, -32'sd863134, -32'sd316253, -32'sd1632248, -32'sd244390, 32'sd1180644, 32'sd1262316, -32'sd222837, 32'sd565748, -32'sd2264341, -32'sd2641719, -32'sd726039, -32'sd1073175, 32'sd742275, 32'sd565955, 32'sd2061860, 32'sd2137687, 32'sd508691, -32'sd400545, 32'sd529738, 32'sd2435642, -32'sd476604, -32'sd876085, 32'sd865869, 32'sd980361, -32'sd115467, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd309219, -32'sd624734, 32'sd148069, 32'sd725588, 32'sd1255634, 32'sd618755, -32'sd509154, -32'sd1672076, 32'sd178621, 32'sd245787, 32'sd399458, 32'sd1156046, 32'sd657543, 32'sd880562, -32'sd545672, -32'sd888679, 32'sd431142, -32'sd1512420, 32'sd1250726, 32'sd1382730, 32'sd799133, -32'sd287429, -32'sd292846, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1436089, 32'sd846511, 32'sd301394, 32'sd1120878, 32'sd270963, 32'sd178769, -32'sd1766410, 32'sd811377, -32'sd958436, 32'sd1145879, 32'sd726773, -32'sd797683, 32'sd783803, 32'sd180443, 32'sd1394483, -32'sd356885, -32'sd1153925, -32'sd35881, 32'sd144261, -32'sd1194552, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd604999, -32'sd705179, 32'sd68369, -32'sd603146, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd762526, 32'sd1341641, 32'sd1054512, -32'sd1718090, 32'sd894511, 32'sd401505, 32'sd234761, 32'sd1066352, -32'sd1165976, -32'sd864305, 32'sd620672, 32'sd1009700, -32'sd434028, 32'sd129183, -32'sd199920, -32'sd267212, 32'sd338271, 32'sd855045, 32'sd483895, 32'sd654516, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1610807, 32'sd539898, -32'sd809180, 32'sd1138850, 32'sd351420, -32'sd864359, 32'sd307644, -32'sd368472, -32'sd262154, 32'sd1262938, 32'sd1907453, 32'sd2606387, -32'sd1163640, 32'sd803350, 32'sd1895258, -32'sd1628981, -32'sd581417, 32'sd1723800, 32'sd993192, -32'sd1041435, 32'sd333854, 32'sd427471, 32'sd954607, 32'sd439177, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1643818, -32'sd470873, 32'sd547388, -32'sd319292, 32'sd1340574, -32'sd704199, -32'sd170305, 32'sd682533, 32'sd2238552, 32'sd991601, 32'sd3545819, 32'sd2538362, 32'sd453615, 32'sd757504, 32'sd2007780, -32'sd842436, -32'sd1910606, -32'sd2147777, 32'sd1142458, 32'sd389917, -32'sd287756, -32'sd875421, 32'sd687285, -32'sd479064, 32'sd727120, 32'sd0, 32'sd0, 32'sd911712, -32'sd1035940, -32'sd787603, -32'sd463622, 32'sd974633, -32'sd883351, -32'sd1404458, -32'sd1001967, 32'sd2770533, 32'sd1275151, 32'sd1465763, 32'sd2790185, 32'sd672428, 32'sd1246535, 32'sd909023, -32'sd724053, 32'sd575709, -32'sd686648, -32'sd1805715, -32'sd222163, 32'sd939558, 32'sd1202434, -32'sd1644472, -32'sd821778, -32'sd1584547, -32'sd126550, 32'sd474147, 32'sd0, 32'sd470377, 32'sd304234, -32'sd348427, 32'sd255527, -32'sd895492, 32'sd633690, -32'sd626384, 32'sd870663, 32'sd213346, 32'sd1223046, 32'sd1536618, -32'sd121416, 32'sd1138217, 32'sd2524134, 32'sd1416652, 32'sd50278, -32'sd169375, 32'sd1305832, 32'sd425954, -32'sd179139, -32'sd514301, 32'sd913864, -32'sd624098, 32'sd91271, 32'sd535652, -32'sd1488755, 32'sd173360, 32'sd0, 32'sd934762, 32'sd486113, 32'sd1758239, -32'sd700173, -32'sd20516, -32'sd796715, -32'sd1333377, 32'sd621219, -32'sd443617, 32'sd956503, -32'sd686617, 32'sd1108025, 32'sd748669, 32'sd861829, 32'sd2199501, 32'sd2004574, -32'sd75834, 32'sd1430897, -32'sd472889, -32'sd369585, 32'sd324024, -32'sd580269, -32'sd1572083, 32'sd648204, 32'sd2356960, 32'sd471487, -32'sd578714, 32'sd1019273, 32'sd1014982, 32'sd1010901, 32'sd1743444, -32'sd1054171, -32'sd139069, -32'sd1044616, -32'sd1014930, -32'sd1686431, 32'sd275919, -32'sd74797, 32'sd1630123, 32'sd1492213, 32'sd940454, 32'sd779659, 32'sd1522498, 32'sd2682288, 32'sd2692972, 32'sd194043, 32'sd3076177, 32'sd1024874, -32'sd433750, -32'sd522650, 32'sd230994, 32'sd910368, -32'sd251910, -32'sd621485, 32'sd579951, 32'sd984704, 32'sd976661, 32'sd485228, -32'sd1579043, -32'sd509300, 32'sd1202758, -32'sd882094, -32'sd885794, -32'sd219396, -32'sd1748681, 32'sd433616, 32'sd326357, 32'sd764152, 32'sd2193752, 32'sd2044687, 32'sd1769036, 32'sd1521414, 32'sd1835981, 32'sd1958619, -32'sd51319, 32'sd2417436, 32'sd1632947, 32'sd1852737, 32'sd764381, 32'sd552612, 32'sd230011, -32'sd153535, -32'sd1406781, 32'sd1085462, -32'sd1269320, -32'sd1914847, -32'sd48338, 32'sd77054, -32'sd1394557, -32'sd2149656, -32'sd72068, -32'sd318816, -32'sd378136, -32'sd1268526, -32'sd16069, 32'sd388742, 32'sd1923787, 32'sd2490397, 32'sd1744729, 32'sd1513452, -32'sd1672311, -32'sd1452235, 32'sd41111, 32'sd776738, 32'sd592518, 32'sd628245, 32'sd886889, 32'sd1742743, 32'sd1658928, -32'sd405288, 32'sd783594, -32'sd627511, 32'sd11933, -32'sd1239766, -32'sd2984131, -32'sd36885, -32'sd1134766, -32'sd906591, -32'sd1687480, -32'sd706796, 32'sd1031607, -32'sd1439830, 32'sd502534, 32'sd1419517, 32'sd2106184, 32'sd1115753, 32'sd112536, 32'sd641931, -32'sd736247, -32'sd2462920, -32'sd1123662, -32'sd384699, -32'sd1144351, 32'sd687109, 32'sd944203, 32'sd1665589, -32'sd2598078, -32'sd1378091, 32'sd1239751, 32'sd747814, 32'sd492025, -32'sd327031, 32'sd1248333, 32'sd382629, -32'sd1214333, 32'sd725822, -32'sd101027, -32'sd1540923, -32'sd2158095, 32'sd1675378, 32'sd1377270, 32'sd3033529, 32'sd2448209, 32'sd213721, -32'sd524532, 32'sd165891, -32'sd1520552, 32'sd1629026, -32'sd278868, -32'sd1395303, -32'sd2818552, -32'sd1431560, -32'sd1260914, 32'sd3668, -32'sd1622052, -32'sd108361, 32'sd937886, -32'sd44334, -32'sd272830, -32'sd798990, 32'sd847013, 32'sd1069095, -32'sd33136, 32'sd1439583, 32'sd701904, 32'sd700521, 32'sd243624, -32'sd270793, 32'sd1093038, 32'sd2583319, 32'sd2516319, 32'sd596693, 32'sd138795, 32'sd235347, -32'sd710972, 32'sd1344937, 32'sd1036929, -32'sd1181331, -32'sd957663, -32'sd845277, 32'sd233298, -32'sd1112217, -32'sd1312036, -32'sd910950, 32'sd1886086, 32'sd803387, -32'sd44167, 32'sd205973, 32'sd2481854, 32'sd2211890, -32'sd1273570, 32'sd89612, 32'sd876320, 32'sd1763902, -32'sd965979, 32'sd739760, 32'sd742195, 32'sd194530, 32'sd860975, 32'sd605062, -32'sd175669, 32'sd2138150, 32'sd1350421, 32'sd2816801, 32'sd1261927, -32'sd901111, -32'sd1230909, -32'sd1224462, 32'sd29454, -32'sd685723, -32'sd841020, -32'sd495194, 32'sd1264771, 32'sd1101479, -32'sd128486, -32'sd1635505, -32'sd459013, 32'sd1223934, -32'sd2268423, -32'sd561996, -32'sd422135, -32'sd260755, -32'sd572021, -32'sd1991396, -32'sd1820085, 32'sd953890, -32'sd127669, 32'sd1212446, -32'sd397420, -32'sd201409, -32'sd855980, 32'sd1431499, 32'sd1723575, 32'sd787231, -32'sd501395, -32'sd499818, 32'sd1593907, 32'sd645632, -32'sd698647, -32'sd1130088, 32'sd1074568, 32'sd1180398, 32'sd420408, 32'sd684480, -32'sd430776, 32'sd1429966, -32'sd2508976, -32'sd3046790, -32'sd3369051, -32'sd4686422, -32'sd5940600, -32'sd4054996, -32'sd1048600, 32'sd774716, -32'sd2005615, -32'sd662490, -32'sd1164822, -32'sd293065, -32'sd539305, 32'sd1867387, 32'sd8856, 32'sd1620474, 32'sd2296504, 32'sd2513060, 32'sd6275, 32'sd195342, 32'sd1991902, 32'sd139868, 32'sd471530, 32'sd872792, 32'sd1155918, 32'sd351048, 32'sd789151, 32'sd1251785, -32'sd893802, -32'sd1150144, -32'sd352900, -32'sd5070135, -32'sd4432874, -32'sd3181484, -32'sd2571411, -32'sd1353157, -32'sd2023493, -32'sd725357, -32'sd669410, -32'sd125661, 32'sd1125332, 32'sd1934971, 32'sd1020245, 32'sd2476612, 32'sd3131228, 32'sd2984956, -32'sd241820, -32'sd157254, -32'sd2577547, -32'sd450173, 32'sd882526, 32'sd0, 32'sd179138, -32'sd560453, -32'sd528327, 32'sd1480700, 32'sd1311964, -32'sd816352, 32'sd1203354, -32'sd65893, -32'sd1853713, -32'sd2432051, -32'sd997513, -32'sd1900496, -32'sd1207621, -32'sd340537, -32'sd1131252, -32'sd1357807, 32'sd1374042, 32'sd1081277, 32'sd136084, 32'sd2618370, 32'sd2462821, -32'sd110392, -32'sd1676477, -32'sd606076, -32'sd2521142, 32'sd547176, -32'sd349938, 32'sd451641, -32'sd6936, -32'sd154689, 32'sd504617, 32'sd2147436, 32'sd1624348, 32'sd2335411, 32'sd2010251, 32'sd2052524, 32'sd932434, -32'sd323376, 32'sd1325430, -32'sd1945099, -32'sd2178234, -32'sd2317720, -32'sd906253, 32'sd396243, 32'sd920061, -32'sd791175, -32'sd183836, 32'sd1217410, 32'sd740911, -32'sd548529, -32'sd1295108, -32'sd839291, -32'sd210543, -32'sd1582748, 32'sd199535, 32'sd485821, -32'sd247660, -32'sd321347, 32'sd952354, -32'sd44702, 32'sd1132936, 32'sd589119, 32'sd167615, 32'sd1355471, 32'sd2715415, 32'sd1155091, 32'sd2367730, 32'sd1308504, 32'sd1963563, 32'sd1883457, 32'sd2211779, 32'sd2062940, 32'sd419425, 32'sd1472768, 32'sd1179973, -32'sd183071, 32'sd364956, -32'sd27192, -32'sd508515, 32'sd199764, -32'sd1070314, -32'sd1522322, 32'sd1003855, 32'sd0, -32'sd1161709, -32'sd2102190, 32'sd1498481, 32'sd500731, -32'sd767558, -32'sd303291, 32'sd556774, 32'sd2892399, 32'sd3546751, 32'sd3197813, 32'sd2582762, 32'sd4145695, 32'sd3625662, 32'sd45164, 32'sd732058, 32'sd61551, 32'sd2154035, 32'sd416633, -32'sd317377, 32'sd708228, 32'sd934007, 32'sd38957, -32'sd125700, 32'sd714091, -32'sd61517, 32'sd19988, 32'sd1020014, 32'sd1451332, 32'sd436015, 32'sd343735, -32'sd346246, 32'sd1224000, -32'sd96075, -32'sd1145198, 32'sd113077, 32'sd1817579, 32'sd1613064, 32'sd526161, 32'sd2039910, 32'sd2387769, 32'sd2082471, 32'sd2336543, 32'sd133236, -32'sd1952545, 32'sd770047, -32'sd1253842, -32'sd1624014, 32'sd558000, -32'sd1343999, 32'sd665173, 32'sd611497, -32'sd1880474, 32'sd777520, 32'sd453918, 32'sd1765562, 32'sd720448, 32'sd982980, -32'sd1318159, -32'sd101717, 32'sd229830, -32'sd613060, 32'sd1078750, -32'sd72687, -32'sd867002, -32'sd869169, -32'sd333345, 32'sd852962, 32'sd1695097, 32'sd2048025, 32'sd990340, 32'sd1903770, 32'sd608396, 32'sd581769, -32'sd770953, -32'sd1095745, -32'sd217634, -32'sd1533715, -32'sd293936, 32'sd381121, 32'sd59210, 32'sd2070130, 32'sd1448063, 32'sd876427, 32'sd0, 32'sd1660634, 32'sd1145238, -32'sd1546938, -32'sd1856218, -32'sd874567, 32'sd1268394, 32'sd432538, 32'sd1255448, 32'sd1347578, 32'sd1366046, 32'sd2201446, 32'sd532686, -32'sd321699, 32'sd563053, 32'sd2095516, 32'sd2065159, 32'sd1847711, 32'sd519323, -32'sd952346, -32'sd555054, -32'sd1374004, -32'sd874166, 32'sd212241, 32'sd944352, -32'sd828457, 32'sd2040508, 32'sd0, 32'sd0, 32'sd0, 32'sd547678, -32'sd365580, -32'sd1578575, 32'sd109930, 32'sd56223, 32'sd2676381, 32'sd1363561, 32'sd1028879, 32'sd1350941, 32'sd1092314, 32'sd2001892, 32'sd1398187, 32'sd2095549, 32'sd518965, -32'sd454285, 32'sd1755953, 32'sd656560, -32'sd314704, 32'sd218565, 32'sd253904, 32'sd414169, 32'sd204101, 32'sd2239946, 32'sd953075, 32'sd797549, 32'sd0, 32'sd0, 32'sd0, 32'sd1635016, 32'sd547954, -32'sd850728, 32'sd183830, -32'sd476821, 32'sd1106497, 32'sd2031895, 32'sd2134218, -32'sd626096, -32'sd1888461, 32'sd1816068, 32'sd1242919, 32'sd1265932, 32'sd153272, 32'sd370378, -32'sd3870470, -32'sd2636900, -32'sd360818, -32'sd212065, -32'sd286812, -32'sd389675, 32'sd850397, 32'sd1195847, 32'sd1561510, -32'sd911831, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1170467, 32'sd913023, 32'sd538253, 32'sd1071145, -32'sd813384, 32'sd152011, 32'sd72677, 32'sd1467310, -32'sd366917, -32'sd346437, -32'sd1407957, 32'sd152918, 32'sd1160824, 32'sd609197, 32'sd1053888, -32'sd1309536, -32'sd389178, 32'sd245745, -32'sd738907, -32'sd114468, -32'sd548799, 32'sd273775, 32'sd588214, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd289986, 32'sd1462249, 32'sd322847, 32'sd1111121, 32'sd945792, 32'sd356485, 32'sd1127684, 32'sd118717, 32'sd313192, 32'sd1027521, 32'sd835255, -32'sd212966, -32'sd383587, 32'sd694946, 32'sd1462, -32'sd91826, 32'sd704095, 32'sd183614, 32'sd1521224, 32'sd501610, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1391809, 32'sd1282197, 32'sd2780896, 32'sd1834815, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2684, 32'sd766681, -32'sd100143, -32'sd1372479, 32'sd361377, -32'sd446658, 32'sd2168623, 32'sd941409, 32'sd1484388, 32'sd1175073, -32'sd354649, 32'sd2127723, 32'sd1400650, 32'sd1501726, 32'sd2199548, 32'sd982298, 32'sd192375, 32'sd1067935, 32'sd1116492, 32'sd1263945, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2216979, 32'sd1399658, 32'sd1422318, -32'sd1185704, 32'sd760982, -32'sd149605, -32'sd590739, 32'sd2251625, -32'sd39222, 32'sd1996867, -32'sd873239, -32'sd2421959, 32'sd126865, 32'sd1900194, -32'sd718010, 32'sd579622, 32'sd311897, 32'sd39223, -32'sd150542, -32'sd283218, 32'sd1434837, 32'sd931456, 32'sd365947, 32'sd2086888, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd449904, 32'sd1357171, -32'sd481889, 32'sd87514, 32'sd291095, -32'sd534696, 32'sd1069530, 32'sd2261734, -32'sd1107476, 32'sd142898, -32'sd1764381, -32'sd517847, -32'sd786546, 32'sd590690, 32'sd491892, 32'sd1962299, 32'sd1178763, 32'sd196327, 32'sd852015, -32'sd207201, 32'sd1519774, 32'sd345844, -32'sd73151, 32'sd605466, 32'sd975719, 32'sd0, 32'sd0, 32'sd1020798, 32'sd698934, -32'sd733561, -32'sd130211, 32'sd244228, -32'sd584112, 32'sd669153, 32'sd1516358, 32'sd1613645, 32'sd1008005, 32'sd118260, -32'sd620426, -32'sd2218047, -32'sd3015775, -32'sd865599, -32'sd2412518, 32'sd898705, 32'sd561860, 32'sd271679, 32'sd294222, -32'sd1203450, -32'sd1202030, 32'sd237006, -32'sd437054, -32'sd1351436, -32'sd1166557, 32'sd1205335, 32'sd0, 32'sd1317741, 32'sd1839315, 32'sd509407, 32'sd317093, -32'sd1418033, -32'sd739209, 32'sd1997292, 32'sd1303648, 32'sd964171, 32'sd1099055, 32'sd193350, -32'sd1744698, 32'sd208572, -32'sd2061122, -32'sd508035, -32'sd2391694, -32'sd1854557, -32'sd1069922, -32'sd620696, -32'sd1329360, -32'sd3622834, -32'sd2027281, -32'sd543467, -32'sd717712, -32'sd802648, -32'sd627004, 32'sd240465, 32'sd0, 32'sd305946, 32'sd973765, -32'sd1232574, -32'sd39878, 32'sd109892, 32'sd137385, 32'sd157779, -32'sd716087, 32'sd1306664, -32'sd896706, -32'sd786755, -32'sd248346, 32'sd737170, 32'sd1286602, 32'sd356637, 32'sd516722, 32'sd1714763, 32'sd916883, 32'sd520056, -32'sd626215, -32'sd1085492, -32'sd508005, -32'sd2765411, -32'sd919152, -32'sd1517000, -32'sd527413, -32'sd86162, 32'sd1390425, 32'sd1016507, 32'sd419713, 32'sd1194032, 32'sd1018238, 32'sd1581276, 32'sd123660, -32'sd1049911, -32'sd22412, -32'sd259445, -32'sd2748363, -32'sd1414825, 32'sd696883, 32'sd2613780, -32'sd169511, -32'sd2021431, -32'sd2438561, 32'sd858000, -32'sd1254068, -32'sd467956, -32'sd1018997, -32'sd2275072, -32'sd1502999, 32'sd949037, 32'sd354576, -32'sd1000499, 32'sd974355, -32'sd830300, 32'sd758719, 32'sd746021, 32'sd936038, 32'sd318022, -32'sd1292790, 32'sd747171, -32'sd318756, 32'sd670345, -32'sd75582, -32'sd1613558, -32'sd236349, 32'sd571793, 32'sd674248, 32'sd226021, 32'sd1969444, -32'sd2476521, -32'sd1787923, -32'sd2473064, 32'sd204272, -32'sd789247, -32'sd1906425, -32'sd2811457, -32'sd2062066, 32'sd177280, 32'sd514105, 32'sd201302, 32'sd388605, 32'sd1008683, 32'sd1934913, 32'sd2451232, -32'sd626898, 32'sd845891, -32'sd50997, 32'sd3137888, 32'sd2488102, 32'sd597366, -32'sd520501, -32'sd886600, 32'sd1193902, 32'sd1898385, 32'sd2749007, 32'sd1492979, 32'sd2157825, -32'sd285167, -32'sd3368076, -32'sd2286315, 32'sd476893, -32'sd1244932, -32'sd1911449, -32'sd1842810, -32'sd981903, -32'sd47824, 32'sd637892, -32'sd713548, -32'sd437291, -32'sd54867, 32'sd589561, 32'sd1203224, 32'sd1132406, 32'sd426576, 32'sd54119, 32'sd2565885, 32'sd1615653, 32'sd684816, -32'sd469226, 32'sd481419, -32'sd1724342, 32'sd1469835, 32'sd1831240, 32'sd2328050, -32'sd6303, -32'sd663949, -32'sd318653, -32'sd2576247, -32'sd417413, 32'sd1830580, 32'sd607078, -32'sd1598290, -32'sd2578499, -32'sd431796, 32'sd2581779, 32'sd402875, -32'sd502074, 32'sd411248, 32'sd92264, -32'sd932767, 32'sd406304, 32'sd1570029, 32'sd60238, -32'sd553799, -32'sd343231, 32'sd2447972, -32'sd239135, -32'sd1861618, -32'sd1830967, -32'sd500271, 32'sd1134425, -32'sd679131, 32'sd1174776, 32'sd1235203, 32'sd1546999, 32'sd66397, 32'sd972007, 32'sd2050910, 32'sd1833798, -32'sd1924993, -32'sd1480963, -32'sd30791, -32'sd1549213, -32'sd1242871, -32'sd1250476, -32'sd861192, 32'sd858820, -32'sd1362305, -32'sd271945, -32'sd689505, -32'sd558108, -32'sd36369, -32'sd2103786, 32'sd666594, -32'sd24033, -32'sd3057971, -32'sd473984, 32'sd392469, -32'sd45820, -32'sd1136833, 32'sd282937, 32'sd2011061, 32'sd2547450, -32'sd772597, 32'sd686250, 32'sd848538, -32'sd248833, 32'sd1331567, -32'sd1676483, -32'sd751315, -32'sd936833, 32'sd1758194, 32'sd742394, 32'sd41454, 32'sd107437, -32'sd225064, 32'sd529574, -32'sd1870567, -32'sd169198, -32'sd398616, -32'sd504717, -32'sd1021370, -32'sd1503841, -32'sd747419, 32'sd90506, 32'sd1659914, 32'sd1671064, 32'sd3177411, 32'sd2581714, 32'sd650126, 32'sd1273759, -32'sd1185308, -32'sd182244, 32'sd727901, 32'sd1100853, 32'sd578631, 32'sd257405, -32'sd151552, 32'sd2878884, 32'sd1514904, -32'sd961253, -32'sd1721254, 32'sd1031404, 32'sd61781, -32'sd1584593, 32'sd688528, 32'sd59832, -32'sd242672, 32'sd190436, 32'sd1263950, 32'sd546624, 32'sd355772, 32'sd2407746, 32'sd1615204, 32'sd1518625, 32'sd684592, 32'sd1025786, 32'sd1360421, 32'sd2033922, 32'sd597985, 32'sd2546776, 32'sd2535671, 32'sd1731928, 32'sd1732749, 32'sd1766886, 32'sd722039, -32'sd533345, -32'sd70149, -32'sd918050, 32'sd2608078, -32'sd367201, 32'sd415583, 32'sd475036, 32'sd282380, -32'sd55266, -32'sd1051332, -32'sd149352, -32'sd908777, 32'sd926273, 32'sd1711898, 32'sd2235765, 32'sd2957782, 32'sd840282, 32'sd686017, -32'sd139086, 32'sd2713271, -32'sd707343, 32'sd1850153, 32'sd2796071, 32'sd1794406, 32'sd896046, 32'sd2001031, -32'sd453696, -32'sd166206, 32'sd1897503, 32'sd643465, 32'sd1429418, 32'sd42683, 32'sd999262, 32'sd428285, 32'sd305633, 32'sd39347, 32'sd599853, -32'sd943760, 32'sd512769, 32'sd972401, 32'sd2334800, 32'sd42022, 32'sd689951, 32'sd3378050, 32'sd204311, 32'sd534423, 32'sd1301071, 32'sd1028895, -32'sd831073, 32'sd650995, 32'sd2256000, -32'sd156156, 32'sd599826, 32'sd2357329, 32'sd650289, 32'sd1393417, -32'sd441753, 32'sd25051, -32'sd1613540, 32'sd362811, 32'sd0, 32'sd401037, -32'sd1748473, -32'sd1598741, 32'sd1080366, 32'sd942521, -32'sd843222, -32'sd1043844, -32'sd756269, 32'sd422527, 32'sd1833390, 32'sd1059121, -32'sd979675, 32'sd369283, 32'sd1291064, 32'sd1074152, -32'sd1025369, -32'sd1088659, -32'sd129977, 32'sd1924325, 32'sd1957883, 32'sd1002378, 32'sd291369, 32'sd1982950, 32'sd780675, 32'sd1529885, -32'sd1255351, -32'sd418062, -32'sd577253, -32'sd607498, -32'sd1191577, -32'sd470194, 32'sd559114, -32'sd1383608, -32'sd2118480, -32'sd1689229, -32'sd761205, 32'sd559408, 32'sd15240, -32'sd1968426, -32'sd1340600, 32'sd160783, -32'sd211412, -32'sd2415473, -32'sd4020855, -32'sd1625591, -32'sd895295, 32'sd53711, -32'sd1743503, -32'sd1191425, -32'sd86349, 32'sd783367, 32'sd595015, -32'sd106106, -32'sd43117, -32'sd518181, 32'sd219717, 32'sd763768, 32'sd229754, -32'sd1274272, -32'sd620998, -32'sd1124388, -32'sd957416, -32'sd1337268, -32'sd2160777, -32'sd1325582, -32'sd1703056, -32'sd166692, -32'sd2141177, -32'sd1403971, 32'sd404779, -32'sd1161330, -32'sd1692848, -32'sd582316, -32'sd2572445, -32'sd1278229, -32'sd2336675, -32'sd2346173, -32'sd1295508, -32'sd982337, 32'sd79380, -32'sd686327, -32'sd429398, 32'sd1069709, 32'sd0, 32'sd8806, -32'sd302628, -32'sd840480, -32'sd375263, -32'sd135613, -32'sd2696807, -32'sd2399225, -32'sd2815585, -32'sd2803268, -32'sd2492763, -32'sd1278796, 32'sd767897, -32'sd2443399, 32'sd223209, -32'sd2174114, -32'sd216255, -32'sd2365408, -32'sd3508746, -32'sd2778486, -32'sd1938492, -32'sd2402843, -32'sd686810, -32'sd1517631, 32'sd881689, 32'sd304651, -32'sd1392416, 32'sd712982, 32'sd477162, -32'sd674091, -32'sd1732167, -32'sd871108, 32'sd369704, -32'sd778093, -32'sd1194428, -32'sd1894844, -32'sd1774388, -32'sd2318810, -32'sd738784, -32'sd1656148, -32'sd614476, -32'sd3317532, -32'sd3598275, -32'sd2037690, -32'sd1138056, -32'sd2249645, -32'sd3683137, -32'sd3064289, -32'sd3087678, -32'sd2003420, -32'sd1043151, -32'sd1887675, -32'sd100229, -32'sd436715, -32'sd623184, -32'sd264169, -32'sd882592, 32'sd643350, -32'sd1293071, 32'sd1037843, -32'sd721272, 32'sd71565, -32'sd15633, 32'sd131778, -32'sd1067685, -32'sd1625934, -32'sd134347, -32'sd2628037, -32'sd1603608, -32'sd1231746, -32'sd1691588, -32'sd1982532, -32'sd837762, -32'sd1388609, -32'sd2027106, -32'sd1587874, -32'sd439452, -32'sd3211167, -32'sd91336, -32'sd482751, -32'sd552968, -32'sd868437, -32'sd44820, 32'sd227233, 32'sd0, 32'sd1095415, -32'sd897641, -32'sd928134, -32'sd1069486, -32'sd2707731, 32'sd1183167, -32'sd534974, -32'sd533197, 32'sd164191, -32'sd869461, -32'sd3293643, -32'sd1386076, -32'sd697559, 32'sd623664, -32'sd1417321, -32'sd1912668, 32'sd208791, -32'sd714220, -32'sd868943, -32'sd2248591, -32'sd3380666, -32'sd1095841, 32'sd1049233, 32'sd852774, -32'sd44142, -32'sd1179436, 32'sd0, 32'sd0, 32'sd0, 32'sd1382264, 32'sd880313, -32'sd1740452, -32'sd310687, -32'sd1447050, 32'sd601803, 32'sd1633434, -32'sd195824, -32'sd1305422, -32'sd1375519, -32'sd265117, -32'sd1103686, -32'sd243568, 32'sd1021717, -32'sd813224, 32'sd913408, -32'sd394002, 32'sd814743, 32'sd1072334, -32'sd955999, -32'sd1733060, 32'sd1184145, -32'sd229173, -32'sd1795087, 32'sd1514988, 32'sd0, 32'sd0, 32'sd0, 32'sd484185, -32'sd125264, -32'sd52215, -32'sd1047406, -32'sd188325, 32'sd1075000, 32'sd766213, -32'sd1196424, -32'sd1265778, -32'sd616262, 32'sd207297, 32'sd696866, 32'sd1467279, 32'sd718354, 32'sd2708855, 32'sd2407454, 32'sd407580, -32'sd730399, 32'sd1442819, 32'sd986200, -32'sd1582874, -32'sd1828205, -32'sd845698, 32'sd1353404, 32'sd1735463, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1873083, 32'sd1063538, -32'sd1149811, 32'sd872586, 32'sd1561823, 32'sd73882, 32'sd789880, 32'sd744409, 32'sd66673, -32'sd98285, 32'sd1251547, 32'sd2841959, -32'sd365783, 32'sd1095032, -32'sd880422, -32'sd325421, 32'sd174671, 32'sd366394, -32'sd265214, 32'sd552933, 32'sd928396, 32'sd477781, 32'sd1277405, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2197422, 32'sd1173046, 32'sd1451031, 32'sd686804, 32'sd305494, 32'sd907006, 32'sd1403338, 32'sd1445240, -32'sd571749, 32'sd1947698, -32'sd420416, 32'sd2028478, 32'sd84504, 32'sd1891330, 32'sd592956, 32'sd204209, -32'sd612969, 32'sd841641, -32'sd359474, 32'sd2900585, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd407367, 32'sd395095, 32'sd2059319, 32'sd240510, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd788838, -32'sd1540559, -32'sd162193, -32'sd386446, -32'sd413790, 32'sd228264, -32'sd76982, 32'sd629737, -32'sd143742, -32'sd751867, 32'sd1415114, 32'sd823286, 32'sd976758, 32'sd97387, -32'sd1276169, 32'sd973608, -32'sd219330, 32'sd2459032, 32'sd1716624, 32'sd883480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1256551, 32'sd885497, -32'sd125025, -32'sd259794, -32'sd1113848, -32'sd1786911, 32'sd396585, 32'sd1456244, 32'sd970482, 32'sd483561, 32'sd415982, 32'sd1012919, 32'sd346756, 32'sd254229, 32'sd1711322, -32'sd1281914, -32'sd1940687, 32'sd478091, -32'sd309966, -32'sd146875, 32'sd137881, 32'sd383402, 32'sd518687, 32'sd1782523, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd347317, 32'sd164011, -32'sd235548, 32'sd72753, -32'sd209656, 32'sd1500930, 32'sd1488414, -32'sd137835, 32'sd1730569, 32'sd1247502, 32'sd249580, 32'sd1106693, -32'sd1976836, -32'sd1603603, -32'sd447075, -32'sd1627955, -32'sd1523791, -32'sd1308315, -32'sd267368, 32'sd28437, 32'sd19261, 32'sd734429, 32'sd233698, 32'sd532348, 32'sd1243427, 32'sd0, 32'sd0, 32'sd918591, 32'sd1422260, 32'sd1815300, -32'sd15361, 32'sd673707, 32'sd184856, 32'sd1203560, 32'sd133398, -32'sd1290193, 32'sd1287465, 32'sd864377, 32'sd1563429, 32'sd592619, 32'sd1609357, -32'sd323089, -32'sd1002885, -32'sd2595496, -32'sd3752292, -32'sd2852569, -32'sd2630956, 32'sd105502, 32'sd254904, -32'sd373057, 32'sd349862, -32'sd1458356, -32'sd13522, 32'sd815690, 32'sd0, 32'sd1532630, -32'sd242645, -32'sd795976, -32'sd576474, 32'sd2276557, 32'sd2185150, -32'sd79632, -32'sd2288, 32'sd806848, 32'sd1257839, 32'sd1079436, 32'sd2384794, 32'sd842306, 32'sd227266, 32'sd1243760, -32'sd1126944, -32'sd2740706, -32'sd2125309, -32'sd1599847, -32'sd3176987, -32'sd1268262, -32'sd681102, -32'sd683060, -32'sd1818462, -32'sd346775, -32'sd1710151, 32'sd1336143, 32'sd0, 32'sd1448812, 32'sd322273, 32'sd853918, -32'sd2035299, 32'sd68848, 32'sd632613, 32'sd422726, 32'sd682344, -32'sd1100859, 32'sd116209, -32'sd433683, 32'sd353686, -32'sd254904, -32'sd4581, -32'sd282202, 32'sd1002380, -32'sd858638, -32'sd1316498, -32'sd2118731, -32'sd3413415, -32'sd2943448, -32'sd4028856, -32'sd2218634, -32'sd882287, 32'sd2031409, -32'sd264067, -32'sd66785, 32'sd1952024, -32'sd499025, 32'sd741039, 32'sd1345363, -32'sd1356291, -32'sd1582106, -32'sd236159, -32'sd356189, 32'sd268392, 32'sd1064214, 32'sd1189952, 32'sd175085, 32'sd775578, 32'sd804668, 32'sd1291749, -32'sd1368216, 32'sd1217724, -32'sd2369684, -32'sd2302244, -32'sd5058910, -32'sd2487069, -32'sd2867029, -32'sd1578198, -32'sd2307656, 32'sd1411756, 32'sd2067128, -32'sd653021, -32'sd843298, 32'sd50705, -32'sd147062, 32'sd793455, 32'sd575900, -32'sd741530, -32'sd1887117, -32'sd116085, -32'sd1747651, -32'sd1017092, -32'sd456575, 32'sd928488, -32'sd585812, 32'sd1751732, 32'sd717071, 32'sd1626306, 32'sd2154375, 32'sd938950, 32'sd910327, -32'sd336670, -32'sd1316635, -32'sd3123412, -32'sd1768110, -32'sd52131, -32'sd1672663, 32'sd727878, -32'sd2172506, 32'sd190248, 32'sd156618, 32'sd955897, 32'sd784550, -32'sd274206, -32'sd1372502, -32'sd692366, 32'sd2570403, -32'sd969173, 32'sd998265, -32'sd1334778, 32'sd1167537, 32'sd1929767, 32'sd246498, 32'sd1658340, 32'sd4277689, 32'sd4053129, 32'sd3803141, 32'sd4553213, 32'sd1341252, -32'sd679070, -32'sd2438928, -32'sd2992423, -32'sd2321630, 32'sd1411834, 32'sd1020715, 32'sd2375900, -32'sd2594968, -32'sd637768, -32'sd577654, -32'sd639643, -32'sd1419213, -32'sd30396, -32'sd1922974, -32'sd212152, 32'sd1976723, -32'sd71885, 32'sd253563, -32'sd1192943, -32'sd355637, 32'sd2948050, 32'sd3170464, 32'sd4399429, 32'sd3654661, 32'sd2957178, 32'sd2145631, 32'sd2316712, 32'sd1020280, -32'sd58749, -32'sd3432022, -32'sd4038943, -32'sd605969, 32'sd2346355, 32'sd2413228, 32'sd1047571, -32'sd2392538, 32'sd105239, 32'sd923032, 32'sd1266450, 32'sd1100672, 32'sd444175, 32'sd116180, -32'sd1400117, -32'sd981007, -32'sd666852, 32'sd1404990, 32'sd156533, 32'sd358507, 32'sd3705316, 32'sd1823928, 32'sd517179, 32'sd2127196, 32'sd1180946, 32'sd772321, -32'sd1247758, 32'sd3439205, 32'sd3170801, -32'sd1339585, -32'sd3532840, -32'sd3696879, -32'sd689174, 32'sd2728948, 32'sd1312633, -32'sd637410, 32'sd232951, -32'sd187452, 32'sd234788, 32'sd1348381, 32'sd100555, 32'sd886496, -32'sd334122, 32'sd444962, -32'sd55270, -32'sd2516328, -32'sd2374304, 32'sd209947, 32'sd109312, -32'sd1789219, -32'sd960577, 32'sd613541, 32'sd1023676, 32'sd563053, 32'sd950730, 32'sd3510293, 32'sd528296, -32'sd3002096, -32'sd4669824, -32'sd3830848, -32'sd1337014, -32'sd199361, 32'sd202815, 32'sd364154, 32'sd558113, 32'sd1018877, 32'sd1162609, 32'sd935542, -32'sd551135, -32'sd1846085, -32'sd425076, -32'sd3017638, -32'sd610804, -32'sd1544561, -32'sd1449865, -32'sd1231874, -32'sd764689, -32'sd160612, -32'sd2244144, -32'sd1265175, 32'sd1083364, 32'sd450951, 32'sd1030927, 32'sd2347993, -32'sd1266444, -32'sd2930163, -32'sd3012779, -32'sd1967436, 32'sd234085, 32'sd657543, 32'sd2638368, 32'sd301850, 32'sd1270511, 32'sd108608, 32'sd527105, -32'sd957259, -32'sd258654, -32'sd1348099, 32'sd846324, -32'sd1457716, -32'sd2870998, -32'sd1542880, -32'sd1882853, -32'sd1170845, 32'sd334439, -32'sd1054624, -32'sd688792, -32'sd1396729, 32'sd167330, -32'sd1289896, 32'sd1729000, 32'sd794293, 32'sd104103, -32'sd2355535, -32'sd2805937, -32'sd98677, -32'sd1174718, 32'sd1710714, 32'sd267410, -32'sd1101515, 32'sd14490, 32'sd290268, 32'sd303802, -32'sd1284593, -32'sd409440, -32'sd627753, 32'sd1538795, -32'sd392058, -32'sd1483317, -32'sd2466229, -32'sd1335145, -32'sd468039, -32'sd1950343, -32'sd920997, -32'sd321860, 32'sd630801, -32'sd797751, 32'sd407610, -32'sd272469, 32'sd998808, -32'sd2208410, -32'sd1769948, -32'sd1190480, -32'sd1773246, -32'sd1213087, 32'sd151038, 32'sd953618, -32'sd1977780, -32'sd896760, 32'sd1561306, 32'sd1447422, 32'sd2236813, -32'sd91017, -32'sd9300, 32'sd222391, -32'sd684815, 32'sd639623, -32'sd404517, -32'sd1075557, 32'sd1171659, 32'sd125897, -32'sd20063, 32'sd1755068, 32'sd862860, 32'sd137791, -32'sd623358, 32'sd848946, -32'sd621149, -32'sd1173989, -32'sd921002, -32'sd1355548, 32'sd185581, 32'sd145279, 32'sd101797, 32'sd1914208, -32'sd534056, -32'sd249335, 32'sd1552395, 32'sd0, 32'sd303509, 32'sd868174, 32'sd1135022, 32'sd467957, 32'sd942237, 32'sd749939, -32'sd1664245, -32'sd510577, 32'sd1849504, -32'sd681548, 32'sd712931, -32'sd600875, -32'sd546472, 32'sd129271, -32'sd267685, 32'sd63854, -32'sd1053302, -32'sd10063, 32'sd474060, -32'sd27703, -32'sd775766, -32'sd1088697, 32'sd1512089, 32'sd149805, 32'sd2021747, 32'sd1369724, 32'sd119285, -32'sd385868, 32'sd320678, 32'sd2528, -32'sd787210, 32'sd55556, 32'sd698140, 32'sd981524, 32'sd119278, -32'sd1180957, -32'sd889323, -32'sd392616, 32'sd827616, -32'sd1073444, 32'sd1066455, -32'sd23959, -32'sd15623, -32'sd13426, -32'sd179620, -32'sd21133, 32'sd878116, -32'sd45072, -32'sd12468, 32'sd2392492, 32'sd2775745, 32'sd936711, 32'sd717347, 32'sd1583425, -32'sd584556, 32'sd376040, 32'sd899348, -32'sd1065260, -32'sd1618546, 32'sd279166, 32'sd724612, 32'sd912515, 32'sd2436122, -32'sd247154, -32'sd2065510, 32'sd578461, -32'sd1588231, -32'sd232846, 32'sd1388989, 32'sd1003007, 32'sd29445, 32'sd1400638, -32'sd359660, 32'sd258274, 32'sd673711, 32'sd1235275, 32'sd539000, 32'sd2224638, 32'sd2206034, -32'sd75998, -32'sd26108, 32'sd869591, -32'sd1317279, 32'sd0, 32'sd410029, 32'sd127238, -32'sd1645569, -32'sd533261, 32'sd1699279, -32'sd400339, -32'sd138928, -32'sd1556795, -32'sd1785422, -32'sd138464, 32'sd201111, 32'sd1882383, 32'sd1677572, -32'sd157992, 32'sd74682, 32'sd1960173, 32'sd160309, 32'sd827151, -32'sd1119405, 32'sd846767, 32'sd1118913, 32'sd2450731, -32'sd37874, 32'sd155298, -32'sd818300, 32'sd94924, 32'sd1095581, 32'sd1640083, 32'sd664990, -32'sd662374, -32'sd487930, 32'sd705440, -32'sd438604, 32'sd2240484, -32'sd1065898, -32'sd621224, -32'sd42800, 32'sd906313, -32'sd924683, 32'sd321108, 32'sd512220, 32'sd595015, 32'sd466147, -32'sd470537, -32'sd1237535, 32'sd1115553, -32'sd1019519, -32'sd398677, 32'sd1791686, 32'sd491578, 32'sd1067480, -32'sd1333388, -32'sd1279409, -32'sd475684, 32'sd1274667, 32'sd717046, 32'sd39510, 32'sd749057, 32'sd1663018, 32'sd1982468, -32'sd502616, -32'sd716320, 32'sd323566, 32'sd1268536, -32'sd425954, 32'sd115040, -32'sd1382562, 32'sd655692, 32'sd165006, 32'sd1203341, -32'sd295461, -32'sd386703, -32'sd1306712, -32'sd715899, -32'sd1760700, 32'sd1234672, 32'sd1605953, 32'sd2213956, 32'sd1770349, 32'sd1146715, -32'sd803481, -32'sd1465887, 32'sd1763025, 32'sd0, 32'sd1310323, 32'sd972101, 32'sd332188, -32'sd450587, 32'sd292359, -32'sd249706, -32'sd878650, -32'sd344938, -32'sd567988, -32'sd912274, -32'sd1244932, 32'sd1098861, 32'sd1161647, -32'sd85074, 32'sd2612710, -32'sd844476, 32'sd827188, 32'sd367075, -32'sd751356, 32'sd1809533, 32'sd1521330, 32'sd44778, 32'sd985672, 32'sd923596, 32'sd1022467, -32'sd1128396, 32'sd0, 32'sd0, 32'sd0, 32'sd1211807, 32'sd1538803, 32'sd252804, 32'sd302422, -32'sd696853, -32'sd1747377, -32'sd748808, -32'sd2402787, -32'sd2754762, -32'sd1188803, 32'sd1073458, -32'sd460357, -32'sd784778, 32'sd984837, 32'sd250874, -32'sd41929, 32'sd1733629, 32'sd589922, 32'sd49291, 32'sd987434, -32'sd591050, 32'sd2605193, -32'sd143607, 32'sd533863, 32'sd706134, 32'sd0, 32'sd0, 32'sd0, 32'sd890095, -32'sd162287, -32'sd1430351, 32'sd999196, 32'sd848909, 32'sd2514529, 32'sd1460270, -32'sd2779938, -32'sd2456561, -32'sd2538141, -32'sd991529, 32'sd140727, -32'sd819254, 32'sd1010731, 32'sd1233989, 32'sd1089308, 32'sd139631, -32'sd1091246, 32'sd132761, -32'sd1177333, -32'sd518494, -32'sd658902, -32'sd1387851, 32'sd369472, -32'sd92385, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1177478, -32'sd1207510, 32'sd1453851, 32'sd849378, 32'sd705353, 32'sd519972, -32'sd971117, 32'sd1580360, -32'sd1246676, 32'sd2535990, 32'sd1931458, -32'sd166535, -32'sd406303, -32'sd1404842, -32'sd340182, -32'sd1851882, 32'sd1104890, -32'sd225599, 32'sd1031343, 32'sd293225, 32'sd285801, 32'sd1394008, 32'sd1269077, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2292131, -32'sd255356, 32'sd1640245, 32'sd661501, 32'sd1107773, 32'sd268236, 32'sd208727, -32'sd631841, 32'sd1747133, 32'sd946246, -32'sd263407, 32'sd12221, 32'sd589250, 32'sd1310917, 32'sd754477, 32'sd532371, 32'sd451330, 32'sd1349598, 32'sd1044212, 32'sd2850019, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd574165, 32'sd1734727, -32'sd316803, 32'sd762242, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd45310, 32'sd709851, -32'sd549710, -32'sd779318, 32'sd395214, 32'sd1129525, -32'sd58070, 32'sd130046, -32'sd1922981, 32'sd229444, 32'sd891605, 32'sd541053, -32'sd366570, 32'sd1975395, 32'sd2042749, 32'sd75625, -32'sd292241, 32'sd203435, 32'sd1114958, -32'sd34427, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd578718, 32'sd1320648, -32'sd573313, 32'sd59227, -32'sd69582, 32'sd603094, -32'sd1079258, -32'sd1361731, 32'sd753627, -32'sd1378500, -32'sd176670, 32'sd1186576, -32'sd1840044, 32'sd219306, 32'sd1126927, 32'sd1880429, 32'sd1273140, -32'sd115497, 32'sd1114836, 32'sd444370, 32'sd210393, -32'sd465455, 32'sd178881, 32'sd724496, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd508882, -32'sd684466, 32'sd1133739, 32'sd520273, -32'sd77885, -32'sd1150056, -32'sd1740329, -32'sd1020766, -32'sd2026615, -32'sd1720767, -32'sd2597995, -32'sd1816119, -32'sd1753499, 32'sd2096297, 32'sd1165116, 32'sd972934, 32'sd732869, -32'sd1370973, 32'sd634769, -32'sd345477, -32'sd642083, 32'sd729792, -32'sd736237, 32'sd873417, -32'sd1174142, 32'sd0, 32'sd0, 32'sd123908, -32'sd636085, -32'sd426572, -32'sd75064, -32'sd1593282, -32'sd1373226, -32'sd368234, -32'sd644792, 32'sd1334509, -32'sd1273372, 32'sd232076, -32'sd144998, -32'sd1004741, -32'sd1282337, -32'sd685883, 32'sd1998324, -32'sd684548, -32'sd1430076, -32'sd403076, 32'sd1553071, 32'sd1809179, 32'sd480235, -32'sd366804, 32'sd508664, -32'sd309393, -32'sd388136, 32'sd301106, 32'sd0, -32'sd124546, 32'sd615455, 32'sd252110, 32'sd262422, 32'sd653529, 32'sd138837, 32'sd528308, 32'sd482506, -32'sd919679, 32'sd10787, 32'sd154784, -32'sd2133995, -32'sd448651, 32'sd141428, 32'sd924666, 32'sd568140, 32'sd943477, 32'sd1791094, 32'sd2964831, -32'sd250910, -32'sd1073895, 32'sd935957, -32'sd2449020, 32'sd381139, 32'sd1327524, 32'sd1328198, 32'sd529295, 32'sd0, 32'sd103116, -32'sd585134, 32'sd1280808, -32'sd804572, 32'sd207049, -32'sd586754, 32'sd217351, 32'sd285991, 32'sd967943, -32'sd1003318, -32'sd1434510, -32'sd1442726, -32'sd2052256, -32'sd2199216, 32'sd549451, -32'sd26827, 32'sd984971, -32'sd1011978, 32'sd844, 32'sd278123, -32'sd676499, 32'sd370909, -32'sd689206, -32'sd726883, -32'sd2579248, -32'sd102233, -32'sd1454760, 32'sd754805, 32'sd537540, 32'sd1275685, -32'sd949639, -32'sd212276, 32'sd505210, -32'sd107724, 32'sd1374716, -32'sd688889, 32'sd1235574, -32'sd1192890, 32'sd32517, 32'sd1597037, -32'sd176190, 32'sd183661, 32'sd1018488, 32'sd3049529, 32'sd1777308, -32'sd325850, -32'sd1025604, -32'sd2336049, 32'sd971264, -32'sd594687, 32'sd1781319, 32'sd1118322, -32'sd168445, -32'sd353591, 32'sd1486769, 32'sd69768, 32'sd471908, 32'sd963231, -32'sd1556366, 32'sd299808, -32'sd1578598, 32'sd710452, -32'sd186113, -32'sd1219186, -32'sd1692028, 32'sd1104920, 32'sd691391, -32'sd1483388, -32'sd1158433, -32'sd1467164, 32'sd1153010, 32'sd404738, 32'sd1482346, -32'sd416605, -32'sd875941, -32'sd849962, -32'sd550297, 32'sd496606, 32'sd991596, -32'sd835148, 32'sd660931, 32'sd2034958, -32'sd866706, 32'sd413256, -32'sd250769, 32'sd1940289, 32'sd818687, -32'sd257321, 32'sd536012, -32'sd514473, 32'sd253578, -32'sd1130521, 32'sd841281, -32'sd958382, -32'sd531224, -32'sd1835163, -32'sd1089936, -32'sd966726, -32'sd2920943, -32'sd1417822, 32'sd745981, -32'sd599164, 32'sd1700818, 32'sd3145697, -32'sd735891, -32'sd389512, 32'sd173105, -32'sd49232, 32'sd2473378, -32'sd640373, 32'sd820756, 32'sd922892, 32'sd1465312, 32'sd1155883, -32'sd591586, -32'sd697679, 32'sd197509, -32'sd30214, -32'sd601358, -32'sd1351396, 32'sd392166, 32'sd656233, 32'sd505693, -32'sd885663, -32'sd1491821, -32'sd2615933, -32'sd2422750, -32'sd1638451, 32'sd303119, 32'sd1065038, 32'sd1586461, 32'sd1438834, 32'sd568765, -32'sd1139486, -32'sd394045, 32'sd1226825, 32'sd2296382, -32'sd160901, -32'sd1223165, 32'sd773568, 32'sd136314, 32'sd79422, 32'sd1900705, -32'sd698338, -32'sd593476, 32'sd1103900, 32'sd1153722, -32'sd755044, -32'sd1575072, 32'sd852520, -32'sd1763748, 32'sd143999, 32'sd1059983, -32'sd943403, -32'sd4618423, -32'sd3043079, -32'sd1704918, 32'sd3580300, 32'sd1917714, 32'sd1347144, 32'sd154056, 32'sd347503, -32'sd6666, 32'sd868140, 32'sd532603, -32'sd712315, -32'sd162064, 32'sd233554, 32'sd1646964, 32'sd344442, -32'sd106599, -32'sd1392027, -32'sd1673321, -32'sd1056358, -32'sd489640, -32'sd865773, -32'sd1379736, 32'sd451230, -32'sd603225, -32'sd117740, 32'sd430103, -32'sd1189754, -32'sd5332588, -32'sd2180420, -32'sd3418149, 32'sd1300515, 32'sd1351047, 32'sd1836713, -32'sd102237, -32'sd1000407, -32'sd1823040, -32'sd908831, -32'sd446887, -32'sd1401665, 32'sd583728, 32'sd680706, 32'sd364765, 32'sd738175, -32'sd807916, -32'sd1112013, 32'sd346621, 32'sd2596765, 32'sd2573756, -32'sd700795, 32'sd1288406, -32'sd419453, 32'sd1453441, 32'sd2736615, -32'sd1503564, -32'sd2747982, -32'sd3730894, -32'sd3039670, -32'sd516858, -32'sd256539, -32'sd828736, -32'sd753362, -32'sd285720, -32'sd1057019, -32'sd325338, -32'sd1014976, -32'sd473727, 32'sd356058, 32'sd1426667, -32'sd640090, -32'sd571953, 32'sd1126490, -32'sd1278767, -32'sd759103, 32'sd586814, 32'sd2406820, 32'sd3369188, 32'sd1037126, 32'sd1072131, 32'sd318372, -32'sd30617, 32'sd750259, -32'sd3002685, -32'sd2696574, -32'sd3093161, -32'sd4494911, -32'sd770975, 32'sd285932, -32'sd1759031, -32'sd677901, 32'sd907930, 32'sd548443, -32'sd144113, -32'sd850046, 32'sd637726, 32'sd1898025, 32'sd1945288, 32'sd773037, 32'sd501700, 32'sd1152027, -32'sd1234765, 32'sd164773, 32'sd971748, 32'sd2501385, 32'sd1063951, 32'sd511786, 32'sd2529268, 32'sd3107739, 32'sd1255282, 32'sd397028, -32'sd4372168, -32'sd2264952, -32'sd1840491, -32'sd929316, 32'sd1653461, 32'sd622915, 32'sd55219, -32'sd546921, 32'sd284617, -32'sd691003, -32'sd978985, 32'sd1782586, -32'sd365794, -32'sd87755, 32'sd757285, 32'sd152479, 32'sd64994, -32'sd741409, -32'sd1442213, 32'sd456502, 32'sd536869, 32'sd438124, -32'sd385470, 32'sd2509749, 32'sd3168001, 32'sd2423427, 32'sd182871, -32'sd899440, -32'sd3787076, -32'sd1775317, 32'sd4352, 32'sd2464213, 32'sd1857320, 32'sd3116716, 32'sd1813324, 32'sd698376, 32'sd2851250, 32'sd1727841, -32'sd638384, 32'sd86312, -32'sd1266117, 32'sd858655, 32'sd419968, 32'sd0, 32'sd121472, 32'sd842402, -32'sd712521, -32'sd373502, -32'sd291490, 32'sd1506079, 32'sd1114011, 32'sd2169022, 32'sd1371691, 32'sd832156, 32'sd53106, -32'sd2403793, -32'sd339708, 32'sd1715775, 32'sd1680224, 32'sd3558070, 32'sd2005377, 32'sd733885, 32'sd710080, -32'sd554795, 32'sd2274534, -32'sd349003, 32'sd858975, 32'sd1038755, -32'sd514377, -32'sd496309, 32'sd1820449, 32'sd632717, 32'sd79370, -32'sd1487825, 32'sd135585, 32'sd1277814, -32'sd79932, 32'sd368074, 32'sd2903234, 32'sd3493662, 32'sd4414131, 32'sd554124, -32'sd755139, -32'sd1044352, -32'sd356746, 32'sd1251304, 32'sd2287723, 32'sd464562, 32'sd9421, 32'sd2697918, 32'sd1463008, 32'sd2799987, 32'sd1262674, 32'sd1278779, 32'sd1796910, 32'sd763192, -32'sd271744, 32'sd618573, 32'sd1177003, -32'sd250442, 32'sd891228, 32'sd477134, -32'sd348245, 32'sd33031, 32'sd371224, 32'sd753153, 32'sd1177364, 32'sd2134802, 32'sd896433, 32'sd465309, -32'sd2331372, -32'sd2705925, 32'sd82312, 32'sd2949920, 32'sd2507553, 32'sd465373, -32'sd327189, -32'sd138651, 32'sd189557, -32'sd470525, 32'sd1807535, -32'sd256398, -32'sd239956, -32'sd1229896, -32'sd516880, 32'sd11969, 32'sd1399002, 32'sd0, 32'sd1227722, 32'sd1316851, 32'sd467210, 32'sd520944, -32'sd1203929, -32'sd810640, 32'sd1877485, 32'sd53991, -32'sd586712, 32'sd754467, 32'sd64551, -32'sd1636957, -32'sd195165, 32'sd718747, -32'sd398630, -32'sd327595, 32'sd577267, -32'sd321174, -32'sd676488, -32'sd665370, 32'sd325493, 32'sd560947, -32'sd403392, -32'sd129745, -32'sd510690, 32'sd458077, 32'sd765866, -32'sd663728, -32'sd1872819, -32'sd653286, 32'sd536542, 32'sd1691647, 32'sd1280060, 32'sd426339, 32'sd1362106, -32'sd410268, 32'sd485202, -32'sd473055, -32'sd524740, 32'sd420700, -32'sd1508948, -32'sd30495, -32'sd107995, -32'sd3197545, -32'sd1125499, -32'sd997667, 32'sd1868385, 32'sd1131517, -32'sd39213, 32'sd2024973, 32'sd63322, -32'sd650885, -32'sd1350912, -32'sd1339866, 32'sd495043, 32'sd617117, -32'sd778274, 32'sd147829, 32'sd656597, 32'sd399136, 32'sd1240123, 32'sd2575763, 32'sd388704, 32'sd1137265, 32'sd1003301, -32'sd1307437, -32'sd203669, 32'sd1091739, -32'sd1773374, -32'sd743757, -32'sd3216744, -32'sd2987293, -32'sd1978993, 32'sd139335, 32'sd1633698, -32'sd220635, -32'sd634979, 32'sd203935, -32'sd973362, 32'sd827099, -32'sd1473403, -32'sd1095987, 32'sd178772, 32'sd0, 32'sd692231, 32'sd565322, 32'sd816715, -32'sd146277, -32'sd943955, -32'sd1038290, 32'sd957876, -32'sd773182, -32'sd974757, 32'sd32505, 32'sd2301723, 32'sd558366, -32'sd326672, -32'sd984615, -32'sd2373159, -32'sd3115792, -32'sd2801126, 32'sd489269, -32'sd29061, 32'sd702432, -32'sd954231, -32'sd1115981, 32'sd295610, -32'sd395766, 32'sd235787, -32'sd101334, 32'sd0, 32'sd0, 32'sd0, -32'sd1558304, -32'sd17455, 32'sd619278, -32'sd196042, -32'sd338522, 32'sd238984, -32'sd1570053, 32'sd1217787, 32'sd134, 32'sd568189, 32'sd161414, 32'sd177242, -32'sd1570150, -32'sd2203317, -32'sd2682624, -32'sd3257378, -32'sd3072415, -32'sd826962, 32'sd80051, 32'sd34243, -32'sd264364, 32'sd36604, 32'sd84621, 32'sd1631777, -32'sd743475, 32'sd0, 32'sd0, 32'sd0, 32'sd118999, 32'sd571956, -32'sd349705, 32'sd2280596, 32'sd1217024, -32'sd1539888, -32'sd1705313, -32'sd1685713, -32'sd1386956, -32'sd1576097, 32'sd36388, -32'sd763957, -32'sd1760380, 32'sd444283, -32'sd1396835, -32'sd1427056, -32'sd2435494, -32'sd939581, -32'sd152649, -32'sd1078918, -32'sd79936, -32'sd1006452, -32'sd931214, 32'sd518912, 32'sd468502, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1185134, -32'sd169652, 32'sd1439436, 32'sd2643912, -32'sd1692831, -32'sd1244403, -32'sd2096846, 32'sd341997, -32'sd1542461, 32'sd975324, -32'sd2357368, -32'sd1460458, -32'sd707151, 32'sd1256068, -32'sd964966, -32'sd1852468, 32'sd597265, -32'sd667284, 32'sd230984, 32'sd66650, 32'sd421801, 32'sd510056, 32'sd1367082, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd465663, -32'sd231572, 32'sd707550, 32'sd1424582, 32'sd194603, 32'sd1404999, 32'sd146644, -32'sd321620, -32'sd887502, 32'sd1058334, 32'sd691607, 32'sd1292537, -32'sd1113911, 32'sd1374133, -32'sd643256, 32'sd536847, 32'sd423694, 32'sd1581122, 32'sd108718, -32'sd94254, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1587991, 32'sd431386, 32'sd2116190, 32'sd2230698, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd511943, 32'sd78959, -32'sd271032, 32'sd1363633, 32'sd1716801, 32'sd179428, -32'sd11847, 32'sd662204, -32'sd21897, -32'sd1029719, -32'sd514577, 32'sd1326922, 32'sd881185, 32'sd656316, -32'sd338607, 32'sd135538, 32'sd544491, -32'sd401012, 32'sd279470, 32'sd1011704, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1825814, 32'sd626811, 32'sd68123, 32'sd791450, 32'sd1457961, -32'sd920421, -32'sd542644, 32'sd1466954, 32'sd309676, -32'sd617810, -32'sd443549, -32'sd1030015, -32'sd21625, -32'sd725407, 32'sd902336, 32'sd539907, 32'sd56893, 32'sd1529980, 32'sd459055, -32'sd668464, -32'sd838921, 32'sd421552, -32'sd78739, 32'sd1104227, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd144733, -32'sd552700, -32'sd1304076, -32'sd137090, -32'sd171521, -32'sd412926, -32'sd761398, -32'sd1544638, 32'sd2317920, -32'sd1097923, -32'sd1289128, -32'sd1161742, -32'sd739313, 32'sd448538, 32'sd1261097, 32'sd1764735, -32'sd596436, 32'sd448558, 32'sd1156737, -32'sd1377099, -32'sd1150426, -32'sd282976, -32'sd1635138, -32'sd1690236, 32'sd291122, 32'sd0, 32'sd0, 32'sd657054, -32'sd168417, 32'sd864305, -32'sd621564, -32'sd1997045, -32'sd903729, -32'sd2284385, -32'sd2801928, -32'sd1886299, 32'sd292899, 32'sd1168270, -32'sd1637094, -32'sd1118069, -32'sd141286, -32'sd260006, 32'sd1665606, 32'sd2948288, 32'sd537903, 32'sd2581877, 32'sd1170632, -32'sd395862, -32'sd23389, -32'sd1642108, -32'sd426787, 32'sd1309194, -32'sd1637487, 32'sd333309, 32'sd0, 32'sd1063296, 32'sd440974, 32'sd704772, -32'sd711508, 32'sd505045, -32'sd296092, -32'sd978159, -32'sd637006, -32'sd1771842, 32'sd1821845, -32'sd467136, 32'sd607351, -32'sd1418950, -32'sd2728308, -32'sd625708, 32'sd957797, 32'sd1249354, 32'sd312059, 32'sd1066286, -32'sd1071055, -32'sd86846, 32'sd1508411, 32'sd342663, -32'sd2693421, 32'sd441575, -32'sd1427361, 32'sd243203, 32'sd0, 32'sd192867, 32'sd2410595, 32'sd1961909, 32'sd1937769, -32'sd612467, -32'sd130227, -32'sd272830, 32'sd775576, 32'sd887998, 32'sd4140106, 32'sd3008959, 32'sd1822216, -32'sd723506, -32'sd903187, 32'sd844808, -32'sd111382, 32'sd396809, 32'sd1565330, 32'sd341366, -32'sd685527, 32'sd990412, 32'sd1372966, -32'sd1047091, -32'sd1219280, 32'sd764268, -32'sd72359, 32'sd648117, 32'sd940880, 32'sd394568, 32'sd170646, -32'sd1105159, 32'sd647008, 32'sd244934, 32'sd1502443, 32'sd2761280, 32'sd2409469, -32'sd70057, 32'sd1687426, 32'sd4146828, 32'sd2015249, -32'sd2032549, -32'sd1768829, 32'sd100213, 32'sd904389, -32'sd365929, 32'sd791630, 32'sd2838802, 32'sd1185136, -32'sd454911, -32'sd1338819, 32'sd1319185, 32'sd2256786, 32'sd1122208, 32'sd1058507, 32'sd65701, 32'sd686731, 32'sd75738, 32'sd990397, 32'sd193772, 32'sd502386, -32'sd1743596, -32'sd1374248, 32'sd1036084, 32'sd1064481, 32'sd787786, -32'sd549732, 32'sd1893450, 32'sd460791, -32'sd209545, -32'sd915424, -32'sd675915, -32'sd967931, 32'sd737395, 32'sd2239278, 32'sd1888185, 32'sd2151859, 32'sd906541, 32'sd1657783, 32'sd61448, -32'sd143604, 32'sd1309766, -32'sd678736, 32'sd345181, 32'sd626458, 32'sd612502, 32'sd450944, 32'sd1327381, -32'sd160767, -32'sd2107601, -32'sd2442105, -32'sd1095482, -32'sd1910432, -32'sd1783912, -32'sd1430804, -32'sd2877567, -32'sd2923890, -32'sd3292107, -32'sd2721224, -32'sd502171, 32'sd1000531, 32'sd1822089, 32'sd2478143, -32'sd5584, 32'sd2053314, -32'sd232735, 32'sd1171, 32'sd441599, -32'sd1741155, -32'sd1521720, -32'sd812130, -32'sd297613, -32'sd209658, 32'sd329330, 32'sd1355666, 32'sd1909739, 32'sd272609, 32'sd392806, -32'sd1100926, -32'sd3651138, -32'sd2315680, -32'sd3765883, -32'sd3756239, -32'sd4014309, -32'sd1713961, -32'sd3229992, -32'sd3589983, -32'sd516192, 32'sd690236, 32'sd520478, 32'sd842406, -32'sd685045, 32'sd2059731, 32'sd1917146, 32'sd1516587, 32'sd104771, -32'sd3535669, 32'sd1189602, -32'sd181158, -32'sd227376, 32'sd12339, 32'sd1593869, 32'sd1066198, 32'sd397142, -32'sd283648, -32'sd2355788, -32'sd3946435, -32'sd1807791, -32'sd3344628, -32'sd4835266, -32'sd4299275, -32'sd2946601, -32'sd2019142, 32'sd624260, -32'sd39930, 32'sd455539, -32'sd2038963, -32'sd44141, 32'sd2128207, -32'sd1209634, -32'sd399695, 32'sd666071, 32'sd1723647, -32'sd699043, -32'sd1217156, -32'sd2000613, 32'sd115615, 32'sd698178, 32'sd1365168, -32'sd551859, -32'sd21531, 32'sd88151, -32'sd533902, 32'sd146008, -32'sd2569166, -32'sd2136683, -32'sd3733783, -32'sd4018825, -32'sd1691633, -32'sd64023, 32'sd1458908, 32'sd1141184, 32'sd68368, -32'sd1487085, 32'sd1690257, 32'sd1302050, 32'sd643563, 32'sd86910, 32'sd734342, -32'sd1854327, -32'sd368882, -32'sd1228339, -32'sd241171, -32'sd1733863, 32'sd742461, -32'sd265597, 32'sd1091299, -32'sd1297882, 32'sd1263248, 32'sd1465436, 32'sd1779781, 32'sd966042, 32'sd163033, -32'sd982848, -32'sd340331, -32'sd1025523, 32'sd543246, 32'sd1314661, 32'sd352529, -32'sd22520, -32'sd352659, -32'sd1993393, -32'sd399026, -32'sd200059, 32'sd833997, -32'sd1065856, 32'sd1308960, 32'sd1062198, -32'sd267898, 32'sd779547, 32'sd450873, 32'sd777645, 32'sd876381, 32'sd999626, 32'sd1434463, 32'sd12011, -32'sd602033, -32'sd1019267, 32'sd1071583, 32'sd1397051, 32'sd480000, 32'sd650753, 32'sd1221009, 32'sd3383860, 32'sd2116727, 32'sd2474738, 32'sd1333932, 32'sd323196, -32'sd1595935, -32'sd690600, 32'sd821735, 32'sd1556186, -32'sd226089, -32'sd99560, 32'sd412241, 32'sd1175077, 32'sd2256758, 32'sd240001, 32'sd404479, -32'sd218821, 32'sd821896, -32'sd388972, -32'sd1383358, -32'sd759050, -32'sd848385, 32'sd2291316, 32'sd557458, 32'sd1330455, 32'sd1565030, 32'sd307988, -32'sd400243, 32'sd2776051, 32'sd1569970, 32'sd2190273, 32'sd2958111, 32'sd2577526, -32'sd137344, 32'sd612862, 32'sd1958326, 32'sd806650, 32'sd44836, -32'sd1345918, 32'sd670891, 32'sd1900835, 32'sd752449, 32'sd103824, 32'sd583728, -32'sd257426, 32'sd359882, 32'sd19159, 32'sd698166, 32'sd960623, 32'sd720991, 32'sd1078758, 32'sd544292, 32'sd2003971, 32'sd1684712, 32'sd148852, 32'sd1032698, 32'sd2693308, 32'sd2193028, 32'sd1868400, 32'sd2748629, 32'sd2873096, 32'sd1625383, 32'sd70100, -32'sd34080, 32'sd817480, 32'sd480295, -32'sd367324, -32'sd793475, 32'sd746094, 32'sd245178, -32'sd240835, 32'sd76281, -32'sd413677, -32'sd282329, 32'sd667032, 32'sd0, 32'sd1259529, -32'sd103316, -32'sd862521, 32'sd1559939, 32'sd1737494, -32'sd1974541, -32'sd1249218, -32'sd995103, -32'sd1392312, -32'sd1776645, -32'sd2532309, -32'sd865365, 32'sd843463, -32'sd888229, 32'sd351438, -32'sd1503281, -32'sd319351, 32'sd727017, -32'sd786230, -32'sd2409046, -32'sd2167820, -32'sd3179892, -32'sd444886, -32'sd663707, -32'sd1098988, -32'sd661955, 32'sd859318, 32'sd238266, 32'sd1082928, 32'sd563424, 32'sd950330, -32'sd501836, -32'sd1508905, -32'sd3108327, -32'sd1154742, -32'sd779419, -32'sd1135136, -32'sd3558235, -32'sd2289988, -32'sd5590418, -32'sd1953986, -32'sd1718350, -32'sd1147037, -32'sd288235, -32'sd899646, -32'sd902928, -32'sd2373263, -32'sd2200246, -32'sd1422753, -32'sd1861501, 32'sd326844, -32'sd815943, -32'sd1235715, -32'sd1071754, -32'sd155969, 32'sd1077834, 32'sd793387, 32'sd795094, -32'sd121160, -32'sd2413969, -32'sd870923, -32'sd707125, -32'sd510533, 32'sd75729, -32'sd725708, -32'sd2686579, -32'sd2052913, -32'sd3620377, -32'sd646951, 32'sd164261, 32'sd873787, 32'sd472632, -32'sd961954, -32'sd1280709, -32'sd2325448, 32'sd562605, -32'sd1254893, -32'sd588489, 32'sd1107546, -32'sd1293214, -32'sd119841, 32'sd102311, 32'sd791469, 32'sd0, -32'sd1475447, 32'sd1109335, 32'sd203971, 32'sd1138715, -32'sd1745999, -32'sd541379, -32'sd284895, 32'sd893942, -32'sd1232842, -32'sd868222, -32'sd825988, -32'sd903440, -32'sd88055, 32'sd2349276, 32'sd604881, 32'sd237951, -32'sd116246, 32'sd686301, -32'sd588191, 32'sd11869, -32'sd1537783, -32'sd922607, -32'sd1299187, 32'sd1229617, -32'sd102466, -32'sd689446, 32'sd794018, 32'sd516400, 32'sd475577, 32'sd17783, 32'sd2059326, 32'sd694838, -32'sd797530, 32'sd385733, 32'sd490744, 32'sd1078662, -32'sd957616, -32'sd1603728, -32'sd965888, -32'sd208728, 32'sd711396, 32'sd354669, 32'sd2557545, -32'sd253717, -32'sd56840, 32'sd346777, 32'sd345840, 32'sd780136, -32'sd761272, -32'sd543586, -32'sd892156, 32'sd2835517, 32'sd2533026, -32'sd97401, 32'sd1092635, 32'sd1601047, 32'sd1210753, 32'sd758828, 32'sd1283923, 32'sd1187526, 32'sd1655359, 32'sd1345090, 32'sd1567671, -32'sd1413438, -32'sd2591846, -32'sd1861662, -32'sd356651, -32'sd1674037, 32'sd1671082, 32'sd105555, 32'sd1961124, -32'sd145470, 32'sd332945, 32'sd913783, 32'sd81730, -32'sd17212, -32'sd2378984, -32'sd815506, -32'sd434039, -32'sd207400, 32'sd972499, 32'sd1708284, 32'sd1619892, 32'sd0, 32'sd1448205, 32'sd817294, -32'sd865149, 32'sd708152, 32'sd381740, 32'sd654010, 32'sd1588322, 32'sd991824, -32'sd691651, -32'sd58255, 32'sd151548, -32'sd1077886, 32'sd674291, -32'sd572466, 32'sd967323, -32'sd301677, -32'sd1751117, -32'sd1411568, 32'sd582190, -32'sd199393, -32'sd1746599, -32'sd197409, 32'sd604962, 32'sd1441991, -32'sd609916, 32'sd1492756, 32'sd0, 32'sd0, 32'sd0, 32'sd532980, -32'sd103164, 32'sd830144, -32'sd94565, -32'sd973441, -32'sd728034, 32'sd1741323, -32'sd1159836, -32'sd1556362, -32'sd991058, -32'sd1538233, 32'sd73905, 32'sd129855, -32'sd1426046, 32'sd958306, 32'sd255916, 32'sd355196, -32'sd1319385, 32'sd782502, -32'sd1040913, 32'sd972277, 32'sd1294827, 32'sd1302790, 32'sd1824849, 32'sd871555, 32'sd0, 32'sd0, 32'sd0, 32'sd362130, 32'sd1142946, 32'sd246445, -32'sd945499, -32'sd1380307, -32'sd69575, -32'sd645398, -32'sd1261775, 32'sd565802, -32'sd159548, -32'sd395023, 32'sd875803, 32'sd1001151, 32'sd527768, 32'sd1642318, -32'sd373150, 32'sd104518, -32'sd942745, -32'sd175492, -32'sd448699, -32'sd1211354, 32'sd1923276, -32'sd496748, 32'sd525166, 32'sd1618152, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1430196, 32'sd1141117, 32'sd458475, 32'sd793897, -32'sd807707, -32'sd1131588, -32'sd828574, 32'sd264676, -32'sd2804845, -32'sd1210317, 32'sd769839, -32'sd1199246, 32'sd618377, 32'sd1461791, 32'sd977072, 32'sd479772, -32'sd1724590, -32'sd931671, -32'sd835385, -32'sd711221, -32'sd407620, 32'sd1061503, 32'sd888091, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd813523, 32'sd696623, 32'sd234393, 32'sd530193, 32'sd1085375, 32'sd565117, 32'sd599690, 32'sd139958, 32'sd897739, 32'sd133554, -32'sd46453, -32'sd1479774, -32'sd699560, 32'sd429175, -32'sd441235, 32'sd740607, 32'sd68235, 32'sd382660, -32'sd539831, 32'sd1486589, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd53114, 32'sd307433, 32'sd1655754, -32'sd602669, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd407778, 32'sd3230, 32'sd1486175, -32'sd632264, -32'sd198374, 32'sd917404, 32'sd1845659, 32'sd991610, 32'sd940081, -32'sd368093, 32'sd1309108, 32'sd810049, 32'sd1765280, 32'sd191360, 32'sd577435, -32'sd466994, 32'sd504206, 32'sd853026, 32'sd970585, 32'sd1018192, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd789369, -32'sd549305, 32'sd349880, 32'sd1111475, 32'sd1571887, 32'sd1003874, -32'sd732298, 32'sd939729, 32'sd723435, -32'sd905311, -32'sd1117664, -32'sd323082, -32'sd57242, -32'sd109990, 32'sd679936, -32'sd256059, 32'sd781835, 32'sd1652367, 32'sd388409, 32'sd1967730, 32'sd1135553, 32'sd1431478, 32'sd289550, 32'sd2473613, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd160532, -32'sd401521, 32'sd1118388, -32'sd1847574, -32'sd2192699, 32'sd66764, -32'sd1478869, -32'sd438813, -32'sd1213615, 32'sd414242, -32'sd326582, -32'sd1296595, -32'sd2629780, -32'sd766458, -32'sd508399, -32'sd1498281, -32'sd458696, -32'sd481658, -32'sd462996, 32'sd2124469, 32'sd1961491, -32'sd1042733, 32'sd225379, 32'sd489288, 32'sd899639, 32'sd0, 32'sd0, 32'sd725085, 32'sd53973, 32'sd225767, -32'sd1373010, -32'sd646738, -32'sd86815, -32'sd791403, -32'sd1435756, -32'sd773199, -32'sd22705, -32'sd328653, 32'sd942799, -32'sd45598, 32'sd64480, -32'sd1145163, 32'sd18679, -32'sd528150, -32'sd533995, -32'sd1889389, 32'sd184394, 32'sd769508, -32'sd478910, 32'sd221749, -32'sd2503139, 32'sd156008, 32'sd182961, 32'sd615292, 32'sd0, 32'sd1822407, 32'sd1174387, 32'sd1373853, 32'sd272811, -32'sd159210, -32'sd1333543, -32'sd1008152, -32'sd828002, -32'sd1526959, 32'sd279990, -32'sd359426, -32'sd1045790, -32'sd1355290, -32'sd650308, -32'sd1042275, 32'sd58410, -32'sd1249160, -32'sd1166410, 32'sd592272, 32'sd891006, 32'sd2457082, 32'sd1134988, 32'sd1373422, -32'sd233516, 32'sd500174, -32'sd302480, 32'sd870589, 32'sd0, 32'sd642722, -32'sd143495, -32'sd368769, 32'sd510670, -32'sd1954442, -32'sd947975, -32'sd1261416, -32'sd833693, 32'sd937033, -32'sd477026, 32'sd530215, -32'sd1087328, 32'sd594065, 32'sd1891673, 32'sd705087, 32'sd935365, 32'sd489516, 32'sd864700, 32'sd336154, -32'sd1553909, 32'sd625829, 32'sd957584, -32'sd548566, -32'sd288439, 32'sd592093, 32'sd1160239, 32'sd116354, 32'sd1674242, 32'sd130554, 32'sd946433, 32'sd223030, 32'sd220197, -32'sd1262952, -32'sd2913168, -32'sd1647282, 32'sd208687, -32'sd268296, -32'sd1680197, 32'sd144194, -32'sd1703865, 32'sd1557224, 32'sd2710361, 32'sd910763, 32'sd2515334, -32'sd629618, -32'sd272614, 32'sd2670242, -32'sd405772, 32'sd842486, 32'sd618608, -32'sd1855360, -32'sd1301488, -32'sd518929, 32'sd301567, 32'sd728535, 32'sd814635, 32'sd241173, -32'sd1122444, 32'sd1022912, -32'sd944048, -32'sd1319408, -32'sd2858247, -32'sd1416531, -32'sd1197810, 32'sd853693, -32'sd801573, 32'sd89200, -32'sd559147, 32'sd2100923, 32'sd2678783, 32'sd2941586, 32'sd615919, -32'sd505243, -32'sd3215517, 32'sd291188, 32'sd6389, -32'sd37235, -32'sd591821, 32'sd300400, -32'sd942967, -32'sd1697410, -32'sd736269, -32'sd511443, 32'sd681090, -32'sd1210264, 32'sd72523, 32'sd1493887, 32'sd2296771, 32'sd502612, -32'sd1546699, 32'sd1001702, -32'sd621479, 32'sd1282226, 32'sd391460, 32'sd92170, -32'sd334896, 32'sd2174685, 32'sd3098380, 32'sd2966685, 32'sd336915, -32'sd216091, -32'sd537138, -32'sd1778714, -32'sd481538, -32'sd847143, -32'sd475835, -32'sd247339, -32'sd301924, 32'sd539601, 32'sd418577, -32'sd79185, -32'sd32243, 32'sd1257035, 32'sd214561, -32'sd1800228, 32'sd462304, 32'sd517933, -32'sd927162, -32'sd1155577, 32'sd187973, -32'sd588916, -32'sd87077, -32'sd166398, -32'sd46841, 32'sd1422213, 32'sd1844345, 32'sd420164, -32'sd506387, -32'sd923630, -32'sd1983184, -32'sd23804, -32'sd1289850, -32'sd747511, -32'sd498584, 32'sd849769, 32'sd684246, -32'sd15305, -32'sd870354, -32'sd460191, 32'sd675889, 32'sd1034178, 32'sd487009, -32'sd565055, -32'sd155132, -32'sd1770757, -32'sd1158448, -32'sd1218386, -32'sd567773, -32'sd943745, 32'sd685393, 32'sd138532, -32'sd2617204, -32'sd3050730, 32'sd793071, 32'sd56362, -32'sd883835, -32'sd3984335, -32'sd2535291, 32'sd317189, 32'sd100600, -32'sd911101, 32'sd1468738, 32'sd2165195, -32'sd490905, -32'sd443018, -32'sd624956, -32'sd35920, 32'sd600332, -32'sd960310, -32'sd372574, -32'sd1933095, -32'sd2278998, -32'sd1970307, -32'sd1723079, -32'sd1949544, -32'sd537564, 32'sd599179, -32'sd37184, -32'sd3663421, -32'sd4414924, -32'sd3419239, 32'sd408797, -32'sd875387, -32'sd2004674, -32'sd2765893, -32'sd1882428, -32'sd2593078, -32'sd80847, 32'sd118371, 32'sd1623083, 32'sd1178452, -32'sd400770, -32'sd1442278, 32'sd784182, -32'sd995745, 32'sd721283, 32'sd637155, 32'sd275426, -32'sd1873025, -32'sd403110, -32'sd2276157, -32'sd1938524, -32'sd1152320, -32'sd1372910, -32'sd1863312, -32'sd3407375, -32'sd3446814, -32'sd653233, -32'sd901542, 32'sd1591644, -32'sd1245114, 32'sd123909, -32'sd2357173, -32'sd2009926, -32'sd696625, -32'sd1110457, -32'sd1411071, 32'sd392034, 32'sd18448, -32'sd805327, 32'sd551811, 32'sd1530041, 32'sd1359727, 32'sd1098180, 32'sd128880, -32'sd515291, 32'sd749149, -32'sd1256609, -32'sd964889, -32'sd909969, -32'sd1471580, -32'sd1222899, -32'sd1779932, -32'sd2220269, -32'sd1182043, 32'sd62557, 32'sd648038, 32'sd3785259, 32'sd725155, -32'sd77553, -32'sd2235366, -32'sd2050261, -32'sd2444450, -32'sd3505885, -32'sd2054621, -32'sd2004912, 32'sd75455, 32'sd1410688, 32'sd811736, 32'sd699954, 32'sd1956530, -32'sd622552, 32'sd1369507, 32'sd285185, 32'sd12981, -32'sd431434, -32'sd488678, -32'sd539670, -32'sd1448090, -32'sd1299893, 32'sd363035, 32'sd2518849, 32'sd2050268, 32'sd3487173, 32'sd5070958, 32'sd804802, -32'sd177467, -32'sd1070677, -32'sd2097644, -32'sd1071885, -32'sd2634944, -32'sd2198280, -32'sd1818670, -32'sd3199480, -32'sd2753746, -32'sd1876030, -32'sd1058463, 32'sd683777, 32'sd212421, 32'sd102831, 32'sd1052691, -32'sd1186478, -32'sd1058738, 32'sd362536, -32'sd1112779, 32'sd1760067, -32'sd711391, -32'sd821425, 32'sd5114628, 32'sd5122838, 32'sd1912300, 32'sd1769307, 32'sd2017122, 32'sd2293309, -32'sd110975, -32'sd1157378, -32'sd2534592, -32'sd1552666, -32'sd3305075, -32'sd2867828, -32'sd425178, -32'sd675637, -32'sd345532, -32'sd628881, 32'sd701394, 32'sd589185, 32'sd396750, 32'sd0, -32'sd902868, -32'sd183087, -32'sd206550, 32'sd263194, -32'sd141164, 32'sd2074990, 32'sd1442722, 32'sd2499546, 32'sd898850, 32'sd1456208, 32'sd1180264, 32'sd1273169, 32'sd1928635, 32'sd2498501, -32'sd709312, -32'sd1057842, -32'sd99628, -32'sd381323, -32'sd651958, -32'sd1348832, 32'sd1505727, -32'sd714032, -32'sd612820, -32'sd1565043, 32'sd233470, 32'sd1956606, 32'sd757921, 32'sd206500, 32'sd1569440, 32'sd287556, -32'sd876664, -32'sd123039, 32'sd1671144, 32'sd959204, 32'sd2017887, 32'sd659857, 32'sd281510, 32'sd1634942, -32'sd796100, 32'sd538047, 32'sd1845212, 32'sd361079, -32'sd1540245, -32'sd1987537, 32'sd1016428, 32'sd2524929, 32'sd2273764, 32'sd1986420, 32'sd2272571, -32'sd665267, 32'sd823739, -32'sd564845, 32'sd840161, -32'sd585626, 32'sd918820, 32'sd1283972, 32'sd767728, 32'sd912659, -32'sd935670, 32'sd1879620, -32'sd207547, 32'sd2022576, 32'sd1969806, 32'sd2212006, 32'sd1229653, -32'sd38570, 32'sd1479893, 32'sd748158, 32'sd896032, -32'sd79241, 32'sd486404, 32'sd583854, 32'sd1696705, 32'sd2115141, 32'sd2366534, 32'sd1635178, 32'sd1613708, 32'sd1419039, 32'sd1750902, -32'sd1730384, 32'sd1658938, 32'sd606254, 32'sd2238425, 32'sd0, -32'sd146364, -32'sd283162, -32'sd871866, 32'sd591437, 32'sd1091685, 32'sd3146777, 32'sd2398534, 32'sd1078232, -32'sd787311, 32'sd50862, -32'sd1058072, -32'sd1149131, -32'sd1527725, -32'sd892215, 32'sd2444548, 32'sd1549505, 32'sd1172733, 32'sd3006355, 32'sd2523939, 32'sd3290089, 32'sd3030062, 32'sd1813704, 32'sd2856750, 32'sd291685, 32'sd546074, 32'sd121349, 32'sd1104104, -32'sd652078, -32'sd1068237, 32'sd1916261, 32'sd1767838, 32'sd458294, 32'sd1724278, 32'sd1080054, -32'sd869676, 32'sd135367, 32'sd237438, -32'sd917492, -32'sd1031051, 32'sd945303, -32'sd171199, 32'sd1300663, 32'sd606313, -32'sd685052, 32'sd1992045, 32'sd875200, 32'sd2338614, 32'sd1847144, 32'sd1986498, 32'sd986933, 32'sd43823, 32'sd1027626, -32'sd451809, -32'sd366025, 32'sd220566, 32'sd417229, -32'sd674622, -32'sd169498, 32'sd886082, 32'sd348555, 32'sd1858907, 32'sd1725338, 32'sd1851029, -32'sd841117, 32'sd536291, -32'sd723958, 32'sd14767, 32'sd1869460, 32'sd2155413, -32'sd1637762, -32'sd630684, -32'sd1008302, -32'sd1545213, -32'sd239656, 32'sd691433, 32'sd2320289, 32'sd114623, 32'sd951728, 32'sd2196549, 32'sd515212, -32'sd22248, 32'sd604590, -32'sd88019, 32'sd0, 32'sd1763329, 32'sd791363, -32'sd971485, 32'sd606415, -32'sd1031846, 32'sd1372030, -32'sd864766, -32'sd222486, -32'sd1543428, 32'sd192391, -32'sd509467, 32'sd1671240, -32'sd620154, -32'sd1557029, 32'sd947276, 32'sd466776, 32'sd248020, -32'sd352542, -32'sd963269, -32'sd393001, 32'sd731915, 32'sd1048967, 32'sd1638762, -32'sd187496, 32'sd681195, 32'sd1408355, 32'sd0, 32'sd0, 32'sd0, -32'sd1048070, 32'sd560134, 32'sd1824488, 32'sd677508, -32'sd1013059, -32'sd779368, 32'sd56398, -32'sd1190088, -32'sd3230211, -32'sd2806167, -32'sd2533527, -32'sd1138352, -32'sd2095140, -32'sd3543991, -32'sd1947011, -32'sd1516454, -32'sd2656955, -32'sd2736833, -32'sd2058590, -32'sd1262044, 32'sd895896, 32'sd344519, -32'sd597686, -32'sd51943, 32'sd505477, 32'sd0, 32'sd0, 32'sd0, 32'sd1025315, 32'sd1027028, 32'sd403104, -32'sd525401, -32'sd742845, -32'sd768067, -32'sd162748, -32'sd2833325, -32'sd3796040, 32'sd36468, -32'sd1056199, -32'sd116116, 32'sd151996, -32'sd610091, -32'sd415787, 32'sd562437, 32'sd654871, -32'sd933234, -32'sd2341073, -32'sd241132, 32'sd341602, -32'sd842864, -32'sd102339, 32'sd1275742, 32'sd934267, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1653514, 32'sd612303, -32'sd256431, 32'sd187578, 32'sd1018879, -32'sd914079, -32'sd451020, -32'sd135211, 32'sd696338, 32'sd373207, 32'sd152218, -32'sd497172, -32'sd518474, -32'sd1989926, -32'sd69133, -32'sd143845, 32'sd321033, -32'sd1207499, 32'sd719215, -32'sd943480, -32'sd1467814, 32'sd131373, 32'sd1049874, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1054296, 32'sd1143999, 32'sd359825, 32'sd1146416, -32'sd1339021, 32'sd406427, 32'sd1746027, 32'sd1672640, 32'sd797623, 32'sd1659990, 32'sd1215041, -32'sd310223, 32'sd1267304, 32'sd192248, -32'sd124781, 32'sd2141998, 32'sd3642858, -32'sd390365, -32'sd772832, 32'sd435073, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd554792, 32'sd277630, -32'sd744888, 32'sd1038432, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd56385, -32'sd673893, -32'sd1116341, -32'sd232835, -32'sd331413, -32'sd747005, 32'sd602611, -32'sd1274363, -32'sd191797, -32'sd248963, 32'sd133910, -32'sd201899, 32'sd1095476, 32'sd1417322, 32'sd1280808, 32'sd1026516, -32'sd232780, 32'sd1214525, -32'sd46297, -32'sd95031, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd151058, 32'sd157078, 32'sd687406, 32'sd1776242, 32'sd716650, -32'sd770457, 32'sd631003, -32'sd1121546, 32'sd95300, 32'sd494407, 32'sd256064, -32'sd1943425, -32'sd1737782, -32'sd1140925, -32'sd1604359, -32'sd86729, 32'sd168665, -32'sd654899, 32'sd267189, 32'sd688565, -32'sd205903, 32'sd266768, 32'sd417110, -32'sd358154, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd265270, -32'sd715679, 32'sd18840, 32'sd1179684, 32'sd538163, -32'sd595456, -32'sd538856, 32'sd2178851, 32'sd1543172, 32'sd222864, -32'sd910104, 32'sd605526, 32'sd129545, -32'sd110476, -32'sd1514134, 32'sd369578, 32'sd1310187, 32'sd674027, 32'sd213842, 32'sd677647, -32'sd678121, 32'sd1064486, 32'sd593105, 32'sd1162304, 32'sd459685, 32'sd0, 32'sd0, 32'sd695272, 32'sd430747, -32'sd930486, -32'sd1260974, -32'sd185676, 32'sd1151267, 32'sd141349, 32'sd425667, 32'sd2306064, 32'sd1415392, -32'sd161726, -32'sd397285, -32'sd1695821, -32'sd1764606, 32'sd306141, 32'sd717127, 32'sd48652, 32'sd1493894, -32'sd563883, -32'sd67606, -32'sd498184, -32'sd1419623, 32'sd728079, 32'sd642459, 32'sd424227, 32'sd1117750, -32'sd279903, 32'sd0, 32'sd251890, 32'sd498701, -32'sd2097944, 32'sd672980, 32'sd1043745, -32'sd510112, 32'sd1135162, 32'sd1432652, 32'sd949236, -32'sd914971, -32'sd541410, -32'sd418972, 32'sd1078697, 32'sd1342018, -32'sd1278548, -32'sd2106492, -32'sd1432142, -32'sd69669, -32'sd691017, 32'sd581937, 32'sd1582396, -32'sd1017223, 32'sd913200, -32'sd236866, -32'sd381206, 32'sd388168, -32'sd16446, 32'sd0, 32'sd373342, -32'sd922649, -32'sd1494858, 32'sd18387, 32'sd546803, -32'sd357509, -32'sd34369, 32'sd959046, -32'sd592326, 32'sd2381037, 32'sd787745, 32'sd1858997, 32'sd692111, 32'sd675036, 32'sd1948707, 32'sd411883, -32'sd1398298, 32'sd1007053, 32'sd1297138, -32'sd25715, 32'sd1972444, 32'sd786608, 32'sd55913, 32'sd720558, 32'sd72993, -32'sd61520, -32'sd655726, 32'sd399245, 32'sd1062094, 32'sd229817, -32'sd3251034, -32'sd1614396, -32'sd1287386, 32'sd478535, 32'sd281333, 32'sd960622, 32'sd1205988, 32'sd2329122, 32'sd3019440, 32'sd1148982, 32'sd4341434, 32'sd2532524, 32'sd2047400, 32'sd1972745, 32'sd615409, -32'sd845781, -32'sd847344, 32'sd1432006, -32'sd792625, -32'sd1174335, -32'sd2185992, -32'sd1425571, -32'sd711709, 32'sd107354, -32'sd183788, 32'sd700982, -32'sd281276, -32'sd1216742, -32'sd735652, -32'sd2082592, -32'sd107832, 32'sd1028389, 32'sd549202, -32'sd460817, 32'sd1539194, 32'sd3523432, 32'sd1747050, 32'sd2938131, 32'sd3226542, 32'sd2794222, 32'sd1192970, 32'sd1042438, -32'sd230947, -32'sd1027887, -32'sd633811, 32'sd175166, -32'sd2291629, -32'sd2617488, -32'sd3231065, -32'sd585875, -32'sd1459578, -32'sd1014739, -32'sd1564086, 32'sd220017, -32'sd1248795, 32'sd1834399, 32'sd281305, 32'sd642205, -32'sd33321, 32'sd962254, 32'sd706716, 32'sd148219, 32'sd3436428, 32'sd126059, -32'sd1233486, 32'sd1029998, 32'sd796287, 32'sd275260, -32'sd954602, -32'sd796117, -32'sd651506, 32'sd2061037, 32'sd576077, -32'sd552700, -32'sd10024, -32'sd752220, -32'sd1735721, 32'sd403156, -32'sd287477, -32'sd1552604, 32'sd1294713, 32'sd249177, -32'sd1746583, 32'sd1959482, -32'sd1248879, 32'sd314819, 32'sd694340, 32'sd2001542, 32'sd113523, 32'sd679305, 32'sd979693, 32'sd1527020, 32'sd279029, -32'sd2445454, 32'sd113064, -32'sd1216569, -32'sd661782, -32'sd575780, 32'sd1730404, 32'sd1875731, -32'sd398428, -32'sd1185402, 32'sd286000, 32'sd1329016, -32'sd424718, -32'sd1277531, -32'sd754346, -32'sd420583, 32'sd28867, 32'sd355059, -32'sd72964, -32'sd351025, -32'sd462610, -32'sd63789, 32'sd1296957, 32'sd1039171, -32'sd721567, 32'sd1088849, 32'sd1083383, 32'sd312663, -32'sd115606, -32'sd2989319, -32'sd2989076, -32'sd3657739, -32'sd1694527, -32'sd292495, -32'sd985169, 32'sd264576, -32'sd17907, 32'sd482162, 32'sd1509153, 32'sd1997524, 32'sd2134604, 32'sd482662, -32'sd1671850, 32'sd548766, 32'sd1224468, 32'sd237144, 32'sd1414952, -32'sd532727, -32'sd822247, 32'sd779254, -32'sd714751, 32'sd1790990, 32'sd595606, -32'sd880182, -32'sd498725, -32'sd989615, -32'sd2607430, -32'sd3032289, -32'sd1433228, -32'sd1140919, -32'sd867757, 32'sd652118, -32'sd1158210, -32'sd235634, -32'sd1247131, 32'sd1282532, 32'sd2146066, 32'sd575751, 32'sd999342, -32'sd1615169, -32'sd787542, 32'sd549475, -32'sd1075205, -32'sd4893, 32'sd378483, 32'sd992630, 32'sd1376123, 32'sd1193351, -32'sd938235, 32'sd981920, 32'sd709194, -32'sd24558, -32'sd1042132, -32'sd702536, -32'sd2463861, -32'sd425465, -32'sd1510562, -32'sd827485, -32'sd2600053, -32'sd1793570, -32'sd1819795, -32'sd1330332, -32'sd403141, 32'sd1974634, -32'sd250100, -32'sd296035, -32'sd1284725, 32'sd1936939, 32'sd2111438, 32'sd316875, 32'sd1051002, -32'sd101664, 32'sd695629, 32'sd1294500, 32'sd1019863, -32'sd1539504, -32'sd2150151, -32'sd1836996, -32'sd1068494, 32'sd445777, -32'sd1185041, -32'sd195699, -32'sd2138510, -32'sd1292200, -32'sd1289285, -32'sd1866968, -32'sd1427183, -32'sd3664418, -32'sd1571105, 32'sd119117, 32'sd182679, 32'sd1982897, -32'sd657130, -32'sd860556, -32'sd222156, 32'sd1065883, -32'sd371902, 32'sd1161176, 32'sd23676, -32'sd143748, -32'sd118511, 32'sd869006, -32'sd6632, 32'sd344992, -32'sd118393, -32'sd2381450, -32'sd1913905, -32'sd889484, -32'sd1161005, 32'sd770655, 32'sd699571, 32'sd362280, 32'sd170448, -32'sd1898090, -32'sd868804, -32'sd2632262, -32'sd1770103, 32'sd1483598, -32'sd821955, 32'sd1572023, 32'sd1802382, 32'sd910621, 32'sd368838, 32'sd1342670, -32'sd1685662, 32'sd1375726, 32'sd196373, 32'sd333412, 32'sd1350614, -32'sd513173, -32'sd1107295, 32'sd365397, 32'sd570725, 32'sd61600, 32'sd113524, -32'sd1036457, -32'sd685523, 32'sd2388715, 32'sd1681386, 32'sd2839639, 32'sd1509083, 32'sd439439, -32'sd2325196, -32'sd3409001, -32'sd1070013, -32'sd1741939, -32'sd42292, 32'sd677617, -32'sd287767, -32'sd529033, 32'sd1419634, -32'sd881958, 32'sd125314, 32'sd42923, -32'sd1557425, 32'sd0, -32'sd293659, -32'sd1014819, 32'sd120852, 32'sd23192, 32'sd1842301, 32'sd352410, -32'sd183553, -32'sd1414698, -32'sd122399, 32'sd195658, -32'sd522547, 32'sd795419, 32'sd1254051, -32'sd1473311, -32'sd2141212, -32'sd1016510, -32'sd2487829, -32'sd1537062, 32'sd960217, 32'sd1018344, -32'sd1498111, 32'sd623490, 32'sd2026893, 32'sd746673, 32'sd339674, -32'sd1168374, 32'sd1273494, 32'sd173467, -32'sd1040052, 32'sd839139, 32'sd111793, -32'sd1794299, 32'sd345020, 32'sd9156, 32'sd1696272, -32'sd611216, -32'sd606558, 32'sd22844, -32'sd709962, -32'sd1144318, -32'sd722154, -32'sd3506175, -32'sd737025, -32'sd220229, -32'sd514385, -32'sd750084, 32'sd1356040, 32'sd1165151, -32'sd439620, 32'sd928698, 32'sd1445788, 32'sd219554, -32'sd332491, -32'sd1432392, 32'sd475814, 32'sd466766, 32'sd142905, 32'sd186225, 32'sd489551, 32'sd685130, 32'sd460309, -32'sd469520, -32'sd513821, -32'sd1595597, -32'sd767976, -32'sd830112, -32'sd826188, -32'sd1939436, -32'sd3923824, -32'sd3822460, -32'sd1100229, -32'sd91196, 32'sd880564, 32'sd1007908, 32'sd38088, 32'sd1958743, -32'sd1800816, 32'sd371511, 32'sd1682247, 32'sd2006094, -32'sd1694445, -32'sd1373963, -32'sd122896, 32'sd0, 32'sd1006800, 32'sd969506, 32'sd575747, 32'sd840042, -32'sd414670, -32'sd1021323, 32'sd116915, 32'sd214104, -32'sd564824, -32'sd2956056, -32'sd3682300, -32'sd2959498, -32'sd2477077, 32'sd926, 32'sd2249078, 32'sd2913061, 32'sd2095969, 32'sd1524572, -32'sd198110, 32'sd12113, -32'sd464914, -32'sd635246, -32'sd114758, -32'sd1077229, -32'sd133831, -32'sd596085, 32'sd622489, -32'sd161442, -32'sd1469871, -32'sd782116, 32'sd1931877, 32'sd621490, -32'sd720121, 32'sd518158, 32'sd1043705, -32'sd1781461, -32'sd1467378, -32'sd1266540, -32'sd1380484, -32'sd1741129, -32'sd702433, 32'sd2947128, 32'sd4006352, 32'sd1094671, -32'sd1004914, -32'sd784310, -32'sd1070861, -32'sd1397400, -32'sd1754944, -32'sd417493, -32'sd2309389, -32'sd2323290, 32'sd1718967, 32'sd1070958, 32'sd421254, -32'sd303948, -32'sd158965, -32'sd1413304, 32'sd632901, 32'sd1727742, 32'sd819046, -32'sd185926, -32'sd1074326, -32'sd791750, -32'sd332801, -32'sd776957, 32'sd831501, 32'sd160404, -32'sd729190, 32'sd1902352, 32'sd1473467, 32'sd851446, 32'sd971823, 32'sd1353557, 32'sd948809, 32'sd11708, -32'sd304281, -32'sd152043, 32'sd39224, -32'sd716408, 32'sd569595, 32'sd1422319, 32'sd140765, 32'sd0, 32'sd795662, -32'sd585053, 32'sd301890, -32'sd1302008, -32'sd908685, 32'sd224328, -32'sd1437802, -32'sd666178, 32'sd86693, 32'sd1288376, 32'sd868585, 32'sd44591, 32'sd697219, 32'sd2261899, 32'sd2779957, 32'sd650717, 32'sd1063155, -32'sd380814, -32'sd30865, -32'sd1465885, -32'sd1742873, -32'sd9647, 32'sd1432515, 32'sd596870, 32'sd1183840, 32'sd1415484, 32'sd0, 32'sd0, 32'sd0, -32'sd433042, 32'sd977663, -32'sd738767, 32'sd1042703, -32'sd598664, 32'sd1843005, 32'sd2366765, 32'sd1575549, 32'sd2005093, 32'sd1394428, 32'sd2695473, 32'sd1398567, 32'sd3406119, 32'sd1616107, 32'sd778973, 32'sd1239929, 32'sd1619775, 32'sd384151, -32'sd162760, 32'sd739578, 32'sd1790254, -32'sd72531, 32'sd243525, 32'sd437381, -32'sd296167, 32'sd0, 32'sd0, 32'sd0, -32'sd101239, 32'sd380418, -32'sd970919, -32'sd259251, 32'sd365491, 32'sd1935460, 32'sd3346761, 32'sd3118664, 32'sd2410219, 32'sd473105, 32'sd3080243, -32'sd1511221, -32'sd1622540, 32'sd1601819, 32'sd43036, -32'sd766661, -32'sd440898, 32'sd1242193, 32'sd927768, 32'sd377189, 32'sd60168, 32'sd112492, 32'sd1608822, -32'sd128567, -32'sd97667, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd799111, -32'sd1598000, 32'sd414751, -32'sd1485619, 32'sd43988, -32'sd1847815, -32'sd864814, 32'sd759652, -32'sd887212, -32'sd596689, 32'sd879491, -32'sd155417, 32'sd2411651, 32'sd1252460, -32'sd629178, -32'sd1500041, 32'sd677606, 32'sd1344538, 32'sd297681, -32'sd485905, 32'sd428209, 32'sd483542, 32'sd718692, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd530821, 32'sd484067, 32'sd481627, 32'sd963422, -32'sd417041, -32'sd142983, 32'sd852547, 32'sd1236685, -32'sd572214, -32'sd731931, -32'sd322358, 32'sd1253597, 32'sd1192194, 32'sd958017, -32'sd225919, -32'sd391503, -32'sd1646442, -32'sd362509, 32'sd1443466, -32'sd1132625, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1759052, 32'sd1785, -32'sd114363, 32'sd755265, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd321926, -32'sd685702, -32'sd442221, 32'sd1988063, 32'sd1526213, 32'sd405963, 32'sd1027788, -32'sd1265180, 32'sd294919, -32'sd412187, -32'sd1374370, -32'sd174044, 32'sd6305, -32'sd235347, 32'sd2068057, 32'sd1323848, 32'sd89821, 32'sd1910271, 32'sd1432103, 32'sd1420714, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd753384, 32'sd241504, 32'sd933481, 32'sd461467, -32'sd1062776, 32'sd1624828, 32'sd1412658, 32'sd1842643, -32'sd1143113, -32'sd856915, -32'sd823898, -32'sd564187, -32'sd459430, 32'sd1946247, 32'sd1083471, 32'sd1524405, -32'sd605756, -32'sd181376, 32'sd740709, 32'sd1381623, -32'sd207098, 32'sd495227, 32'sd1146469, 32'sd1626984, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd84553, 32'sd351951, -32'sd1571807, -32'sd68148, 32'sd313800, -32'sd300439, 32'sd2799842, -32'sd1341420, -32'sd440612, 32'sd1935737, -32'sd473359, 32'sd792998, 32'sd843782, -32'sd268963, 32'sd1995887, 32'sd471118, -32'sd848268, -32'sd647580, -32'sd2026850, -32'sd298171, -32'sd695498, 32'sd650399, 32'sd264216, 32'sd449488, 32'sd250712, 32'sd0, 32'sd0, 32'sd319388, 32'sd246614, 32'sd1798374, -32'sd1412772, -32'sd839078, -32'sd47798, 32'sd790685, 32'sd1824921, 32'sd1819272, -32'sd34987, -32'sd420248, 32'sd125739, 32'sd667477, -32'sd340098, 32'sd1745806, -32'sd306929, 32'sd268655, -32'sd312652, -32'sd883574, -32'sd1520011, -32'sd97507, -32'sd1319871, -32'sd1717908, -32'sd516284, 32'sd457608, 32'sd766060, -32'sd120368, 32'sd0, 32'sd1365069, 32'sd638941, 32'sd543379, 32'sd293780, -32'sd239593, -32'sd2009007, -32'sd794887, -32'sd1672985, 32'sd822369, -32'sd511422, 32'sd2646955, -32'sd636768, 32'sd340175, 32'sd3162407, 32'sd1298231, 32'sd79029, 32'sd234205, -32'sd2413409, 32'sd14543, 32'sd190068, -32'sd2456384, -32'sd1446329, -32'sd1569748, -32'sd1063403, -32'sd1990578, -32'sd905006, 32'sd1379270, 32'sd0, 32'sd677160, -32'sd364872, 32'sd408716, 32'sd1059377, 32'sd1248064, 32'sd264213, 32'sd78179, 32'sd501049, -32'sd435244, 32'sd1023441, 32'sd2043225, 32'sd94386, 32'sd1357378, 32'sd1878074, 32'sd3159896, -32'sd292980, -32'sd2809338, -32'sd1325952, -32'sd2257978, 32'sd438387, -32'sd1484711, -32'sd2411831, -32'sd2441980, -32'sd1590486, -32'sd1983851, 32'sd1706324, 32'sd886956, 32'sd383985, 32'sd245382, -32'sd1213279, -32'sd1093202, 32'sd170715, 32'sd825466, 32'sd1361125, -32'sd1109907, -32'sd802146, -32'sd2075167, 32'sd842545, 32'sd1311683, -32'sd416073, 32'sd2148186, 32'sd2027535, 32'sd545692, -32'sd2052160, -32'sd3364072, -32'sd1454141, -32'sd2280994, 32'sd122645, -32'sd1292279, 32'sd202471, -32'sd2030964, -32'sd1802928, -32'sd2108543, 32'sd313008, -32'sd317329, 32'sd427764, 32'sd421166, 32'sd1441634, 32'sd991714, 32'sd426079, -32'sd1056246, -32'sd1116113, -32'sd1603452, -32'sd2410827, -32'sd2040676, -32'sd362765, 32'sd1656969, 32'sd1926484, 32'sd1364848, 32'sd224494, -32'sd3180937, -32'sd725353, -32'sd1521786, -32'sd1930562, 32'sd465787, -32'sd1163407, -32'sd755825, -32'sd1099526, -32'sd2763566, 32'sd124305, -32'sd7079, 32'sd1607188, 32'sd959000, 32'sd1575611, 32'sd821509, 32'sd1008545, 32'sd665285, -32'sd1561182, 32'sd31276, 32'sd396488, -32'sd1399781, -32'sd890765, 32'sd1817341, -32'sd182668, 32'sd2026744, 32'sd1551501, 32'sd1328537, -32'sd840687, -32'sd3804520, -32'sd1332842, 32'sd258580, -32'sd238785, -32'sd1260952, 32'sd710842, 32'sd1161626, -32'sd112357, -32'sd2678188, -32'sd2102724, 32'sd468475, 32'sd309990, 32'sd158990, -32'sd528911, 32'sd108079, -32'sd387899, 32'sd714210, -32'sd186155, -32'sd1630188, -32'sd1231962, 32'sd301340, 32'sd1968394, 32'sd863802, 32'sd215343, -32'sd234698, 32'sd220462, -32'sd2482644, -32'sd4771666, -32'sd2889465, -32'sd228362, 32'sd323127, 32'sd767463, 32'sd717445, -32'sd378662, 32'sd1301595, 32'sd141589, 32'sd252722, -32'sd2819092, -32'sd1690375, -32'sd163003, 32'sd671046, -32'sd252515, 32'sd1785876, -32'sd901656, -32'sd832442, -32'sd1140080, -32'sd1203083, -32'sd639366, -32'sd1263915, 32'sd890408, 32'sd594590, 32'sd1159145, 32'sd37322, 32'sd322639, -32'sd2926897, -32'sd5184347, -32'sd1175454, 32'sd670567, 32'sd300714, -32'sd40048, -32'sd467805, 32'sd199634, 32'sd1995825, -32'sd1154277, -32'sd345186, -32'sd984328, -32'sd280721, 32'sd412132, -32'sd560601, 32'sd256526, 32'sd227136, -32'sd399195, 32'sd465847, -32'sd388998, 32'sd1535844, 32'sd350975, 32'sd1650341, -32'sd141566, 32'sd539484, 32'sd643874, -32'sd656372, -32'sd1821783, -32'sd2516827, -32'sd1699428, 32'sd2301699, 32'sd1328351, 32'sd2209054, 32'sd1274599, 32'sd1042541, 32'sd1731395, 32'sd2856542, 32'sd202861, 32'sd1718637, 32'sd654217, -32'sd1185715, 32'sd1088467, -32'sd332446, 32'sd368055, -32'sd522904, -32'sd1138270, -32'sd572664, -32'sd457763, -32'sd441140, 32'sd1646997, 32'sd3324750, 32'sd1872564, -32'sd809225, 32'sd1598093, -32'sd1463164, -32'sd722059, -32'sd1442060, 32'sd504850, 32'sd480727, 32'sd1186268, 32'sd310578, -32'sd73862, 32'sd1571640, -32'sd124444, 32'sd1380394, 32'sd1772517, 32'sd1377715, 32'sd562889, -32'sd658551, -32'sd454745, 32'sd49926, -32'sd1043028, -32'sd240651, -32'sd39976, -32'sd230076, 32'sd62476, 32'sd2149567, -32'sd55960, 32'sd1123767, 32'sd1401383, 32'sd1889321, -32'sd211426, -32'sd224322, -32'sd1157507, -32'sd1285947, -32'sd1412667, 32'sd2909976, 32'sd2344029, -32'sd1065107, 32'sd1564847, 32'sd321079, -32'sd56150, -32'sd162317, 32'sd843029, 32'sd1150296, 32'sd1189255, -32'sd1641366, -32'sd337117, -32'sd526523, 32'sd194679, 32'sd1041074, 32'sd368195, -32'sd611458, -32'sd2098502, 32'sd1108589, 32'sd1132818, 32'sd2997357, 32'sd983314, -32'sd78684, 32'sd2019444, 32'sd1905916, -32'sd533791, -32'sd1808562, -32'sd1533985, -32'sd356808, 32'sd816615, -32'sd336998, 32'sd754748, -32'sd146502, -32'sd92854, -32'sd132266, 32'sd1739194, 32'sd1735034, 32'sd1323421, 32'sd356098, -32'sd2295706, 32'sd527739, 32'sd656952, -32'sd1343175, -32'sd604368, -32'sd547792, -32'sd1246122, -32'sd809325, 32'sd145070, 32'sd1669615, 32'sd1651830, 32'sd1449904, 32'sd1645812, 32'sd1709616, 32'sd1369733, 32'sd224244, -32'sd443779, -32'sd225995, -32'sd3873587, -32'sd2159557, -32'sd697945, -32'sd149466, 32'sd186400, -32'sd1301938, -32'sd166886, 32'sd471468, 32'sd2056748, -32'sd538680, -32'sd405429, 32'sd554576, 32'sd0, 32'sd1250472, 32'sd42434, -32'sd932743, 32'sd515765, -32'sd97844, -32'sd243087, 32'sd1163397, 32'sd1586553, 32'sd1470471, 32'sd1489063, 32'sd1977477, 32'sd1082356, 32'sd1464861, 32'sd1512012, -32'sd2291689, -32'sd2830394, -32'sd2450318, -32'sd2151383, 32'sd901916, 32'sd1568649, -32'sd251424, 32'sd1722834, 32'sd2086597, 32'sd1455089, -32'sd903515, -32'sd1779127, -32'sd899127, 32'sd391321, -32'sd601412, 32'sd373431, -32'sd565847, -32'sd727589, 32'sd1129426, -32'sd1269425, -32'sd1452060, 32'sd941103, 32'sd1504502, 32'sd1857987, 32'sd4992206, 32'sd4099524, 32'sd941880, -32'sd1498046, 32'sd214821, -32'sd1146908, -32'sd2646084, -32'sd16148, 32'sd1457692, 32'sd626722, -32'sd641098, 32'sd1869929, 32'sd655099, 32'sd441204, -32'sd1378290, 32'sd197367, 32'sd612213, 32'sd618373, -32'sd79283, 32'sd108487, 32'sd283564, -32'sd890632, -32'sd997841, -32'sd1698343, -32'sd1405156, -32'sd2573618, -32'sd661531, 32'sd848462, 32'sd2476292, 32'sd3730065, 32'sd1105605, -32'sd933723, 32'sd404861, -32'sd552930, 32'sd567037, 32'sd1294322, 32'sd1034130, 32'sd703735, 32'sd1290446, 32'sd444330, -32'sd986134, 32'sd256478, -32'sd1912338, 32'sd703334, -32'sd1444893, 32'sd0, 32'sd107245, 32'sd597757, 32'sd717827, -32'sd21770, 32'sd6013, -32'sd1591085, -32'sd546244, -32'sd1641436, -32'sd1702101, -32'sd964270, 32'sd107716, 32'sd1219, 32'sd1391889, 32'sd1029365, 32'sd1825193, 32'sd600890, 32'sd787215, 32'sd185844, 32'sd1058081, -32'sd29424, 32'sd1710118, 32'sd1114390, -32'sd422167, 32'sd64324, -32'sd123182, 32'sd1008629, 32'sd628512, 32'sd241838, -32'sd168156, -32'sd1277783, 32'sd890305, 32'sd244150, -32'sd376729, 32'sd1096720, -32'sd689171, -32'sd1130153, -32'sd1951143, -32'sd1934373, -32'sd1577737, -32'sd749934, -32'sd1194435, 32'sd3140728, 32'sd3449693, 32'sd1008920, 32'sd1133876, 32'sd1000559, -32'sd1118419, 32'sd736873, 32'sd351607, 32'sd470738, -32'sd887754, -32'sd1821943, -32'sd942706, 32'sd346941, 32'sd365925, 32'sd338776, -32'sd798075, -32'sd1000314, -32'sd832784, -32'sd627151, 32'sd692576, 32'sd491624, -32'sd37039, -32'sd596076, 32'sd25973, -32'sd3021333, -32'sd2206811, -32'sd808786, 32'sd785238, 32'sd1545018, 32'sd1102598, 32'sd2319191, 32'sd1243624, -32'sd315935, -32'sd184680, -32'sd51525, 32'sd1365370, -32'sd663099, -32'sd2398465, -32'sd1655190, -32'sd1594272, 32'sd1464434, 32'sd333958, 32'sd0, -32'sd571754, 32'sd575911, 32'sd235309, -32'sd17878, 32'sd172588, -32'sd198019, 32'sd667741, -32'sd921155, -32'sd234638, 32'sd550326, -32'sd653823, -32'sd1445811, -32'sd83561, 32'sd2584997, -32'sd896276, -32'sd1312955, 32'sd265495, -32'sd106209, 32'sd503303, 32'sd1390911, 32'sd95086, -32'sd388166, -32'sd1215711, -32'sd1778564, -32'sd542779, 32'sd715693, 32'sd0, 32'sd0, 32'sd0, -32'sd85699, 32'sd607494, -32'sd416800, -32'sd406671, 32'sd1436831, 32'sd1057850, 32'sd381666, 32'sd282495, -32'sd274259, -32'sd241548, -32'sd428863, 32'sd3333183, 32'sd588908, 32'sd628492, 32'sd2924915, 32'sd8635, 32'sd626063, -32'sd887109, -32'sd1607250, 32'sd433426, -32'sd886370, 32'sd1593063, -32'sd334012, 32'sd547820, 32'sd183203, 32'sd0, 32'sd0, 32'sd0, -32'sd903424, -32'sd918030, 32'sd69221, 32'sd439009, -32'sd1080058, 32'sd237469, 32'sd2079637, 32'sd723966, -32'sd291324, 32'sd87326, 32'sd263166, 32'sd1824372, 32'sd538301, -32'sd187623, -32'sd246136, -32'sd287593, -32'sd50242, 32'sd1416321, -32'sd443477, -32'sd139512, -32'sd320542, 32'sd2118479, -32'sd76009, 32'sd605686, 32'sd892038, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd644441, 32'sd260571, -32'sd145863, -32'sd1330269, 32'sd189318, 32'sd752751, -32'sd1553370, -32'sd2647503, -32'sd1112246, -32'sd747177, -32'sd1972787, 32'sd181880, -32'sd1079186, 32'sd906103, -32'sd1434138, -32'sd1357910, 32'sd1040321, 32'sd1538107, -32'sd308495, -32'sd2120102, -32'sd1594353, -32'sd180543, 32'sd1285053, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1725923, 32'sd59199, 32'sd989332, 32'sd1449627, 32'sd1526985, -32'sd104453, 32'sd1096093, 32'sd278270, 32'sd1415074, -32'sd474032, -32'sd708381, -32'sd784236, 32'sd136365, 32'sd310332, 32'sd122660, -32'sd167874, 32'sd226027, -32'sd683571, 32'sd183331, 32'sd1169707, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd132268, -32'sd90549, -32'sd158403, 32'sd1144127, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1213200, 32'sd484632, 32'sd693014, 32'sd1628875, -32'sd350521, -32'sd1107208, -32'sd600165, -32'sd146501, 32'sd617097, -32'sd633126, -32'sd348023, 32'sd180486, -32'sd397292, 32'sd1180910, 32'sd341423, 32'sd751378, -32'sd514723, 32'sd1820477, 32'sd809548, 32'sd647437, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1883225, 32'sd994495, 32'sd1573552, -32'sd264227, -32'sd208779, 32'sd607356, 32'sd1690504, 32'sd1097875, -32'sd133758, -32'sd567128, -32'sd2019897, -32'sd154833, -32'sd2275290, -32'sd613131, 32'sd536782, 32'sd3116638, 32'sd3102183, 32'sd304562, 32'sd1164745, -32'sd1285855, 32'sd1080430, 32'sd1006094, 32'sd1385095, 32'sd1186558, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1311238, 32'sd421804, -32'sd272403, 32'sd738129, 32'sd2329378, -32'sd205778, 32'sd1018794, 32'sd309420, -32'sd921738, -32'sd618264, -32'sd1304937, 32'sd1483806, 32'sd406206, 32'sd41004, 32'sd1426530, -32'sd931143, 32'sd1313679, 32'sd604770, -32'sd787501, 32'sd1177747, -32'sd168539, 32'sd428253, -32'sd1284498, 32'sd1554485, -32'sd550698, 32'sd0, 32'sd0, 32'sd1226835, 32'sd355511, 32'sd487008, 32'sd1091940, 32'sd666959, 32'sd1214846, 32'sd811650, -32'sd327169, -32'sd1351427, 32'sd57585, 32'sd79336, 32'sd106853, -32'sd1805039, 32'sd1383008, 32'sd965511, 32'sd118738, 32'sd1028782, 32'sd1488142, 32'sd1090260, 32'sd1569754, 32'sd1025316, -32'sd1870653, 32'sd1225750, 32'sd1829068, -32'sd547228, 32'sd413808, 32'sd10543, 32'sd0, 32'sd593269, 32'sd436147, -32'sd2221313, -32'sd84773, -32'sd440064, 32'sd214333, -32'sd1627709, 32'sd200752, -32'sd1202239, 32'sd1527098, 32'sd1379965, 32'sd2476346, 32'sd912470, 32'sd1162628, 32'sd2409593, 32'sd3403108, 32'sd2428439, 32'sd3295143, 32'sd1315379, 32'sd1611011, 32'sd3099005, 32'sd1579687, 32'sd2103152, 32'sd2839093, -32'sd924096, -32'sd734522, 32'sd1003098, 32'sd0, 32'sd318540, -32'sd443911, -32'sd1193986, 32'sd326055, -32'sd1095102, -32'sd616570, 32'sd1579903, 32'sd1670858, -32'sd481355, 32'sd965814, 32'sd3614888, 32'sd1262159, 32'sd911379, 32'sd973913, 32'sd3651519, 32'sd3043461, 32'sd2442475, 32'sd2422559, 32'sd2668806, 32'sd731944, 32'sd54261, 32'sd34380, 32'sd21853, 32'sd2458383, -32'sd291797, -32'sd672504, 32'sd220006, 32'sd455444, 32'sd1996457, -32'sd889514, -32'sd1124128, -32'sd441568, 32'sd1152086, 32'sd1041703, -32'sd481078, 32'sd738018, 32'sd413472, 32'sd526156, 32'sd1334847, 32'sd1204818, 32'sd248511, 32'sd2225314, 32'sd282995, 32'sd1649044, -32'sd387517, -32'sd324950, -32'sd703376, -32'sd2239374, -32'sd1357761, -32'sd281160, -32'sd3356461, -32'sd1883155, 32'sd667153, 32'sd325966, 32'sd999181, 32'sd1297426, 32'sd516895, -32'sd16878, -32'sd408536, -32'sd355545, -32'sd920267, 32'sd298930, -32'sd384473, 32'sd436330, 32'sd47221, 32'sd737403, 32'sd1421675, 32'sd1207438, -32'sd386752, 32'sd959481, -32'sd2721429, -32'sd3427506, -32'sd2312618, -32'sd657843, -32'sd2198372, -32'sd3605488, -32'sd1799233, -32'sd363192, -32'sd3365548, -32'sd3039469, -32'sd1329829, 32'sd337095, -32'sd212908, 32'sd432203, -32'sd498554, -32'sd124127, -32'sd87766, -32'sd322856, -32'sd457194, 32'sd1928677, -32'sd74133, 32'sd459790, -32'sd264893, 32'sd1474920, -32'sd910063, -32'sd994555, -32'sd151131, -32'sd1260465, -32'sd3567481, -32'sd4208188, -32'sd1277750, -32'sd1474918, -32'sd3824861, -32'sd2973472, -32'sd1436163, -32'sd1910297, -32'sd4992498, -32'sd994919, -32'sd1085006, -32'sd528267, 32'sd581528, 32'sd244121, -32'sd1712905, -32'sd929310, -32'sd1374120, -32'sd614343, 32'sd1230326, 32'sd2286425, -32'sd7757, 32'sd168927, 32'sd1812, -32'sd1254695, -32'sd1952482, -32'sd2235224, -32'sd2464734, -32'sd4357100, -32'sd3571074, -32'sd3925786, -32'sd4452881, -32'sd2531643, -32'sd2869514, -32'sd1980557, -32'sd2149151, -32'sd3628527, -32'sd786652, -32'sd2386834, -32'sd1147494, -32'sd1008083, -32'sd38643, 32'sd277962, -32'sd287195, 32'sd581906, -32'sd99850, 32'sd1535511, 32'sd286950, 32'sd1062102, -32'sd978292, -32'sd1071980, -32'sd2136212, -32'sd318271, -32'sd2936284, -32'sd161126, -32'sd2685524, -32'sd1648970, 32'sd566844, -32'sd1837244, -32'sd631755, -32'sd445033, -32'sd2796891, -32'sd2711930, 32'sd46692, 32'sd142709, -32'sd839837, 32'sd730894, -32'sd713133, -32'sd497112, -32'sd281893, 32'sd425666, 32'sd759442, -32'sd982434, 32'sd2217751, -32'sd208636, 32'sd101868, -32'sd754652, -32'sd1894106, -32'sd976122, -32'sd1142057, -32'sd957675, -32'sd1515292, -32'sd1342329, -32'sd3130611, -32'sd350907, 32'sd1627092, 32'sd742326, 32'sd1235944, -32'sd689162, 32'sd867634, 32'sd711283, -32'sd789069, -32'sd567036, 32'sd1151354, 32'sd1835207, -32'sd1077735, -32'sd1891733, -32'sd361459, 32'sd333624, -32'sd1672047, -32'sd99406, 32'sd288228, -32'sd289459, -32'sd1628738, -32'sd42360, 32'sd1269176, 32'sd513827, -32'sd951004, 32'sd333412, 32'sd419911, -32'sd1307931, -32'sd1087873, 32'sd971472, 32'sd124824, 32'sd1224124, 32'sd1191906, 32'sd1235824, 32'sd3219662, 32'sd3732155, -32'sd1501730, -32'sd1249646, 32'sd125039, 32'sd1080397, 32'sd75526, 32'sd173136, -32'sd160339, 32'sd2130480, 32'sd1078451, 32'sd195735, 32'sd863551, 32'sd825902, 32'sd999389, 32'sd474051, -32'sd412579, -32'sd149949, -32'sd852405, 32'sd1571431, 32'sd1313409, -32'sd1286568, -32'sd840541, 32'sd30915, -32'sd1060715, 32'sd371248, 32'sd187188, 32'sd1259450, 32'sd2044167, 32'sd1749233, 32'sd73479, -32'sd1358380, -32'sd586722, 32'sd699146, -32'sd815477, -32'sd264234, 32'sd461469, 32'sd862401, 32'sd181091, 32'sd385063, 32'sd76958, -32'sd839914, -32'sd180951, 32'sd2267930, 32'sd1526387, 32'sd1938293, 32'sd84488, -32'sd1761779, -32'sd2213538, -32'sd1563937, -32'sd538706, -32'sd357731, -32'sd1819878, 32'sd231297, 32'sd926548, 32'sd516185, 32'sd1467878, 32'sd1404095, 32'sd491496, -32'sd2462573, 32'sd945872, 32'sd248092, 32'sd1446577, 32'sd640060, -32'sd912229, 32'sd1159164, 32'sd1353249, -32'sd663695, 32'sd1293694, 32'sd1438244, -32'sd111381, -32'sd927660, 32'sd32332, -32'sd727667, -32'sd784857, -32'sd527682, -32'sd1033215, 32'sd449833, 32'sd1029839, -32'sd110835, 32'sd1389331, 32'sd1548158, 32'sd1615750, 32'sd1785795, 32'sd578647, 32'sd667585, -32'sd342934, -32'sd657173, 32'sd1501196, -32'sd1045553, 32'sd617658, -32'sd743442, 32'sd585602, 32'sd0, -32'sd387805, 32'sd133538, 32'sd1277873, 32'sd1005746, -32'sd458778, -32'sd886254, -32'sd2547169, -32'sd1042718, 32'sd275205, 32'sd307003, 32'sd221419, 32'sd2369765, -32'sd228715, -32'sd794496, 32'sd1135796, 32'sd2001851, -32'sd407941, -32'sd379226, 32'sd43606, 32'sd164759, 32'sd675540, 32'sd841547, -32'sd1128273, -32'sd1224132, 32'sd248960, -32'sd1694667, 32'sd989306, 32'sd969660, 32'sd1315042, 32'sd138948, -32'sd14383, 32'sd296833, 32'sd1585297, 32'sd1411867, -32'sd2650092, -32'sd1218096, -32'sd1760309, 32'sd2016597, 32'sd2557394, 32'sd1663032, 32'sd346268, 32'sd596195, 32'sd1502023, 32'sd747873, -32'sd50363, -32'sd134974, 32'sd307685, -32'sd623471, -32'sd891339, 32'sd1132637, 32'sd100039, -32'sd43883, 32'sd812463, -32'sd308499, 32'sd1179671, 32'sd1009431, 32'sd760381, 32'sd30013, -32'sd686548, 32'sd94314, 32'sd863332, 32'sd37353, -32'sd1654446, -32'sd575724, -32'sd272699, 32'sd3328828, 32'sd2755401, 32'sd2310801, 32'sd1035022, -32'sd400507, -32'sd749339, 32'sd608284, 32'sd429521, 32'sd2262738, 32'sd206102, -32'sd1007291, -32'sd1606656, 32'sd827618, 32'sd703975, 32'sd420530, 32'sd2142001, 32'sd1643558, -32'sd881965, 32'sd0, -32'sd1229078, 32'sd1074147, -32'sd247619, 32'sd2935746, 32'sd1217196, 32'sd1686433, -32'sd302927, -32'sd1419904, 32'sd1591169, 32'sd955055, -32'sd12952, 32'sd2085485, 32'sd379599, -32'sd232829, -32'sd386581, -32'sd814288, 32'sd562249, 32'sd1035469, -32'sd225957, -32'sd592899, 32'sd421884, 32'sd979353, 32'sd1593017, 32'sd894901, 32'sd559539, -32'sd1156526, 32'sd601905, 32'sd1732112, 32'sd795245, -32'sd1142008, 32'sd1127488, 32'sd1704262, 32'sd769480, 32'sd2341865, -32'sd893398, 32'sd590719, 32'sd1689052, 32'sd1229827, 32'sd1725265, 32'sd1918916, 32'sd1247724, -32'sd6534, 32'sd1949390, 32'sd1790811, 32'sd230816, 32'sd1096671, 32'sd406321, -32'sd513856, 32'sd35231, -32'sd180005, 32'sd1257527, 32'sd1293122, -32'sd854225, -32'sd724583, 32'sd1180457, -32'sd84951, -32'sd89940, -32'sd726384, 32'sd784990, 32'sd1161399, 32'sd1191335, -32'sd903999, -32'sd178090, 32'sd470720, 32'sd1384532, -32'sd492234, -32'sd462503, 32'sd1503111, -32'sd147741, 32'sd1001527, -32'sd436223, -32'sd1213482, -32'sd1996795, 32'sd410298, -32'sd1131538, -32'sd670150, 32'sd480526, 32'sd1385074, 32'sd1673172, 32'sd192038, 32'sd684248, -32'sd407236, 32'sd615004, 32'sd0, 32'sd620026, -32'sd1473531, -32'sd388600, -32'sd255651, 32'sd1487917, -32'sd1579892, 32'sd342431, 32'sd882121, -32'sd1313550, -32'sd259825, -32'sd2424617, 32'sd137677, -32'sd865240, -32'sd618295, -32'sd19022, -32'sd1202260, -32'sd1421486, -32'sd1078154, -32'sd284035, 32'sd105412, 32'sd1323870, 32'sd832450, 32'sd1386461, 32'sd1248728, 32'sd1524033, -32'sd459596, 32'sd0, 32'sd0, 32'sd0, -32'sd454126, -32'sd392849, -32'sd386667, 32'sd430268, -32'sd1634506, -32'sd545563, -32'sd620176, 32'sd212011, 32'sd324755, -32'sd1019653, -32'sd1916383, 32'sd76713, -32'sd195942, -32'sd431961, -32'sd614005, 32'sd264093, 32'sd1708573, 32'sd588305, 32'sd1268844, 32'sd1201242, -32'sd241722, -32'sd281012, 32'sd694125, -32'sd457762, 32'sd445834, 32'sd0, 32'sd0, 32'sd0, 32'sd1553536, 32'sd631690, -32'sd1525205, 32'sd396016, -32'sd1401528, -32'sd558039, -32'sd2094864, -32'sd2276032, -32'sd994821, -32'sd204332, 32'sd992059, -32'sd1770990, 32'sd552838, -32'sd1308362, 32'sd780207, 32'sd179407, 32'sd746985, 32'sd943972, 32'sd826139, -32'sd59532, 32'sd587732, 32'sd1786648, 32'sd1509655, 32'sd838204, 32'sd426501, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd622141, 32'sd25181, -32'sd228363, -32'sd859873, 32'sd714037, 32'sd1594625, -32'sd240092, 32'sd1015169, 32'sd146491, 32'sd23668, -32'sd352045, 32'sd58611, -32'sd337101, -32'sd1197975, -32'sd83422, 32'sd785463, 32'sd1382348, 32'sd1931800, 32'sd197409, 32'sd418620, 32'sd511196, 32'sd2270306, 32'sd841082, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd535232, 32'sd1595692, -32'sd6895, 32'sd908265, 32'sd100778, -32'sd108991, 32'sd1134364, 32'sd1010468, 32'sd90808, 32'sd614585, 32'sd1877676, 32'sd1008714, 32'sd650267, -32'sd785710, 32'sd269009, -32'sd31841, 32'sd13518, 32'sd621684, 32'sd538523, -32'sd314355, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd456730, -32'sd1494461, -32'sd26119, 32'sd554422, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd96700, -32'sd396524, -32'sd215597, 32'sd41297, -32'sd1512199, -32'sd353005, 32'sd361927, -32'sd1808610, -32'sd1323888, -32'sd535903, 32'sd298359, -32'sd2093344, 32'sd1436129, 32'sd393128, 32'sd1420524, 32'sd1707256, -32'sd732029, 32'sd1287014, 32'sd393970, 32'sd137792, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd471751, -32'sd768914, 32'sd410375, 32'sd498855, -32'sd658349, 32'sd280719, -32'sd1072047, -32'sd616710, -32'sd2109941, 32'sd599440, -32'sd2531342, -32'sd1177666, 32'sd471246, 32'sd1103446, -32'sd449492, 32'sd2968607, 32'sd1046437, 32'sd1506109, -32'sd182081, 32'sd1570688, 32'sd1892615, -32'sd192925, 32'sd323616, -32'sd738883, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd348683, -32'sd310220, 32'sd1390083, -32'sd1550057, -32'sd868276, 32'sd65056, 32'sd1103474, -32'sd2014968, -32'sd1631324, 32'sd156242, -32'sd1913177, -32'sd197745, 32'sd1317974, -32'sd1858826, 32'sd232933, 32'sd813766, 32'sd102235, 32'sd1157621, -32'sd870781, 32'sd1137530, -32'sd24145, 32'sd1325028, 32'sd270439, -32'sd334810, -32'sd678592, 32'sd0, 32'sd0, 32'sd680724, -32'sd1658310, -32'sd715905, -32'sd501045, 32'sd1061784, -32'sd135608, -32'sd247648, -32'sd2969709, -32'sd2804899, -32'sd2927071, -32'sd559136, -32'sd777336, -32'sd188255, 32'sd1255624, 32'sd952406, 32'sd1673819, 32'sd1882282, 32'sd1575052, -32'sd368038, 32'sd342712, 32'sd1603302, -32'sd644439, -32'sd10245, -32'sd772101, -32'sd484886, 32'sd349120, -32'sd502295, 32'sd0, -32'sd1008069, 32'sd1398777, 32'sd76852, -32'sd1414540, -32'sd1304251, -32'sd1746187, -32'sd3382848, -32'sd2142510, -32'sd1449136, -32'sd1892547, 32'sd999164, 32'sd233894, -32'sd2018504, -32'sd1533764, -32'sd773330, -32'sd428190, 32'sd118231, 32'sd860649, 32'sd2095141, -32'sd51004, -32'sd1793421, -32'sd1661506, -32'sd1538004, -32'sd997339, -32'sd522401, -32'sd526372, 32'sd262851, 32'sd0, -32'sd983377, 32'sd561171, 32'sd238738, -32'sd1560473, -32'sd2093392, -32'sd1510708, -32'sd1693041, -32'sd3022782, -32'sd2178483, -32'sd306697, -32'sd952436, -32'sd1574726, 32'sd483315, 32'sd2435822, 32'sd2548830, 32'sd304713, 32'sd594701, 32'sd1566952, 32'sd1852086, 32'sd2072281, 32'sd470609, -32'sd2110779, -32'sd1804482, -32'sd1965968, 32'sd985945, -32'sd559523, 32'sd847521, -32'sd368139, -32'sd1188405, -32'sd59798, 32'sd125548, -32'sd266444, -32'sd2780711, -32'sd3702084, -32'sd3027987, -32'sd3726759, -32'sd2882589, 32'sd946681, -32'sd772011, -32'sd49172, 32'sd1230070, 32'sd2462237, 32'sd2378783, -32'sd208044, -32'sd1170496, 32'sd658655, -32'sd458324, 32'sd2283101, 32'sd2513505, -32'sd638011, -32'sd2215667, 32'sd326044, 32'sd235751, -32'sd529220, -32'sd1156984, -32'sd463218, 32'sd618908, 32'sd1693717, 32'sd57279, -32'sd2098554, -32'sd4189819, -32'sd2640690, -32'sd2928767, -32'sd2343468, -32'sd1908012, 32'sd366267, 32'sd2227160, 32'sd890076, 32'sd2959640, 32'sd750229, 32'sd476428, 32'sd674140, -32'sd762607, -32'sd20413, -32'sd279561, -32'sd1299911, 32'sd1513354, -32'sd1794542, -32'sd1776129, 32'sd753586, -32'sd1172227, -32'sd242887, -32'sd1206514, -32'sd988851, -32'sd1690671, 32'sd501924, 32'sd1080927, -32'sd2671079, -32'sd2758495, -32'sd3548700, -32'sd3830113, -32'sd1929328, 32'sd831925, 32'sd2806371, 32'sd63995, 32'sd572957, 32'sd2442713, 32'sd1693523, 32'sd529941, 32'sd150464, -32'sd3515129, -32'sd1321340, -32'sd1818140, -32'sd762936, -32'sd1878541, 32'sd63059, 32'sd675425, 32'sd789091, 32'sd1197, -32'sd1120812, -32'sd1678955, 32'sd382573, -32'sd1398337, 32'sd1029726, 32'sd41527, -32'sd2728240, -32'sd2931561, -32'sd2360866, 32'sd31227, -32'sd736168, 32'sd649204, 32'sd729603, -32'sd347706, -32'sd1116160, 32'sd280453, 32'sd2616304, -32'sd1177482, -32'sd1551237, -32'sd1872220, -32'sd2167828, -32'sd3572838, -32'sd203490, -32'sd1055067, -32'sd1647309, 32'sd788712, 32'sd926531, -32'sd309289, -32'sd1104838, -32'sd898751, -32'sd944044, -32'sd1934243, -32'sd948094, -32'sd539450, -32'sd2702327, -32'sd1741700, -32'sd3587025, 32'sd1133133, 32'sd1316005, 32'sd2720137, 32'sd310720, -32'sd1513828, 32'sd407053, 32'sd2196623, -32'sd8731, -32'sd2189443, -32'sd4990894, -32'sd4059354, 32'sd19405, -32'sd2763931, -32'sd467273, -32'sd460481, -32'sd378039, -32'sd342551, 32'sd1159919, 32'sd1900211, 32'sd422108, -32'sd1115510, 32'sd87389, -32'sd481591, -32'sd2235250, 32'sd328283, -32'sd1203966, -32'sd3456855, -32'sd3075385, -32'sd96449, 32'sd1968480, 32'sd337847, -32'sd1050952, 32'sd1403613, 32'sd1037447, -32'sd190852, -32'sd1141548, -32'sd4929559, -32'sd2004886, -32'sd2157645, -32'sd1068416, 32'sd197895, 32'sd1534262, 32'sd2027073, 32'sd600257, 32'sd2642781, 32'sd1848395, -32'sd12683, 32'sd654818, -32'sd1198280, -32'sd195310, -32'sd1199444, -32'sd1414732, 32'sd236799, -32'sd927475, -32'sd2154133, 32'sd862630, 32'sd462420, 32'sd1700312, -32'sd449496, 32'sd83915, 32'sd1142372, 32'sd833848, -32'sd832246, -32'sd2002973, -32'sd693440, 32'sd1222362, 32'sd56754, 32'sd170415, 32'sd2779888, 32'sd1811094, 32'sd231281, 32'sd3316440, 32'sd1831414, -32'sd664169, -32'sd2052575, -32'sd230481, -32'sd1138486, -32'sd556146, -32'sd584902, 32'sd339373, -32'sd817439, -32'sd1229286, 32'sd345094, 32'sd569111, -32'sd55145, 32'sd24967, 32'sd92235, -32'sd747998, -32'sd1203569, -32'sd2098731, -32'sd1615762, 32'sd224545, -32'sd574293, 32'sd3073151, 32'sd720120, 32'sd362518, 32'sd1711366, 32'sd1448080, 32'sd1296010, 32'sd1518079, -32'sd458018, -32'sd930762, -32'sd266917, 32'sd289769, 32'sd380927, -32'sd733277, 32'sd87809, 32'sd1066947, -32'sd1417251, -32'sd2411676, -32'sd271894, -32'sd294306, 32'sd2140958, 32'sd2620382, -32'sd834607, 32'sd1103324, -32'sd1439782, -32'sd1103384, -32'sd280644, 32'sd79923, 32'sd304802, 32'sd1620523, 32'sd40349, -32'sd544654, 32'sd752680, 32'sd793059, -32'sd1525607, 32'sd245881, -32'sd516931, -32'sd1391229, 32'sd632690, -32'sd693304, 32'sd501123, 32'sd72564, 32'sd469427, 32'sd229055, -32'sd1233337, -32'sd2344653, -32'sd784221, -32'sd983372, 32'sd2433739, 32'sd2391017, -32'sd368156, -32'sd404138, 32'sd1026205, -32'sd1201287, -32'sd315239, -32'sd580397, 32'sd726368, -32'sd272110, -32'sd634917, -32'sd230371, -32'sd56025, 32'sd1570217, 32'sd89661, -32'sd1777827, 32'sd883224, -32'sd766951, 32'sd1450002, 32'sd887365, 32'sd393331, 32'sd0, -32'sd1104154, -32'sd111908, 32'sd485343, 32'sd259287, -32'sd37323, 32'sd1210726, 32'sd345312, 32'sd190099, -32'sd118003, -32'sd1709713, -32'sd1884781, 32'sd699784, -32'sd398375, 32'sd696672, -32'sd1929581, -32'sd1120176, 32'sd1060713, -32'sd855339, -32'sd1400006, 32'sd1402576, 32'sd958616, 32'sd1047172, -32'sd628867, 32'sd121992, -32'sd2377035, -32'sd307765, 32'sd940038, -32'sd427603, -32'sd1060659, 32'sd362217, 32'sd777472, -32'sd1925604, -32'sd758086, -32'sd1686262, 32'sd1882981, 32'sd2482557, 32'sd1890478, -32'sd81849, -32'sd1676449, 32'sd1061127, 32'sd820134, -32'sd601683, -32'sd1698227, -32'sd622062, 32'sd2312083, -32'sd1535981, -32'sd235648, 32'sd461053, 32'sd1137312, 32'sd840897, 32'sd1161207, -32'sd80815, 32'sd510036, -32'sd591982, 32'sd154212, -32'sd639172, -32'sd31523, -32'sd861565, -32'sd1345217, -32'sd1030252, 32'sd323605, -32'sd897926, 32'sd2470558, 32'sd3577162, 32'sd2161111, 32'sd2329016, 32'sd217370, -32'sd994666, -32'sd26582, -32'sd265848, -32'sd1268457, -32'sd1695878, -32'sd438544, 32'sd230660, -32'sd1095845, -32'sd1146306, 32'sd2981768, 32'sd4101533, 32'sd3413758, -32'sd97846, -32'sd2066715, -32'sd393109, 32'sd675953, 32'sd0, -32'sd887950, -32'sd666013, -32'sd691470, -32'sd1446954, 32'sd1586824, -32'sd64809, 32'sd142203, 32'sd920894, 32'sd3631037, 32'sd3880269, 32'sd770586, -32'sd1087702, 32'sd692903, -32'sd974699, -32'sd556988, -32'sd1035546, 32'sd906283, -32'sd935388, -32'sd715309, 32'sd2123654, 32'sd2500924, 32'sd2352353, 32'sd1694480, -32'sd739316, 32'sd108059, 32'sd1295174, -32'sd566758, -32'sd27499, 32'sd265476, 32'sd943505, -32'sd476276, 32'sd174753, -32'sd947006, -32'sd1160607, 32'sd586327, 32'sd52122, 32'sd1983915, 32'sd2372946, 32'sd773154, 32'sd732053, 32'sd2655522, 32'sd20363, 32'sd45447, -32'sd278775, -32'sd139539, -32'sd483784, -32'sd406383, 32'sd2150999, 32'sd881338, -32'sd104179, 32'sd1852452, 32'sd1628294, -32'sd1697585, 32'sd411765, -32'sd945826, -32'sd512679, -32'sd502495, -32'sd1120782, 32'sd1857518, 32'sd1564247, 32'sd270832, 32'sd359594, 32'sd357389, -32'sd557022, -32'sd1082290, -32'sd704049, -32'sd1920006, 32'sd2036893, 32'sd2496283, 32'sd2318681, 32'sd3159733, -32'sd153739, -32'sd1613994, -32'sd458516, 32'sd203333, -32'sd1004398, 32'sd1549239, -32'sd1089208, 32'sd1110093, 32'sd968581, -32'sd282141, 32'sd1714389, 32'sd117070, 32'sd0, -32'sd57636, 32'sd1109076, 32'sd374927, 32'sd531835, 32'sd3302570, 32'sd306255, -32'sd877864, -32'sd903442, -32'sd2954355, -32'sd1573175, -32'sd1856792, 32'sd189043, 32'sd1246155, 32'sd617408, 32'sd2294730, 32'sd1344555, 32'sd1702719, 32'sd1600463, -32'sd239367, -32'sd525451, -32'sd2282928, -32'sd327983, -32'sd537870, 32'sd721788, 32'sd65599, 32'sd482231, 32'sd0, 32'sd0, 32'sd0, -32'sd482999, -32'sd1987377, 32'sd187583, 32'sd1352401, -32'sd1315322, -32'sd261661, -32'sd964727, -32'sd1372838, 32'sd913153, -32'sd801584, -32'sd660971, -32'sd2332625, -32'sd1440757, -32'sd243756, 32'sd1599515, -32'sd304193, -32'sd1933041, -32'sd1823241, -32'sd2344120, -32'sd2650826, 32'sd153752, 32'sd1370990, -32'sd705104, 32'sd165145, -32'sd615123, 32'sd0, 32'sd0, 32'sd0, 32'sd1073830, -32'sd1085651, -32'sd1760969, 32'sd1124034, -32'sd1165445, -32'sd2575510, 32'sd516171, 32'sd909899, -32'sd457734, 32'sd912145, -32'sd111712, -32'sd247824, -32'sd1608250, 32'sd280613, 32'sd1030694, 32'sd1124762, -32'sd1992293, 32'sd675410, 32'sd893216, -32'sd1100489, -32'sd954107, 32'sd937547, -32'sd234507, -32'sd831116, -32'sd876925, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd431059, -32'sd853849, -32'sd2088694, -32'sd522239, 32'sd110976, -32'sd945774, -32'sd1940793, 32'sd211012, 32'sd699347, -32'sd1520176, -32'sd3274312, -32'sd3015729, -32'sd2596239, -32'sd1055673, -32'sd2367667, 32'sd424568, -32'sd863248, 32'sd725716, 32'sd1000752, -32'sd1766210, 32'sd951053, -32'sd581750, -32'sd339060, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd17524, 32'sd353936, 32'sd637146, -32'sd70808, -32'sd1186983, 32'sd293263, -32'sd1412597, -32'sd1951914, -32'sd920373, -32'sd1042227, 32'sd913457, 32'sd1030444, -32'sd300508, 32'sd1042183, -32'sd1103171, -32'sd697937, -32'sd1172214, -32'sd708071, 32'sd116879, 32'sd749998, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1314352, 32'sd494126, 32'sd888467, 32'sd1538508, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1651722, 32'sd1136182, 32'sd1088868, 32'sd1186580, 32'sd1929987, 32'sd914925, 32'sd3333172, 32'sd2240159, 32'sd1817628, 32'sd466089, -32'sd444867, 32'sd300478, 32'sd1093017, 32'sd1246815, 32'sd1901704, 32'sd86117, 32'sd1463733, 32'sd1328714, 32'sd2168041, 32'sd1555011, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1094224, 32'sd1214205, -32'sd768727, 32'sd1370330, -32'sd324215, 32'sd53274, -32'sd657473, -32'sd671575, 32'sd477940, 32'sd974055, 32'sd1805852, -32'sd985378, 32'sd1093315, 32'sd2008461, 32'sd2159155, 32'sd964535, 32'sd2196834, -32'sd42441, 32'sd574302, 32'sd1388945, 32'sd823842, 32'sd1510419, 32'sd1696651, 32'sd1454384, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1624578, 32'sd1226040, 32'sd223811, 32'sd1693955, 32'sd761859, 32'sd1333488, 32'sd126334, 32'sd1642857, 32'sd510940, -32'sd710296, -32'sd164949, -32'sd446433, -32'sd378467, 32'sd1632677, 32'sd45705, -32'sd176814, 32'sd220106, -32'sd850023, 32'sd1676293, 32'sd1434620, -32'sd478810, 32'sd224155, 32'sd54764, 32'sd368161, -32'sd603941, 32'sd0, 32'sd0, 32'sd1306945, -32'sd457784, 32'sd647248, -32'sd519584, 32'sd296526, 32'sd1484761, 32'sd1259208, 32'sd1666006, 32'sd706354, 32'sd1529146, 32'sd876610, 32'sd415073, 32'sd169467, 32'sd692681, 32'sd189312, 32'sd1644872, -32'sd1291616, 32'sd954811, -32'sd1079325, 32'sd449061, 32'sd1079671, -32'sd431195, -32'sd1494143, -32'sd607779, 32'sd1099845, -32'sd256467, -32'sd244683, 32'sd0, 32'sd576456, 32'sd392391, 32'sd1207468, 32'sd883154, 32'sd2119269, -32'sd508895, 32'sd960424, 32'sd693059, 32'sd393157, 32'sd1337200, 32'sd1475958, -32'sd850051, 32'sd621894, -32'sd626517, -32'sd1550410, -32'sd1460930, -32'sd1489766, 32'sd1780689, 32'sd146970, 32'sd1055680, 32'sd1382293, 32'sd1439096, -32'sd1290597, -32'sd1022037, 32'sd1048670, 32'sd213134, 32'sd1163080, 32'sd0, 32'sd94663, -32'sd34917, 32'sd1254213, 32'sd79410, 32'sd2375822, 32'sd1444522, 32'sd1753596, 32'sd572626, -32'sd903460, -32'sd31779, 32'sd792874, 32'sd1365681, -32'sd199617, 32'sd191042, -32'sd1085920, -32'sd2067684, -32'sd306931, 32'sd1406242, -32'sd6034, 32'sd1166111, 32'sd118144, 32'sd901191, -32'sd532464, 32'sd1998737, 32'sd1891501, 32'sd1099684, 32'sd390008, 32'sd1319371, 32'sd1175011, 32'sd250340, -32'sd318351, 32'sd1216397, 32'sd1499285, 32'sd1456319, 32'sd944597, 32'sd892912, 32'sd51010, 32'sd1902839, 32'sd1275400, 32'sd1871754, 32'sd635855, 32'sd1627705, -32'sd489936, 32'sd250259, 32'sd1241609, -32'sd32241, 32'sd1034587, 32'sd3856358, 32'sd2253678, 32'sd1721771, -32'sd107335, -32'sd42577, -32'sd129550, -32'sd73779, -32'sd357159, 32'sd1485877, -32'sd249272, 32'sd167991, 32'sd940100, -32'sd1593939, 32'sd216599, -32'sd1195176, 32'sd779714, -32'sd75613, 32'sd1498758, 32'sd275116, 32'sd24190, 32'sd2192117, 32'sd1510802, 32'sd29710, 32'sd1623336, -32'sd723710, -32'sd1464740, -32'sd1157705, -32'sd1098844, 32'sd792822, 32'sd332889, 32'sd1530904, -32'sd1304544, 32'sd1515263, -32'sd1296533, 32'sd833210, 32'sd1168672, 32'sd37908, -32'sd342666, 32'sd1434969, -32'sd665524, 32'sd412008, 32'sd933212, 32'sd308323, 32'sd1037940, -32'sd100837, 32'sd1935262, 32'sd2199117, 32'sd9490, 32'sd1048319, 32'sd1445513, 32'sd1716844, 32'sd1145765, -32'sd1071926, -32'sd2477259, -32'sd500755, -32'sd1848555, -32'sd760828, -32'sd957317, -32'sd223195, 32'sd204632, 32'sd723813, -32'sd667282, -32'sd805841, -32'sd52595, -32'sd387658, 32'sd227152, 32'sd61476, -32'sd1215607, -32'sd1994061, -32'sd2354715, 32'sd1028194, 32'sd218142, -32'sd15406, 32'sd1168875, 32'sd2062732, 32'sd90753, -32'sd1006842, 32'sd1093686, -32'sd60574, -32'sd637546, -32'sd2382611, -32'sd1080398, -32'sd137408, -32'sd2867309, -32'sd2663684, -32'sd338945, -32'sd1562047, -32'sd2710713, -32'sd1963660, -32'sd850247, -32'sd836191, -32'sd567250, 32'sd493574, -32'sd551988, -32'sd619390, -32'sd712018, 32'sd883651, -32'sd103177, -32'sd1636441, -32'sd163980, 32'sd313691, -32'sd312622, -32'sd1420033, -32'sd3268687, -32'sd2297113, -32'sd1399289, -32'sd298920, -32'sd2481483, -32'sd3213304, -32'sd1139605, -32'sd18649, -32'sd2232186, -32'sd3446607, -32'sd2714182, -32'sd2093490, 32'sd757740, 32'sd1769151, 32'sd131349, 32'sd2332585, -32'sd885098, 32'sd1259350, 32'sd779512, 32'sd1119049, 32'sd683886, -32'sd441953, -32'sd1568548, 32'sd1847, 32'sd70781, 32'sd285469, 32'sd1306969, -32'sd2196229, -32'sd2076034, -32'sd338001, -32'sd1277037, -32'sd342329, -32'sd3511550, -32'sd608724, 32'sd51617, 32'sd589358, -32'sd854563, 32'sd542499, -32'sd1090237, -32'sd3566847, 32'sd946979, -32'sd244064, 32'sd1366228, 32'sd2298079, -32'sd1081163, -32'sd189810, 32'sd203075, 32'sd686105, 32'sd100728, -32'sd1391914, 32'sd116019, -32'sd340833, 32'sd1477073, 32'sd2105497, -32'sd1339906, -32'sd2129105, -32'sd1934179, -32'sd2339156, -32'sd72936, 32'sd194352, -32'sd2660128, -32'sd2851962, -32'sd1283638, -32'sd1264539, 32'sd690297, -32'sd1123576, -32'sd789780, -32'sd2729207, -32'sd1352210, -32'sd180608, 32'sd186555, -32'sd289684, 32'sd1018358, 32'sd1343638, 32'sd1045505, 32'sd50899, 32'sd616515, 32'sd178637, -32'sd164476, 32'sd1470611, 32'sd2569565, 32'sd259469, -32'sd626472, -32'sd2349905, -32'sd2514791, -32'sd2140262, -32'sd473891, 32'sd1562478, -32'sd370404, -32'sd2563334, -32'sd3328768, -32'sd1295571, -32'sd2414317, 32'sd293219, -32'sd704801, 32'sd63964, 32'sd1528122, -32'sd282586, -32'sd136571, -32'sd206124, -32'sd431279, 32'sd426026, -32'sd496206, 32'sd2732450, 32'sd759665, -32'sd1662740, 32'sd720057, 32'sd174974, 32'sd530473, -32'sd1982081, -32'sd1394300, -32'sd994406, -32'sd2795896, -32'sd191928, -32'sd142594, -32'sd1255804, -32'sd1517896, -32'sd2328615, -32'sd3198231, -32'sd2535710, -32'sd3317422, -32'sd825062, 32'sd1521927, -32'sd732679, 32'sd384765, 32'sd652984, 32'sd97858, -32'sd1978344, 32'sd791388, 32'sd879382, 32'sd962412, 32'sd51458, -32'sd1465989, -32'sd2790484, -32'sd2700353, -32'sd2669928, -32'sd2934623, -32'sd3164990, -32'sd2314403, -32'sd2250245, -32'sd1780064, -32'sd530545, 32'sd196538, 32'sd1740, -32'sd961871, -32'sd1400340, -32'sd1102450, -32'sd2601527, -32'sd1892868, -32'sd1728371, 32'sd407277, 32'sd1789851, 32'sd1270000, 32'sd687529, -32'sd1105250, 32'sd1556229, 32'sd1339347, 32'sd0, 32'sd1241041, 32'sd813960, -32'sd201007, -32'sd1096726, -32'sd347765, -32'sd451315, -32'sd1037366, -32'sd2241253, -32'sd1899311, -32'sd2994907, -32'sd4272279, -32'sd3213243, -32'sd1896065, -32'sd496372, -32'sd670687, -32'sd1120524, -32'sd996741, -32'sd2439111, -32'sd2183672, 32'sd712535, 32'sd1641678, 32'sd1780432, 32'sd880753, 32'sd229921, -32'sd724231, 32'sd328798, -32'sd303103, 32'sd460830, 32'sd385051, 32'sd2093738, 32'sd1457072, -32'sd307956, -32'sd1633126, -32'sd1260530, -32'sd1963643, -32'sd1987977, -32'sd3312111, -32'sd2110169, -32'sd2516250, -32'sd2950097, -32'sd1887599, -32'sd1290366, -32'sd3307458, -32'sd210069, -32'sd879175, -32'sd1571438, -32'sd154017, 32'sd593456, 32'sd2212943, 32'sd1709659, 32'sd1798129, 32'sd1296435, 32'sd409101, -32'sd2229882, 32'sd1369880, 32'sd1160238, -32'sd1102127, 32'sd1785422, 32'sd1926390, 32'sd302936, -32'sd9322, 32'sd1204583, 32'sd74823, -32'sd1829611, -32'sd2839374, -32'sd4234229, -32'sd2081328, -32'sd2349486, -32'sd521279, -32'sd2391499, -32'sd2168516, -32'sd9012, -32'sd849762, 32'sd869783, 32'sd714710, 32'sd828225, 32'sd32763, 32'sd1872390, -32'sd326663, 32'sd97774, 32'sd931476, -32'sd764723, 32'sd445692, 32'sd0, -32'sd762030, -32'sd376097, 32'sd1155957, 32'sd1381989, 32'sd1520723, 32'sd1498685, 32'sd80669, 32'sd839149, -32'sd366995, 32'sd46138, 32'sd979029, 32'sd442707, 32'sd1216827, 32'sd54290, -32'sd512111, 32'sd1849245, 32'sd568146, -32'sd205291, 32'sd2679320, -32'sd168658, -32'sd146922, 32'sd451258, -32'sd352097, 32'sd837505, -32'sd618164, -32'sd446835, 32'sd1025161, 32'sd1555194, -32'sd111404, 32'sd259134, 32'sd586463, 32'sd2683408, 32'sd2358887, 32'sd778145, 32'sd2142435, 32'sd2611112, 32'sd2465999, 32'sd1024595, 32'sd1805770, 32'sd2313753, 32'sd2174969, 32'sd3894678, 32'sd1613476, -32'sd1631693, -32'sd273661, 32'sd1315008, -32'sd849414, -32'sd228928, 32'sd93853, 32'sd334302, -32'sd591419, 32'sd30054, 32'sd1812656, -32'sd1551927, 32'sd929635, 32'sd888797, 32'sd946534, 32'sd1166115, 32'sd1528065, 32'sd1150583, 32'sd111377, 32'sd222990, -32'sd327657, 32'sd1564515, 32'sd303619, 32'sd1223472, 32'sd2492356, 32'sd831410, 32'sd896180, 32'sd1961199, 32'sd2222755, 32'sd386767, -32'sd786051, -32'sd14966, 32'sd131030, 32'sd1775090, -32'sd525829, -32'sd229265, 32'sd1334193, -32'sd264520, 32'sd413418, 32'sd1014732, 32'sd835200, 32'sd0, 32'sd1975430, -32'sd22095, -32'sd575665, 32'sd622832, 32'sd3160648, 32'sd866662, 32'sd1225236, -32'sd477707, -32'sd1065016, 32'sd1132708, -32'sd77356, -32'sd1067097, 32'sd678980, 32'sd1549257, 32'sd1287536, 32'sd1534971, 32'sd432089, 32'sd2150031, 32'sd496008, 32'sd1166294, 32'sd622744, 32'sd1372657, -32'sd204792, 32'sd582812, 32'sd1557949, -32'sd181932, 32'sd0, 32'sd0, 32'sd0, 32'sd798935, 32'sd369972, -32'sd990226, -32'sd958660, 32'sd852367, 32'sd1864114, 32'sd114567, 32'sd171214, -32'sd160970, 32'sd474284, 32'sd94585, -32'sd719078, 32'sd1808903, -32'sd7974, -32'sd767125, 32'sd1727773, 32'sd2854588, 32'sd1116767, -32'sd1167092, -32'sd316202, 32'sd1014064, 32'sd864352, -32'sd462649, -32'sd440070, 32'sd430838, 32'sd0, 32'sd0, 32'sd0, -32'sd12582, -32'sd355947, 32'sd224919, -32'sd797537, 32'sd729524, 32'sd950125, -32'sd327800, 32'sd447452, -32'sd486361, 32'sd1958796, 32'sd628769, 32'sd3596435, 32'sd302721, -32'sd1106769, 32'sd1626108, 32'sd972207, 32'sd1017668, 32'sd1243203, 32'sd200441, 32'sd409760, 32'sd1390212, 32'sd747277, 32'sd91523, 32'sd1183405, 32'sd1403599, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1881454, 32'sd816206, -32'sd644856, 32'sd527131, -32'sd423653, 32'sd351113, 32'sd159837, 32'sd308892, 32'sd560876, 32'sd1258989, 32'sd1568239, 32'sd336755, 32'sd1475532, 32'sd737642, -32'sd13887, -32'sd1138234, -32'sd1741926, 32'sd206982, -32'sd702510, 32'sd199298, -32'sd980159, 32'sd1439866, 32'sd1312027, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1999995, 32'sd219275, 32'sd366421, 32'sd1498398, 32'sd522758, 32'sd737513, 32'sd1631359, 32'sd785845, -32'sd25316, 32'sd1328998, 32'sd1189811, 32'sd1832291, 32'sd1800972, 32'sd1092011, 32'sd810415, -32'sd730196, 32'sd1144436, 32'sd138525, -32'sd1771918, 32'sd2225077, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1330607, 32'sd614843, 32'sd1650191, 32'sd383560, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd540438, 32'sd5148, -32'sd641260, 32'sd1054989, -32'sd1684194, 32'sd874825, 32'sd1425474, -32'sd287632, -32'sd17978, 32'sd2640164, 32'sd1698799, 32'sd343805, 32'sd1338751, 32'sd428641, -32'sd365881, -32'sd771448, -32'sd783251, -32'sd742250, 32'sd1109318, -32'sd328673, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd520682, -32'sd268541, -32'sd515893, 32'sd1295888, -32'sd1016196, -32'sd24915, -32'sd220901, 32'sd1439407, 32'sd787251, 32'sd1323576, 32'sd44605, -32'sd516656, 32'sd458392, -32'sd356428, -32'sd1857565, 32'sd1906540, -32'sd344481, -32'sd2014842, 32'sd415390, 32'sd172715, 32'sd803124, 32'sd379900, 32'sd209679, -32'sd745720, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd999718, -32'sd429217, 32'sd872488, 32'sd126137, 32'sd1979220, 32'sd1740716, 32'sd950525, -32'sd731371, 32'sd1662363, 32'sd652542, 32'sd294436, 32'sd737670, -32'sd135443, -32'sd77436, -32'sd1271332, -32'sd681685, -32'sd391234, -32'sd358694, 32'sd399556, -32'sd577459, 32'sd1588019, 32'sd825733, -32'sd735666, 32'sd572246, 32'sd1141997, 32'sd0, 32'sd0, 32'sd1193941, 32'sd1145094, 32'sd202556, 32'sd256344, 32'sd974499, -32'sd1297133, 32'sd181810, 32'sd819635, -32'sd1017881, 32'sd3049131, 32'sd1298980, 32'sd1047688, -32'sd631170, 32'sd1559638, -32'sd1654109, 32'sd135363, 32'sd1751367, 32'sd664194, 32'sd1204358, 32'sd43488, 32'sd634510, 32'sd306121, 32'sd159941, 32'sd1758903, 32'sd332104, 32'sd889344, -32'sd52170, 32'sd0, -32'sd115674, 32'sd1449533, 32'sd1744257, 32'sd406963, 32'sd495551, -32'sd1249761, -32'sd321711, 32'sd807402, -32'sd1024166, -32'sd200550, 32'sd739992, 32'sd1818425, 32'sd3554096, 32'sd2546557, -32'sd31912, 32'sd1192926, -32'sd618554, 32'sd84692, 32'sd28531, 32'sd379645, -32'sd1074794, -32'sd1352104, -32'sd2062543, 32'sd754429, 32'sd1624111, 32'sd1396306, 32'sd248895, 32'sd0, 32'sd120201, -32'sd4491, -32'sd1435956, -32'sd1748878, -32'sd992581, 32'sd408627, 32'sd1066645, 32'sd1540485, 32'sd636342, 32'sd578857, 32'sd1076067, 32'sd3002408, 32'sd3987754, 32'sd2470080, 32'sd1948520, -32'sd647933, -32'sd1217392, -32'sd1671307, -32'sd1448031, -32'sd767346, -32'sd415728, -32'sd1149949, 32'sd679997, -32'sd2074998, -32'sd914975, -32'sd667175, -32'sd281267, 32'sd410056, -32'sd621457, 32'sd1000051, -32'sd936315, -32'sd11160, -32'sd1377484, -32'sd469077, 32'sd133001, 32'sd2044225, 32'sd404871, 32'sd888605, 32'sd2297179, 32'sd1327604, 32'sd1489245, 32'sd716649, 32'sd769547, -32'sd1254507, 32'sd453036, -32'sd1241059, -32'sd725732, -32'sd497161, 32'sd228917, 32'sd23303, 32'sd714760, -32'sd183961, -32'sd709444, -32'sd1488629, -32'sd443761, -32'sd15178, -32'sd273686, 32'sd1285700, 32'sd1996001, 32'sd1766377, 32'sd1508271, 32'sd47121, 32'sd436890, 32'sd1723462, 32'sd491671, 32'sd3051999, 32'sd2153067, 32'sd2060800, 32'sd1080820, -32'sd803963, -32'sd610554, 32'sd774103, 32'sd264, -32'sd638510, -32'sd1519418, -32'sd264769, -32'sd203486, -32'sd820735, -32'sd671675, -32'sd2468422, 32'sd307778, -32'sd382765, 32'sd459613, -32'sd766403, 32'sd382014, 32'sd224150, 32'sd849684, 32'sd148981, 32'sd775911, -32'sd1165, 32'sd859776, -32'sd577893, 32'sd1412464, 32'sd597162, -32'sd1943490, -32'sd2238467, -32'sd777955, 32'sd1010729, -32'sd600613, 32'sd352406, 32'sd766051, 32'sd169585, 32'sd390831, 32'sd1923156, -32'sd395579, 32'sd139845, -32'sd456392, -32'sd2702005, -32'sd1496420, 32'sd811240, 32'sd255761, 32'sd516443, -32'sd1002151, -32'sd595441, 32'sd2898441, 32'sd867278, 32'sd135641, 32'sd1578795, -32'sd1731313, -32'sd271645, -32'sd317674, -32'sd1626064, -32'sd2985847, -32'sd3647042, -32'sd2900123, 32'sd170158, 32'sd632248, 32'sd2656496, 32'sd1967044, 32'sd1188684, -32'sd177926, 32'sd1313971, -32'sd1011060, 32'sd465919, -32'sd646642, -32'sd1984894, -32'sd131729, 32'sd501334, -32'sd1198563, -32'sd14831, 32'sd202354, 32'sd1167452, 32'sd1745400, 32'sd22547, -32'sd131274, -32'sd377294, -32'sd1471652, -32'sd1300424, -32'sd305520, -32'sd545452, 32'sd1005985, -32'sd215477, 32'sd588819, 32'sd805988, -32'sd813409, 32'sd1717310, 32'sd1890686, 32'sd856230, 32'sd64497, 32'sd131043, 32'sd390487, 32'sd939492, -32'sd2341383, -32'sd863500, 32'sd178083, 32'sd1145271, 32'sd637328, 32'sd364260, -32'sd770248, -32'sd964166, -32'sd227130, 32'sd1247413, -32'sd74137, 32'sd249691, -32'sd1244757, -32'sd1321219, -32'sd472720, -32'sd3456033, 32'sd485534, 32'sd584154, -32'sd802867, 32'sd159750, 32'sd1519561, -32'sd675246, 32'sd753904, -32'sd1463602, 32'sd2041904, -32'sd779678, -32'sd302863, -32'sd2211604, -32'sd2408402, -32'sd790266, 32'sd1098397, -32'sd874314, -32'sd1375534, 32'sd362082, 32'sd683885, 32'sd2207429, -32'sd1852846, -32'sd1701390, 32'sd767742, 32'sd48288, -32'sd967857, -32'sd1287769, -32'sd571419, -32'sd1038611, 32'sd271772, -32'sd1209615, 32'sd477975, 32'sd2074561, 32'sd1602349, -32'sd882427, -32'sd1831675, -32'sd1296525, -32'sd1667866, -32'sd791605, -32'sd1645460, -32'sd2007619, -32'sd924562, -32'sd1149053, 32'sd922375, -32'sd2456773, -32'sd110644, 32'sd40777, 32'sd425451, 32'sd1169992, 32'sd705377, -32'sd2128419, 32'sd49229, -32'sd1697499, -32'sd777185, -32'sd2181949, -32'sd2366982, -32'sd1942843, 32'sd845465, 32'sd185094, 32'sd1323588, 32'sd4078753, 32'sd2369060, -32'sd854302, -32'sd2199331, -32'sd2205577, -32'sd2025914, -32'sd1271630, -32'sd384633, -32'sd3026096, -32'sd1030918, -32'sd2494913, 32'sd130918, -32'sd214019, 32'sd726789, -32'sd457863, 32'sd1374760, 32'sd208775, 32'sd179731, -32'sd2154559, 32'sd733026, 32'sd473299, -32'sd627882, -32'sd753838, -32'sd2857209, -32'sd2934266, 32'sd1928328, 32'sd2862214, 32'sd3524338, 32'sd4614487, 32'sd2482367, -32'sd241971, -32'sd126248, -32'sd643867, -32'sd2569277, -32'sd1809494, -32'sd701232, -32'sd2788314, -32'sd617144, -32'sd520742, 32'sd360110, -32'sd1656068, -32'sd661127, -32'sd404559, -32'sd260981, 32'sd1035490, 32'sd462220, -32'sd1253489, -32'sd1022577, 32'sd186929, -32'sd203449, -32'sd488092, 32'sd404948, 32'sd151792, 32'sd967754, 32'sd410340, 32'sd1991965, 32'sd3081970, 32'sd183867, 32'sd941633, 32'sd1463107, 32'sd306160, -32'sd180782, -32'sd83593, -32'sd87507, -32'sd1714180, 32'sd847449, 32'sd299352, 32'sd816147, 32'sd508163, 32'sd650123, 32'sd0, -32'sd559784, 32'sd87364, -32'sd196829, -32'sd939595, -32'sd2244896, 32'sd226617, -32'sd2756945, -32'sd2082991, 32'sd192804, -32'sd644211, 32'sd161514, -32'sd80934, 32'sd2134459, 32'sd1317501, 32'sd848112, -32'sd98620, 32'sd1027555, -32'sd450491, -32'sd46136, 32'sd1328463, 32'sd686550, 32'sd384792, 32'sd371320, 32'sd2025734, 32'sd1595576, -32'sd481017, 32'sd837814, -32'sd156463, -32'sd560472, 32'sd1039916, 32'sd1291002, -32'sd556501, -32'sd1733426, -32'sd1129052, -32'sd2749787, 32'sd60713, 32'sd1889675, 32'sd462811, -32'sd41487, 32'sd1231826, -32'sd1720221, -32'sd910801, 32'sd748929, 32'sd1627753, 32'sd1096610, 32'sd1725670, 32'sd1889206, 32'sd1987183, 32'sd1443650, 32'sd1305800, -32'sd296028, -32'sd526830, 32'sd2065334, 32'sd1832120, -32'sd107744, 32'sd2406, 32'sd225867, 32'sd515795, 32'sd1807798, -32'sd2603558, -32'sd2945979, -32'sd3394552, 32'sd632011, 32'sd1240093, 32'sd1616257, 32'sd1927145, -32'sd1241850, -32'sd1966690, -32'sd1588468, -32'sd1235195, -32'sd124913, -32'sd528467, -32'sd621885, 32'sd1283815, 32'sd178146, 32'sd1790480, -32'sd503968, 32'sd778585, -32'sd979821, 32'sd544756, -32'sd530079, 32'sd1159470, -32'sd1286922, 32'sd0, 32'sd107504, -32'sd689560, -32'sd878299, -32'sd1383975, -32'sd2103634, -32'sd2251875, 32'sd1105246, 32'sd2332682, 32'sd2515407, 32'sd2507699, 32'sd389025, -32'sd1493094, -32'sd986751, -32'sd1412548, 32'sd1098620, -32'sd1096238, -32'sd2333607, -32'sd1100681, 32'sd926372, 32'sd1892562, -32'sd589228, -32'sd888581, 32'sd1553166, 32'sd1258574, -32'sd1243937, -32'sd1838719, -32'sd194498, -32'sd287448, 32'sd480413, 32'sd977922, 32'sd1677265, 32'sd35047, -32'sd1755277, -32'sd323621, 32'sd434550, 32'sd2127343, -32'sd531874, 32'sd103268, -32'sd897425, -32'sd781939, -32'sd169614, -32'sd60447, -32'sd910163, -32'sd1369372, -32'sd1836418, 32'sd479268, -32'sd16441, 32'sd632698, 32'sd892697, -32'sd87755, 32'sd1506417, -32'sd6198, -32'sd1962340, -32'sd2027672, 32'sd119852, -32'sd5053, 32'sd292575, -32'sd330624, 32'sd2145020, -32'sd1059965, 32'sd835445, 32'sd724808, 32'sd2104586, 32'sd1300057, 32'sd1517041, -32'sd1131897, -32'sd818009, 32'sd1662911, -32'sd88961, 32'sd245077, 32'sd2153316, 32'sd738239, -32'sd418981, 32'sd1043435, 32'sd1145659, -32'sd731704, 32'sd326018, 32'sd459645, 32'sd1822984, 32'sd936198, -32'sd66656, -32'sd1811061, -32'sd589348, 32'sd0, 32'sd605069, 32'sd1303824, -32'sd681753, 32'sd338189, 32'sd734846, 32'sd838059, 32'sd2063907, 32'sd1163106, 32'sd2258189, -32'sd572414, 32'sd794034, 32'sd1227101, -32'sd832397, 32'sd629180, 32'sd436617, 32'sd320738, 32'sd1924070, 32'sd1432189, 32'sd905342, 32'sd1662812, -32'sd1331774, 32'sd1305596, 32'sd1318397, -32'sd649748, 32'sd554552, -32'sd1381981, 32'sd0, 32'sd0, 32'sd0, 32'sd1142897, 32'sd965061, -32'sd150187, -32'sd360602, 32'sd1599191, 32'sd608684, 32'sd1104462, -32'sd67369, -32'sd1181724, 32'sd1031864, 32'sd1249558, -32'sd731209, -32'sd523594, -32'sd49092, -32'sd174568, -32'sd310189, 32'sd111718, -32'sd1445480, -32'sd456308, -32'sd774952, 32'sd1335723, -32'sd407730, 32'sd168606, 32'sd1206289, -32'sd751723, 32'sd0, 32'sd0, 32'sd0, -32'sd194538, 32'sd369336, 32'sd1149709, 32'sd396029, 32'sd534062, 32'sd1248414, -32'sd988223, -32'sd1733332, -32'sd468909, -32'sd1255690, -32'sd620092, 32'sd489007, 32'sd945813, 32'sd2250558, 32'sd1984989, 32'sd2284753, 32'sd728056, -32'sd1465237, 32'sd3299, -32'sd534068, -32'sd558584, -32'sd654638, -32'sd1087020, 32'sd1001202, 32'sd1000008, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd464242, 32'sd600615, -32'sd198411, -32'sd54723, -32'sd771508, 32'sd1727803, 32'sd1195645, -32'sd770783, -32'sd154308, 32'sd1483466, -32'sd231554, -32'sd517189, -32'sd238750, 32'sd268720, 32'sd276236, 32'sd1328436, 32'sd566559, -32'sd532042, -32'sd284053, 32'sd1057483, -32'sd1055372, 32'sd240882, -32'sd535551, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd56200, 32'sd220662, 32'sd562855, -32'sd31385, 32'sd550251, -32'sd660700, -32'sd34668, 32'sd231202, -32'sd153225, -32'sd655408, -32'sd1026019, -32'sd373108, 32'sd568134, 32'sd1443153, -32'sd322818, 32'sd3887, 32'sd284673, -32'sd2133888, -32'sd370894, -32'sd623841, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1305441, -32'sd108464, -32'sd816978, -32'sd35905, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1586074, 32'sd123843, -32'sd404729, 32'sd869289, 32'sd607029, -32'sd514957, -32'sd2113954, -32'sd2089937, -32'sd698651, -32'sd808345, 32'sd863411, -32'sd1504011, -32'sd2617131, -32'sd160453, -32'sd1928315, 32'sd697286, -32'sd52121, 32'sd1042072, 32'sd261259, -32'sd485470, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd432097, -32'sd1450135, -32'sd88319, -32'sd606038, -32'sd211631, 32'sd596692, 32'sd914077, 32'sd426968, -32'sd1802222, 32'sd1328183, 32'sd1245225, 32'sd1746353, 32'sd2727860, 32'sd1161413, -32'sd901080, -32'sd463914, 32'sd505150, -32'sd2368826, -32'sd301246, -32'sd411110, 32'sd786007, 32'sd502093, 32'sd428141, 32'sd257331, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd726224, 32'sd316876, 32'sd290812, -32'sd176126, -32'sd27397, 32'sd1041711, -32'sd478563, -32'sd1810290, -32'sd1051653, 32'sd1389692, -32'sd72151, 32'sd1618713, 32'sd3025495, 32'sd2315764, 32'sd3087394, 32'sd84670, 32'sd596698, -32'sd195783, 32'sd1363125, 32'sd1723151, 32'sd54998, 32'sd660471, -32'sd738914, -32'sd1826063, 32'sd571481, 32'sd0, 32'sd0, -32'sd185263, 32'sd32125, 32'sd122924, 32'sd32523, 32'sd557601, 32'sd659091, 32'sd792484, -32'sd1378499, 32'sd531100, 32'sd1332710, -32'sd1210450, 32'sd602705, -32'sd987308, 32'sd616653, 32'sd2352198, -32'sd407253, 32'sd419648, 32'sd551670, 32'sd56731, 32'sd500242, 32'sd2922330, -32'sd1199922, 32'sd1757310, 32'sd2124949, -32'sd329974, -32'sd3280975, 32'sd242286, 32'sd0, 32'sd254226, -32'sd6476, 32'sd1087932, 32'sd1066745, -32'sd133044, 32'sd2201693, -32'sd273519, -32'sd2684308, -32'sd917036, -32'sd884140, -32'sd1491415, 32'sd1068805, 32'sd1732218, -32'sd124790, -32'sd1153398, -32'sd1666339, 32'sd1383482, 32'sd1339789, 32'sd615978, 32'sd245981, 32'sd1279283, -32'sd881461, 32'sd1403782, 32'sd1578595, -32'sd1577045, -32'sd1528168, -32'sd523760, 32'sd0, 32'sd872387, 32'sd889566, -32'sd82931, 32'sd792650, -32'sd1222525, -32'sd641915, -32'sd446470, 32'sd2387, -32'sd917652, -32'sd1857745, 32'sd768646, -32'sd676027, -32'sd935424, -32'sd987731, -32'sd1089258, -32'sd582759, 32'sd1511315, 32'sd111886, -32'sd820243, -32'sd250464, -32'sd563271, 32'sd1812269, 32'sd1281356, 32'sd1356371, 32'sd1145095, -32'sd572204, -32'sd211022, -32'sd539674, 32'sd561866, 32'sd65062, -32'sd972876, -32'sd976633, -32'sd2285148, -32'sd217877, -32'sd1622809, -32'sd880947, -32'sd2055952, -32'sd137410, 32'sd1353200, 32'sd484891, -32'sd1289756, 32'sd290965, 32'sd836111, 32'sd1120076, 32'sd1711881, -32'sd982944, -32'sd2452682, -32'sd392685, -32'sd970539, 32'sd2307491, -32'sd587046, 32'sd2417758, 32'sd2061672, -32'sd1427601, -32'sd1154739, -32'sd540576, 32'sd765768, -32'sd319795, -32'sd2870098, -32'sd1874156, -32'sd2028889, 32'sd608571, -32'sd963806, -32'sd702007, -32'sd24288, -32'sd1107300, -32'sd2063559, -32'sd401249, 32'sd529985, 32'sd1792872, -32'sd453336, 32'sd1221498, -32'sd453157, -32'sd1318209, -32'sd1518275, -32'sd2673963, -32'sd677825, -32'sd1724804, -32'sd1022500, 32'sd446120, 32'sd1737307, -32'sd28818, 32'sd356848, -32'sd192265, 32'sd874921, 32'sd796475, -32'sd2004137, -32'sd211809, 32'sd289618, 32'sd383504, 32'sd77478, -32'sd1898988, -32'sd1917271, -32'sd3194652, -32'sd1066051, 32'sd1499094, 32'sd543246, -32'sd664717, -32'sd1963726, 32'sd771028, 32'sd1088578, -32'sd865170, 32'sd367636, -32'sd1086722, 32'sd1302850, -32'sd2771918, -32'sd1405913, -32'sd1486178, 32'sd641140, -32'sd1501455, -32'sd1088648, -32'sd459175, 32'sd812818, -32'sd926574, 32'sd103713, 32'sd1551851, 32'sd2541643, 32'sd742645, -32'sd360503, -32'sd1246725, 32'sd351889, -32'sd1065169, -32'sd966542, -32'sd1389790, -32'sd2344450, -32'sd1563105, -32'sd3050854, -32'sd1487533, -32'sd840237, -32'sd485492, -32'sd928682, -32'sd1639315, -32'sd1332696, -32'sd2162635, -32'sd807528, -32'sd8552, -32'sd217882, -32'sd713514, -32'sd127769, -32'sd779131, -32'sd21098, 32'sd950917, 32'sd1227190, -32'sd555734, -32'sd366221, 32'sd1926905, 32'sd1396503, 32'sd1200667, -32'sd51254, -32'sd278868, -32'sd1111492, -32'sd3286147, -32'sd4418675, -32'sd2960018, -32'sd2400721, -32'sd1132346, -32'sd1340960, -32'sd567451, -32'sd138608, 32'sd1107805, -32'sd322535, -32'sd3058216, -32'sd2111480, -32'sd2730032, -32'sd1673374, -32'sd1131293, -32'sd794086, 32'sd55192, -32'sd726355, 32'sd312297, -32'sd533503, -32'sd726502, 32'sd665115, 32'sd1477726, -32'sd649152, 32'sd990059, 32'sd329685, 32'sd2296550, -32'sd838811, -32'sd2651539, -32'sd2150725, -32'sd1829889, -32'sd1803748, -32'sd585531, -32'sd1300827, 32'sd637610, 32'sd695720, -32'sd1743445, -32'sd2195510, -32'sd584334, 32'sd292548, -32'sd165951, 32'sd1135573, 32'sd196019, -32'sd1016883, 32'sd152194, 32'sd564056, -32'sd986869, 32'sd1345346, -32'sd397080, -32'sd1178667, 32'sd797596, -32'sd347599, 32'sd79834, 32'sd2470915, 32'sd4310714, 32'sd1188871, -32'sd322, -32'sd1315080, -32'sd936076, -32'sd1169652, 32'sd1946452, 32'sd122498, -32'sd1563817, 32'sd391528, -32'sd563920, -32'sd1219531, -32'sd954297, -32'sd1994120, 32'sd164920, -32'sd1285036, 32'sd538540, -32'sd32925, 32'sd100720, 32'sd146061, 32'sd301804, 32'sd1330608, -32'sd997572, 32'sd19830, 32'sd1423514, 32'sd359858, 32'sd844715, 32'sd306291, 32'sd1270246, 32'sd1613705, 32'sd2027225, 32'sd2199490, 32'sd506021, 32'sd617465, 32'sd1687610, 32'sd1427041, -32'sd1164645, -32'sd1025157, -32'sd2233887, -32'sd1224626, -32'sd946780, -32'sd456447, -32'sd656491, 32'sd132215, 32'sd935395, -32'sd601127, -32'sd817833, -32'sd380768, -32'sd1118738, 32'sd1347876, 32'sd35828, 32'sd96841, 32'sd1133605, 32'sd1385916, 32'sd1548242, 32'sd885307, 32'sd960573, 32'sd817152, 32'sd1980533, 32'sd2159775, 32'sd1583528, 32'sd2528358, 32'sd3492178, -32'sd180777, -32'sd1749740, -32'sd1047164, -32'sd2346643, -32'sd856249, 32'sd1005408, 32'sd879225, 32'sd753805, -32'sd634955, 32'sd205255, -32'sd176228, 32'sd838005, 32'sd591679, -32'sd94754, 32'sd202707, 32'sd490149, 32'sd803509, 32'sd2542918, 32'sd2861892, 32'sd2554569, 32'sd1318703, 32'sd666097, 32'sd1945089, 32'sd3897747, 32'sd2689396, -32'sd291053, 32'sd1449497, 32'sd1446625, 32'sd1516094, -32'sd835191, 32'sd582212, -32'sd65164, -32'sd1183664, 32'sd348803, -32'sd343341, -32'sd463993, 32'sd51876, 32'sd842401, 32'sd144872, 32'sd0, 32'sd1096774, 32'sd192865, 32'sd1701872, -32'sd1132137, 32'sd462432, 32'sd807035, 32'sd916084, 32'sd998265, 32'sd2070539, 32'sd3620143, 32'sd1542596, 32'sd2728095, 32'sd972547, -32'sd517813, -32'sd92579, 32'sd1083796, 32'sd735345, -32'sd2059816, -32'sd243524, -32'sd779381, 32'sd493983, -32'sd1350582, -32'sd666480, 32'sd923189, -32'sd268179, -32'sd637901, -32'sd798157, -32'sd43723, -32'sd1698767, -32'sd1478381, 32'sd1175056, -32'sd812952, -32'sd2852861, -32'sd519429, 32'sd1714328, 32'sd3170487, 32'sd2926321, 32'sd179207, 32'sd2166123, 32'sd2439576, 32'sd2140144, -32'sd901626, 32'sd1223733, 32'sd408300, 32'sd281273, -32'sd858073, -32'sd1316330, -32'sd1007217, -32'sd568047, -32'sd293798, 32'sd632406, 32'sd1817682, 32'sd1715471, -32'sd2758265, -32'sd984734, 32'sd900827, -32'sd819498, -32'sd2056873, 32'sd741095, 32'sd1588919, -32'sd356133, -32'sd2130503, -32'sd878785, -32'sd813948, -32'sd948536, -32'sd1468610, -32'sd720563, 32'sd1733882, 32'sd1486421, 32'sd410944, 32'sd84691, 32'sd720208, 32'sd2120623, -32'sd123028, -32'sd435488, -32'sd1899654, 32'sd862943, -32'sd225646, 32'sd385529, 32'sd1392036, 32'sd897702, 32'sd108113, -32'sd1202117, 32'sd0, 32'sd777359, 32'sd664398, 32'sd52814, -32'sd2798511, -32'sd2344983, -32'sd1673655, -32'sd588704, -32'sd62515, 32'sd310305, -32'sd2337793, -32'sd1379874, -32'sd987740, 32'sd1141798, 32'sd1304898, 32'sd169866, -32'sd857540, 32'sd1679436, 32'sd2182262, -32'sd873062, 32'sd907287, 32'sd476213, 32'sd996882, -32'sd1366201, 32'sd431317, -32'sd536153, -32'sd110445, 32'sd411699, -32'sd704319, 32'sd1446629, 32'sd207610, -32'sd181073, -32'sd2107883, -32'sd994054, -32'sd1315078, -32'sd1814802, -32'sd376550, 32'sd32008, -32'sd458984, -32'sd1539109, -32'sd914010, 32'sd2241961, -32'sd776134, 32'sd1148882, -32'sd171497, 32'sd2135300, 32'sd2381543, 32'sd200694, 32'sd78569, -32'sd856804, 32'sd1344592, 32'sd275968, -32'sd1820514, -32'sd1439553, -32'sd882949, 32'sd634657, 32'sd220678, -32'sd122878, 32'sd142442, 32'sd1486413, 32'sd447022, -32'sd509865, -32'sd3620757, -32'sd2664301, -32'sd2044016, 32'sd74968, 32'sd462045, 32'sd653400, -32'sd335991, -32'sd9392, -32'sd1009966, 32'sd1714194, 32'sd3120853, 32'sd706754, 32'sd2826444, 32'sd1619757, 32'sd1862390, 32'sd1454586, 32'sd461922, -32'sd2446933, -32'sd727556, -32'sd1223038, 32'sd375491, -32'sd297684, 32'sd0, 32'sd1123379, -32'sd488237, 32'sd1935911, 32'sd686584, 32'sd103916, -32'sd866178, -32'sd3678138, -32'sd605394, -32'sd683679, 32'sd922088, -32'sd241535, -32'sd1172371, -32'sd2071157, 32'sd312901, 32'sd2018773, -32'sd330778, 32'sd1203919, 32'sd1489527, 32'sd1827456, 32'sd845652, 32'sd1048043, -32'sd175687, -32'sd378044, -32'sd339338, -32'sd1510333, -32'sd387272, 32'sd0, 32'sd0, 32'sd0, -32'sd1033535, -32'sd709909, -32'sd2365218, -32'sd1599075, 32'sd419058, -32'sd146460, 32'sd1095604, -32'sd273000, -32'sd270961, 32'sd2588556, -32'sd382889, 32'sd1178113, 32'sd1605060, -32'sd433701, 32'sd501723, -32'sd1966947, -32'sd384623, 32'sd1514412, 32'sd2511528, -32'sd654754, -32'sd134452, 32'sd1089233, -32'sd1585736, 32'sd241618, 32'sd926607, 32'sd0, 32'sd0, 32'sd0, -32'sd506981, -32'sd547782, -32'sd891282, 32'sd1101085, -32'sd448120, -32'sd18200, -32'sd1283919, 32'sd346415, -32'sd928629, 32'sd811702, 32'sd2718148, 32'sd1756927, -32'sd1634356, -32'sd1605007, -32'sd2088085, -32'sd1972154, 32'sd651894, 32'sd1866615, 32'sd1194173, -32'sd1334537, -32'sd589579, -32'sd1133085, -32'sd261756, 32'sd1330254, 32'sd328298, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd337148, 32'sd734321, 32'sd670229, 32'sd1543226, 32'sd593268, 32'sd51909, -32'sd887548, -32'sd2002504, 32'sd509271, 32'sd966492, 32'sd1559745, 32'sd967609, 32'sd481900, 32'sd194653, -32'sd1823836, -32'sd179937, -32'sd524495, -32'sd872431, 32'sd792690, 32'sd779774, -32'sd330790, 32'sd1359825, -32'sd528826, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd674588, -32'sd745914, -32'sd613933, 32'sd893659, 32'sd1178131, -32'sd108923, 32'sd731996, 32'sd813422, 32'sd1549063, 32'sd131796, 32'sd1035693, 32'sd780927, 32'sd95765, -32'sd252758, -32'sd1131556, 32'sd480240, 32'sd866243, 32'sd682332, 32'sd563788, 32'sd9488, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2232608, 32'sd1003227, 32'sd1682360, 32'sd621706, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd454683, 32'sd457775, -32'sd75039, 32'sd2510073, 32'sd2265961, 32'sd1167570, 32'sd217284, 32'sd709827, 32'sd1887399, 32'sd844331, -32'sd90217, 32'sd1073469, 32'sd801412, 32'sd17905, -32'sd1388921, 32'sd896997, 32'sd839766, 32'sd1644305, 32'sd407084, 32'sd316994, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd885969, 32'sd1528275, 32'sd6504, -32'sd77849, 32'sd1004164, -32'sd453705, 32'sd1829744, 32'sd2210513, 32'sd328875, 32'sd388102, 32'sd1586504, 32'sd1378158, 32'sd722225, 32'sd1490139, 32'sd1003366, 32'sd1715069, 32'sd450729, 32'sd548575, 32'sd1407760, 32'sd1295451, 32'sd1342245, 32'sd1189644, -32'sd179938, 32'sd1393787, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1251337, 32'sd1666660, 32'sd611801, 32'sd442925, -32'sd5198, 32'sd1814736, 32'sd1367687, 32'sd2654373, 32'sd26791, 32'sd1319170, -32'sd1573889, 32'sd506459, 32'sd504135, -32'sd291373, 32'sd146836, -32'sd1269612, -32'sd1630330, -32'sd1703854, -32'sd2316062, 32'sd469668, -32'sd951343, 32'sd475664, 32'sd264609, 32'sd128810, 32'sd1675206, 32'sd0, 32'sd0, 32'sd787860, 32'sd1072274, -32'sd316679, 32'sd805185, 32'sd1335893, -32'sd951277, 32'sd337492, 32'sd780238, -32'sd555379, 32'sd1061735, -32'sd1205520, 32'sd311884, -32'sd1346042, -32'sd204945, 32'sd1381094, 32'sd1903913, 32'sd492036, -32'sd962814, -32'sd219088, -32'sd24045, 32'sd527804, 32'sd2642724, -32'sd519518, -32'sd1034939, -32'sd2049575, 32'sd731656, 32'sd610583, 32'sd0, 32'sd1195316, -32'sd1478271, 32'sd432496, 32'sd1363338, -32'sd34654, -32'sd251150, 32'sd287123, 32'sd400482, -32'sd761951, -32'sd2837315, -32'sd2215336, -32'sd910652, -32'sd2139390, 32'sd60120, 32'sd370369, -32'sd143477, 32'sd905516, -32'sd1694903, -32'sd519440, -32'sd224695, 32'sd787549, 32'sd1661255, 32'sd2868744, -32'sd1302217, -32'sd360413, -32'sd3334557, 32'sd49895, 32'sd0, 32'sd694101, -32'sd5059, -32'sd1163360, 32'sd614127, 32'sd1552302, 32'sd829326, 32'sd1454581, 32'sd2764399, 32'sd858572, -32'sd3977268, -32'sd2085578, -32'sd3267700, -32'sd4053867, -32'sd2581287, -32'sd396580, 32'sd815365, -32'sd389994, 32'sd576752, 32'sd360392, -32'sd415166, -32'sd229555, 32'sd143669, -32'sd616397, 32'sd632044, -32'sd809514, 32'sd351763, -32'sd1314752, 32'sd1897298, -32'sd1332161, -32'sd1713908, -32'sd156953, 32'sd1170179, 32'sd183301, 32'sd3472, 32'sd276016, 32'sd415356, -32'sd2533572, -32'sd2292581, -32'sd2622737, -32'sd1960570, -32'sd2000183, -32'sd1156331, 32'sd231944, 32'sd2171082, -32'sd233935, -32'sd2406672, 32'sd2326551, 32'sd1744710, 32'sd32701, -32'sd1551281, -32'sd731916, -32'sd260825, -32'sd430191, 32'sd147565, 32'sd696570, -32'sd216364, -32'sd1029042, -32'sd235121, -32'sd984135, 32'sd892525, -32'sd334823, 32'sd2175764, 32'sd95661, -32'sd62292, -32'sd1830438, -32'sd864455, -32'sd592238, -32'sd589126, -32'sd1799516, 32'sd2161107, 32'sd233094, 32'sd1034163, -32'sd1465816, -32'sd1147233, 32'sd1432475, 32'sd790258, -32'sd319932, -32'sd846497, -32'sd2268400, 32'sd68963, -32'sd32219, 32'sd862736, 32'sd1075434, 32'sd716332, -32'sd67639, 32'sd27479, 32'sd133920, 32'sd349669, 32'sd344668, 32'sd1722621, 32'sd720466, -32'sd669870, 32'sd26492, 32'sd1131106, -32'sd1557989, -32'sd1743807, -32'sd2582537, 32'sd202726, 32'sd1310412, 32'sd1486595, -32'sd634546, -32'sd1424089, -32'sd727100, -32'sd917524, 32'sd1535065, -32'sd1437870, -32'sd715465, -32'sd757132, -32'sd68382, 32'sd793001, 32'sd1274678, 32'sd262284, 32'sd1429216, -32'sd1116238, -32'sd196749, -32'sd611147, 32'sd329276, -32'sd556162, 32'sd528201, -32'sd957197, 32'sd876153, 32'sd343344, -32'sd1864608, -32'sd3459711, -32'sd1478105, -32'sd23402, 32'sd1124279, -32'sd321379, -32'sd472451, -32'sd402045, -32'sd202560, -32'sd1963874, -32'sd122262, -32'sd246314, -32'sd949477, -32'sd264779, -32'sd1036854, -32'sd787612, 32'sd1316618, 32'sd3677, 32'sd151345, 32'sd748600, -32'sd223673, 32'sd388106, -32'sd1167696, 32'sd747621, -32'sd966192, 32'sd1453800, 32'sd3119807, 32'sd663757, -32'sd1627308, -32'sd2181814, -32'sd2592805, 32'sd767815, -32'sd561572, 32'sd801076, -32'sd2324355, -32'sd1711641, 32'sd704249, -32'sd2299090, -32'sd380671, -32'sd2007650, 32'sd921320, -32'sd2089569, -32'sd701262, 32'sd365209, -32'sd22523, 32'sd837102, -32'sd403315, 32'sd824337, 32'sd423383, -32'sd254215, 32'sd128672, -32'sd1156154, -32'sd45461, 32'sd1905566, 32'sd1662556, 32'sd553758, -32'sd1624934, 32'sd930062, -32'sd183529, -32'sd355225, -32'sd966156, 32'sd178957, -32'sd1117093, -32'sd126711, -32'sd813420, -32'sd1079279, -32'sd372888, -32'sd161262, -32'sd743023, -32'sd1095400, 32'sd687952, -32'sd761504, -32'sd55209, 32'sd541692, 32'sd366859, -32'sd115497, -32'sd1753047, -32'sd2135021, -32'sd350177, -32'sd1340282, 32'sd1370884, 32'sd1615480, 32'sd3478689, 32'sd2247391, -32'sd733641, 32'sd236535, -32'sd1023613, -32'sd736405, 32'sd1960761, 32'sd42176, 32'sd319375, 32'sd1051308, -32'sd746599, -32'sd1405231, -32'sd490391, 32'sd85468, -32'sd224651, -32'sd501946, -32'sd452264, -32'sd374100, 32'sd1731213, 32'sd1050851, 32'sd367489, 32'sd559629, 32'sd414701, -32'sd916691, -32'sd556333, -32'sd1052998, 32'sd54421, 32'sd1750765, 32'sd963288, 32'sd1173898, -32'sd647865, -32'sd1730874, -32'sd530717, 32'sd2198376, 32'sd1352033, 32'sd2699992, 32'sd481652, 32'sd527327, 32'sd87319, -32'sd507880, -32'sd2114634, -32'sd632451, -32'sd138790, 32'sd1356245, -32'sd418575, 32'sd450954, 32'sd2662643, -32'sd1297514, 32'sd965890, -32'sd176699, 32'sd765213, 32'sd111342, 32'sd1772101, -32'sd59604, -32'sd109460, 32'sd1130919, 32'sd628317, 32'sd134830, -32'sd1123698, -32'sd1487446, 32'sd106841, 32'sd1928016, -32'sd452820, 32'sd1180996, 32'sd1283915, 32'sd133665, -32'sd1495297, 32'sd1270532, -32'sd1071297, 32'sd416019, 32'sd1220584, 32'sd1297217, -32'sd1861673, -32'sd2269684, 32'sd1333679, 32'sd455269, -32'sd1623359, -32'sd252641, -32'sd404483, -32'sd1183704, 32'sd112361, -32'sd196338, -32'sd308794, -32'sd22984, 32'sd376607, 32'sd514833, -32'sd456960, 32'sd188300, 32'sd146818, -32'sd889153, 32'sd2709384, 32'sd2183911, -32'sd254475, 32'sd554677, -32'sd124793, 32'sd784402, 32'sd1163666, 32'sd606428, -32'sd468155, 32'sd493848, 32'sd1248193, 32'sd139054, 32'sd1159889, 32'sd0, -32'sd944934, -32'sd361299, -32'sd825756, 32'sd910, 32'sd1329781, -32'sd598916, 32'sd439464, 32'sd1006578, -32'sd2040030, -32'sd370715, -32'sd1408480, -32'sd1299274, 32'sd299779, 32'sd1932207, 32'sd2961495, 32'sd2796256, 32'sd235122, -32'sd832974, -32'sd1840708, -32'sd2465482, -32'sd682229, 32'sd2536259, 32'sd241147, -32'sd1573794, -32'sd463061, -32'sd1006479, -32'sd499877, 32'sd748927, 32'sd990368, -32'sd1737000, 32'sd1710434, -32'sd504779, -32'sd103990, -32'sd1731482, -32'sd599313, 32'sd59747, 32'sd308458, -32'sd789050, -32'sd142207, 32'sd1517800, 32'sd1631525, 32'sd3103852, 32'sd1524850, -32'sd234035, 32'sd206726, -32'sd506797, -32'sd1052114, -32'sd1812625, -32'sd1573122, 32'sd745390, -32'sd1842760, -32'sd1847774, -32'sd1144455, -32'sd1339175, 32'sd728943, 32'sd1075251, -32'sd511624, -32'sd1468943, 32'sd1748019, 32'sd230062, -32'sd318537, -32'sd650286, 32'sd61671, -32'sd571673, -32'sd1291473, 32'sd481981, 32'sd1537734, 32'sd2282009, 32'sd2472199, 32'sd3084624, 32'sd1425198, 32'sd1423942, -32'sd1015170, -32'sd733675, -32'sd713867, -32'sd305502, -32'sd1528299, -32'sd483055, -32'sd794375, -32'sd2246006, 32'sd241453, -32'sd441978, 32'sd131012, 32'sd0, 32'sd131427, -32'sd1240530, 32'sd1180950, 32'sd344662, -32'sd1368161, -32'sd2036934, -32'sd560840, -32'sd268605, -32'sd636477, -32'sd617891, 32'sd1731984, 32'sd1555049, 32'sd293395, 32'sd3728607, 32'sd1740344, 32'sd2960410, -32'sd33599, 32'sd197978, -32'sd679602, -32'sd1469046, -32'sd2204098, -32'sd2742639, -32'sd1376984, 32'sd522385, 32'sd1301576, -32'sd940637, -32'sd253519, 32'sd1650729, 32'sd445887, 32'sd806451, 32'sd994189, 32'sd578922, -32'sd1053592, -32'sd2360448, -32'sd1929729, -32'sd2058215, -32'sd468683, -32'sd789825, -32'sd914072, -32'sd1243470, 32'sd1336928, 32'sd1317069, -32'sd368790, -32'sd66500, 32'sd158741, 32'sd1701268, 32'sd1110125, -32'sd996961, -32'sd1145222, 32'sd449093, 32'sd950964, 32'sd558805, 32'sd1430582, -32'sd1613801, -32'sd857488, 32'sd1724464, 32'sd1527916, 32'sd294395, -32'sd615466, 32'sd515646, 32'sd411624, -32'sd807709, -32'sd1175075, -32'sd2074692, -32'sd1102890, -32'sd36432, 32'sd373258, -32'sd1307250, 32'sd1670979, 32'sd1770057, -32'sd990246, 32'sd37600, -32'sd278129, 32'sd2573312, 32'sd2302284, 32'sd1898132, 32'sd2416532, 32'sd1023517, -32'sd341444, -32'sd1492148, -32'sd455861, 32'sd669184, 32'sd1012599, 32'sd0, 32'sd1259254, 32'sd543380, 32'sd396969, -32'sd295744, -32'sd1539910, -32'sd1235235, -32'sd965655, -32'sd1170273, -32'sd524426, 32'sd588197, -32'sd903108, 32'sd1948080, 32'sd1994168, 32'sd2505433, -32'sd1234196, 32'sd1263673, 32'sd452880, 32'sd2285057, 32'sd84612, 32'sd1588532, 32'sd1442148, 32'sd903423, -32'sd1614957, -32'sd1341009, 32'sd808146, 32'sd449875, 32'sd0, 32'sd0, 32'sd0, -32'sd1152431, -32'sd851813, -32'sd1461569, -32'sd354099, -32'sd166331, 32'sd1559515, 32'sd805840, -32'sd870207, -32'sd186901, -32'sd1176075, 32'sd702753, 32'sd314176, 32'sd1597838, 32'sd1514875, -32'sd1013662, -32'sd1422573, 32'sd959480, 32'sd540737, 32'sd1481174, -32'sd393242, -32'sd1267708, -32'sd981918, -32'sd74094, 32'sd422019, 32'sd1719983, 32'sd0, 32'sd0, 32'sd0, 32'sd1057899, 32'sd1087854, -32'sd606152, 32'sd452349, -32'sd1349953, 32'sd14747, 32'sd150675, 32'sd564225, -32'sd1891370, -32'sd101433, 32'sd1819875, 32'sd1282598, 32'sd1599985, 32'sd779518, 32'sd181057, -32'sd1308968, -32'sd1149466, 32'sd7529, 32'sd403953, 32'sd1117637, 32'sd394744, 32'sd273225, 32'sd167560, 32'sd1041878, -32'sd889859, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1399262, 32'sd895540, -32'sd113662, 32'sd260370, -32'sd1138256, -32'sd991817, -32'sd1555916, 32'sd561441, 32'sd68989, -32'sd1371157, -32'sd2433313, -32'sd49827, -32'sd1224241, 32'sd383506, 32'sd455843, 32'sd1469553, 32'sd1413983, -32'sd1410614, -32'sd1492491, -32'sd2181852, 32'sd1136487, 32'sd705234, 32'sd705022, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1127690, 32'sd355393, 32'sd894101, -32'sd141151, -32'sd1010608, -32'sd90891, -32'sd40387, -32'sd602202, 32'sd320920, -32'sd467947, -32'sd1009717, 32'sd852075, -32'sd1034892, 32'sd409155, 32'sd465126, 32'sd64393, -32'sd1336208, 32'sd1119268, 32'sd858438, 32'sd28768, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1299375, 32'sd1363136, 32'sd730084, 32'sd925372, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1684350, -32'sd1280683, 32'sd628092, 32'sd879562, 32'sd550470, -32'sd68222, 32'sd12136, 32'sd809740, 32'sd584146, 32'sd365696, 32'sd818605, -32'sd912691, 32'sd1121351, 32'sd529330, 32'sd1991591, 32'sd151085, -32'sd529409, 32'sd81591, 32'sd103158, 32'sd1101868, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd590432, 32'sd468074, 32'sd754255, 32'sd713216, 32'sd861826, -32'sd1494580, 32'sd435232, 32'sd271926, 32'sd832974, 32'sd584379, -32'sd1090899, -32'sd378796, 32'sd577073, -32'sd1868839, -32'sd2960097, -32'sd672469, -32'sd452220, 32'sd77309, 32'sd119906, 32'sd1575261, 32'sd845571, -32'sd1458725, 32'sd1060901, 32'sd768856, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd58850, 32'sd405673, 32'sd605545, 32'sd687067, 32'sd1748708, 32'sd588803, -32'sd1146971, -32'sd53218, -32'sd621860, -32'sd1004228, -32'sd1918100, -32'sd2954561, -32'sd1063276, -32'sd1735640, -32'sd1576830, -32'sd1147122, -32'sd3562989, -32'sd869933, -32'sd2149235, -32'sd1545792, -32'sd339657, 32'sd281132, 32'sd1388220, 32'sd115006, -32'sd772474, 32'sd0, 32'sd0, 32'sd1084307, 32'sd541859, -32'sd383746, 32'sd353618, 32'sd524224, -32'sd112470, 32'sd1122163, 32'sd2524466, 32'sd724677, 32'sd307926, -32'sd1275512, -32'sd134814, 32'sd1031184, -32'sd2110217, -32'sd2696944, -32'sd3031350, -32'sd998844, -32'sd1296274, -32'sd1208706, -32'sd68350, -32'sd47578, 32'sd2005939, 32'sd1529315, -32'sd970726, -32'sd194321, -32'sd489869, 32'sd1694071, 32'sd0, 32'sd673461, 32'sd2099393, 32'sd478828, 32'sd533204, 32'sd2001371, 32'sd1710871, 32'sd628321, 32'sd1897031, 32'sd1825147, 32'sd851223, -32'sd941205, -32'sd2492698, -32'sd3268479, -32'sd2248138, -32'sd1461802, -32'sd792696, -32'sd256721, -32'sd1293071, -32'sd1408978, -32'sd1459919, 32'sd181560, 32'sd1181617, 32'sd1949824, -32'sd552086, -32'sd143798, -32'sd197584, -32'sd22957, 32'sd0, -32'sd388574, -32'sd653513, -32'sd33303, 32'sd990838, 32'sd50746, -32'sd2097203, -32'sd20187, 32'sd1346845, 32'sd868622, 32'sd96333, -32'sd1425885, -32'sd1124407, -32'sd3495428, -32'sd3266800, -32'sd2935477, -32'sd2189667, -32'sd1928745, -32'sd1052912, -32'sd229390, 32'sd230993, -32'sd1561646, -32'sd2210427, -32'sd1043308, -32'sd811517, -32'sd1296499, 32'sd1754772, 32'sd327590, 32'sd579740, 32'sd760181, -32'sd1080493, -32'sd2383578, -32'sd182691, 32'sd574279, -32'sd2194051, 32'sd1256157, 32'sd1343055, 32'sd2706402, -32'sd237270, -32'sd529967, -32'sd1141459, -32'sd3682745, -32'sd4360330, -32'sd2959006, 32'sd8034, -32'sd1325784, -32'sd2371081, -32'sd1902541, 32'sd656757, -32'sd2112426, -32'sd1261474, -32'sd2036259, 32'sd815995, -32'sd99435, -32'sd235895, -32'sd994915, 32'sd781793, -32'sd104032, -32'sd671354, -32'sd972798, 32'sd2173626, 32'sd435644, -32'sd120034, 32'sd1433121, 32'sd598, 32'sd1707684, 32'sd945962, 32'sd864964, -32'sd1962005, -32'sd3342810, -32'sd3004478, -32'sd1741205, -32'sd116650, 32'sd77891, -32'sd685932, -32'sd735456, -32'sd393839, -32'sd1686815, -32'sd473915, -32'sd380418, 32'sd1786933, -32'sd159595, 32'sd299701, -32'sd1505536, 32'sd1215130, 32'sd813904, 32'sd1389548, 32'sd522112, 32'sd345352, -32'sd2225920, -32'sd2173233, -32'sd493809, -32'sd252690, 32'sd642329, 32'sd1549761, 32'sd686359, -32'sd2710110, -32'sd4773644, -32'sd3624802, -32'sd1624972, 32'sd1470698, 32'sd1725782, 32'sd176861, 32'sd1106156, 32'sd352057, 32'sd1492525, -32'sd1204886, -32'sd403416, 32'sd439881, -32'sd718687, 32'sd463496, 32'sd1246547, 32'sd504161, 32'sd724470, 32'sd1980948, -32'sd689859, -32'sd1234586, -32'sd1523030, -32'sd1736736, 32'sd638917, 32'sd997354, 32'sd863313, 32'sd777056, 32'sd799344, -32'sd2842908, -32'sd3077798, -32'sd3135038, 32'sd1580190, 32'sd1581545, 32'sd1140046, 32'sd521374, 32'sd247688, -32'sd1741730, 32'sd595726, 32'sd136369, -32'sd751118, 32'sd2707125, 32'sd1161700, 32'sd1483902, -32'sd421277, 32'sd621300, 32'sd1875601, -32'sd1066168, -32'sd750089, 32'sd55855, 32'sd1181920, 32'sd275680, -32'sd12280, -32'sd725884, 32'sd220766, -32'sd565595, -32'sd329460, -32'sd1878519, -32'sd2862757, -32'sd1428440, 32'sd1669561, -32'sd337331, -32'sd1321171, -32'sd165928, 32'sd1263959, -32'sd99250, 32'sd502617, -32'sd33050, 32'sd605888, 32'sd1538091, -32'sd111743, -32'sd1139465, -32'sd4009, 32'sd1450623, 32'sd177150, 32'sd64496, -32'sd101067, 32'sd157801, -32'sd604526, -32'sd739429, -32'sd924981, -32'sd1637223, -32'sd1497203, 32'sd590664, -32'sd672416, -32'sd146853, 32'sd516751, 32'sd1972341, 32'sd2127602, 32'sd2676407, -32'sd777649, -32'sd1658240, 32'sd603115, 32'sd1871081, 32'sd1704078, 32'sd1982903, -32'sd30003, -32'sd466265, 32'sd1710730, -32'sd481311, 32'sd154245, 32'sd491425, 32'sd1902690, -32'sd828333, -32'sd467156, -32'sd181545, 32'sd574038, -32'sd1353074, 32'sd527604, 32'sd897134, -32'sd431101, 32'sd1256380, -32'sd70637, -32'sd932379, 32'sd225263, 32'sd1562945, 32'sd1338994, -32'sd211767, 32'sd1090258, 32'sd897488, 32'sd3086521, 32'sd2853745, 32'sd2554554, 32'sd2542479, 32'sd1835122, -32'sd95060, -32'sd309497, 32'sd592251, -32'sd1318690, 32'sd433294, 32'sd227485, 32'sd193988, -32'sd1772451, 32'sd1774656, 32'sd2566711, 32'sd1135431, 32'sd2493768, 32'sd1187059, 32'sd1573983, 32'sd797330, 32'sd39433, 32'sd3255145, 32'sd2736680, 32'sd1051045, -32'sd162492, 32'sd878942, 32'sd1433482, -32'sd349660, 32'sd2792404, -32'sd9721, 32'sd754068, 32'sd1188869, 32'sd851094, 32'sd2004684, 32'sd922686, -32'sd952209, 32'sd791698, -32'sd373246, -32'sd261110, 32'sd370211, 32'sd988389, -32'sd638868, 32'sd1108296, 32'sd803709, 32'sd2938016, 32'sd1916761, 32'sd1082003, 32'sd2840048, 32'sd1866068, 32'sd2001177, 32'sd3131979, 32'sd2520849, 32'sd214960, -32'sd113410, 32'sd1820672, -32'sd658118, 32'sd606115, 32'sd847678, -32'sd1320410, 32'sd1563990, -32'sd7853, 32'sd531909, 32'sd1643537, -32'sd816314, 32'sd1171799, 32'sd453633, 32'sd1947392, -32'sd630189, 32'sd164556, -32'sd1347465, 32'sd900471, 32'sd1325750, 32'sd1693787, 32'sd940171, -32'sd318898, 32'sd136208, 32'sd184717, 32'sd1280267, -32'sd621349, -32'sd619513, 32'sd3412642, 32'sd314058, 32'sd895109, 32'sd1861939, 32'sd1208383, 32'sd1683773, 32'sd431547, -32'sd686484, -32'sd1036438, -32'sd2988599, -32'sd1007683, -32'sd1116128, 32'sd697462, 32'sd0, 32'sd496921, -32'sd791666, -32'sd412149, -32'sd633612, 32'sd1598605, 32'sd571154, 32'sd242698, 32'sd1004607, -32'sd172462, 32'sd1291709, -32'sd276749, 32'sd110166, 32'sd85947, 32'sd1339578, 32'sd1288709, -32'sd35338, -32'sd218178, -32'sd91700, 32'sd405622, 32'sd1776967, 32'sd911270, -32'sd206280, -32'sd397776, -32'sd2208633, -32'sd630976, -32'sd239169, -32'sd893603, 32'sd120485, 32'sd864887, -32'sd952016, 32'sd845176, 32'sd25391, -32'sd80600, 32'sd1375174, -32'sd1135144, -32'sd646750, 32'sd1198342, 32'sd653507, 32'sd2100661, 32'sd470328, 32'sd190941, 32'sd2423421, 32'sd806227, -32'sd102711, 32'sd523485, 32'sd1594595, 32'sd1489414, 32'sd2276497, 32'sd941521, -32'sd557569, -32'sd1733871, -32'sd878683, 32'sd365019, 32'sd350762, 32'sd1519662, 32'sd457243, 32'sd601806, 32'sd535734, 32'sd1301915, 32'sd1277908, 32'sd1323486, 32'sd1798243, 32'sd1311854, 32'sd881343, 32'sd668315, 32'sd1053457, -32'sd21887, -32'sd2351307, -32'sd1376513, -32'sd813125, 32'sd411860, 32'sd917118, -32'sd923917, 32'sd835089, -32'sd1795845, -32'sd66490, 32'sd870818, -32'sd439095, -32'sd10022, -32'sd1924908, -32'sd1558284, -32'sd1030117, 32'sd472215, 32'sd0, 32'sd518719, -32'sd375655, 32'sd902301, 32'sd1256319, 32'sd421650, 32'sd2509353, 32'sd1220828, -32'sd607654, 32'sd132296, -32'sd2108112, -32'sd396096, -32'sd3373267, -32'sd3255294, -32'sd463055, -32'sd463432, 32'sd993807, -32'sd1827198, -32'sd711316, -32'sd3128151, -32'sd1468006, -32'sd241656, -32'sd364787, -32'sd1245008, -32'sd1238357, -32'sd2878603, 32'sd397587, 32'sd369584, 32'sd1412207, 32'sd1500050, 32'sd160904, 32'sd52338, 32'sd1470681, 32'sd1167423, -32'sd622861, -32'sd431707, -32'sd657833, -32'sd827552, -32'sd1497679, -32'sd3043649, -32'sd1983331, -32'sd2366681, -32'sd918568, -32'sd1017122, -32'sd314223, -32'sd1443894, -32'sd2297682, 32'sd104926, -32'sd875665, 32'sd415018, 32'sd733988, 32'sd18104, -32'sd909408, 32'sd854372, 32'sd1399632, 32'sd456415, 32'sd1250017, 32'sd2498502, 32'sd986119, 32'sd1273717, -32'sd503869, -32'sd322307, -32'sd1238325, 32'sd1417361, 32'sd571215, -32'sd193237, -32'sd1179437, -32'sd721342, -32'sd1757967, -32'sd7499, -32'sd2447491, -32'sd1980799, -32'sd1059315, -32'sd659767, -32'sd1353751, -32'sd634891, -32'sd411636, -32'sd382052, 32'sd1475205, -32'sd136332, 32'sd1663912, -32'sd950183, -32'sd161030, 32'sd113905, 32'sd0, 32'sd630385, 32'sd1174753, 32'sd530387, -32'sd284441, 32'sd137705, -32'sd303055, 32'sd1394104, 32'sd6695, -32'sd795567, -32'sd674812, -32'sd1149499, 32'sd100570, -32'sd908429, -32'sd1288281, -32'sd1257760, -32'sd175842, 32'sd76763, -32'sd1188877, -32'sd969599, -32'sd2051644, 32'sd442233, -32'sd236684, -32'sd823352, -32'sd1291536, -32'sd2604525, -32'sd834207, 32'sd0, 32'sd0, 32'sd0, -32'sd1148035, -32'sd502714, -32'sd487061, -32'sd6859, -32'sd1299102, -32'sd679599, -32'sd260980, -32'sd138480, -32'sd1510817, -32'sd1759038, -32'sd625173, -32'sd722056, 32'sd356607, -32'sd1485431, -32'sd614527, 32'sd251382, -32'sd511968, -32'sd1521460, -32'sd1162746, -32'sd1621889, -32'sd668879, 32'sd1156016, 32'sd468001, 32'sd173649, 32'sd1619379, 32'sd0, 32'sd0, 32'sd0, 32'sd151883, 32'sd66517, -32'sd1124063, -32'sd1398373, 32'sd577530, -32'sd2087707, -32'sd80416, -32'sd845755, -32'sd1666455, 32'sd516405, 32'sd692139, -32'sd887120, -32'sd1179350, 32'sd1022599, -32'sd262835, -32'sd416172, -32'sd537161, 32'sd369188, 32'sd1233099, -32'sd1560438, -32'sd1922566, -32'sd152348, 32'sd331143, 32'sd1214735, 32'sd624709, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1709521, 32'sd94455, -32'sd298114, -32'sd2266375, -32'sd833103, -32'sd1991697, -32'sd1888577, -32'sd2587518, -32'sd1596966, -32'sd2935937, -32'sd2912799, -32'sd512522, -32'sd1867111, -32'sd2732436, -32'sd1202191, -32'sd689793, 32'sd919856, 32'sd576395, -32'sd2012350, -32'sd349970, -32'sd1807588, 32'sd609536, 32'sd1347513, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd869309, 32'sd303495, 32'sd796326, 32'sd496453, 32'sd826037, -32'sd1149926, -32'sd1172053, -32'sd1402515, 32'sd66458, -32'sd1932642, -32'sd240971, -32'sd842594, -32'sd174082, -32'sd543562, 32'sd662347, 32'sd694738, 32'sd1014059, 32'sd547001, -32'sd284879, 32'sd52031, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd137959, -32'sd1263986, -32'sd566650, -32'sd1082046, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd955661, -32'sd923186, -32'sd554712, 32'sd48686, 32'sd444850, -32'sd680869, 32'sd780373, 32'sd493799, -32'sd280145, 32'sd497413, -32'sd781092, -32'sd956749, -32'sd1540047, -32'sd799270, -32'sd1913493, -32'sd210319, -32'sd99843, -32'sd19909, 32'sd145231, -32'sd862835, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd90959, -32'sd1066687, -32'sd1339917, -32'sd998824, -32'sd763170, 32'sd1388320, -32'sd707142, -32'sd207237, 32'sd80377, -32'sd1349958, -32'sd388082, -32'sd1144094, 32'sd520852, -32'sd1464350, -32'sd1490223, 32'sd201200, 32'sd314320, -32'sd1125353, -32'sd2170314, -32'sd1175977, -32'sd1554414, -32'sd292437, 32'sd971120, -32'sd203953, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1285237, -32'sd1147052, -32'sd436525, -32'sd176897, 32'sd655075, 32'sd316616, -32'sd188716, -32'sd137887, 32'sd703827, -32'sd2143831, -32'sd1239268, -32'sd2556756, -32'sd509675, -32'sd1635113, 32'sd721663, -32'sd646280, 32'sd1649073, -32'sd894046, -32'sd193940, 32'sd956061, -32'sd1781320, 32'sd161644, 32'sd430231, -32'sd1125282, -32'sd954535, 32'sd0, 32'sd0, -32'sd717859, -32'sd1148148, -32'sd1127901, -32'sd1919495, 32'sd1392305, 32'sd109425, -32'sd22015, -32'sd1234835, -32'sd2350135, -32'sd2922080, -32'sd2880530, -32'sd166137, 32'sd292641, -32'sd192954, -32'sd376933, 32'sd628325, 32'sd2812965, 32'sd2051791, -32'sd1011122, -32'sd598228, -32'sd699346, -32'sd668922, 32'sd1931059, 32'sd435635, 32'sd648435, -32'sd965271, 32'sd688620, 32'sd0, -32'sd1169092, -32'sd1002549, -32'sd1955496, -32'sd1874227, 32'sd695388, 32'sd13061, -32'sd256403, -32'sd1988241, -32'sd2187221, -32'sd1447891, -32'sd516979, -32'sd746035, -32'sd283830, -32'sd9475, 32'sd454469, 32'sd493243, 32'sd2259047, 32'sd730457, 32'sd1710748, -32'sd1001979, -32'sd1775354, -32'sd2276151, -32'sd2562730, -32'sd514203, 32'sd1614153, -32'sd786835, -32'sd708759, 32'sd0, -32'sd540870, -32'sd1667469, 32'sd193758, -32'sd919404, -32'sd1244395, -32'sd1745457, -32'sd1622181, -32'sd3284989, -32'sd2005021, -32'sd1564515, -32'sd450927, 32'sd383002, 32'sd142872, 32'sd1143525, 32'sd1686667, -32'sd144441, 32'sd1254675, 32'sd2009680, 32'sd227005, 32'sd409479, 32'sd1028823, 32'sd345923, 32'sd1908725, 32'sd2365219, -32'sd76088, 32'sd777767, -32'sd825954, -32'sd1145547, 32'sd599453, 32'sd555366, -32'sd347198, 32'sd1553392, -32'sd2393573, -32'sd2071555, -32'sd2008346, -32'sd2324768, -32'sd1612015, 32'sd2110828, 32'sd2218794, 32'sd3903130, 32'sd2440356, -32'sd143173, 32'sd1290796, 32'sd195579, -32'sd455912, 32'sd2880752, 32'sd887829, -32'sd1295293, -32'sd1137175, -32'sd667877, -32'sd924582, 32'sd2083723, -32'sd157811, -32'sd798499, 32'sd47080, 32'sd903149, -32'sd984900, -32'sd1362209, -32'sd186264, -32'sd1598525, -32'sd1344420, -32'sd2081162, -32'sd2050119, -32'sd880500, 32'sd310851, 32'sd2581009, 32'sd4322732, 32'sd2936350, 32'sd807494, 32'sd1264734, -32'sd460088, 32'sd692197, 32'sd599077, 32'sd777382, 32'sd1760599, 32'sd1703736, 32'sd479420, 32'sd251021, -32'sd91465, 32'sd160652, -32'sd779363, 32'sd642079, 32'sd529213, -32'sd621630, -32'sd1386930, -32'sd1380685, -32'sd976536, 32'sd2120591, 32'sd1010034, -32'sd1763656, -32'sd525409, 32'sd899320, 32'sd1252619, 32'sd1310981, 32'sd1349536, 32'sd1909989, 32'sd2037357, -32'sd336658, 32'sd99032, -32'sd447587, 32'sd672979, 32'sd864326, 32'sd881984, 32'sd3651331, 32'sd1589621, -32'sd966279, 32'sd1123453, 32'sd281203, 32'sd2158595, 32'sd171416, -32'sd680824, -32'sd1605263, 32'sd14398, 32'sd1052759, -32'sd109303, 32'sd487885, 32'sd1409501, 32'sd612856, 32'sd1602643, -32'sd600322, -32'sd396745, 32'sd479984, 32'sd1432563, 32'sd1229348, -32'sd44527, 32'sd154534, -32'sd2094310, -32'sd1514099, 32'sd875485, 32'sd1805644, 32'sd678313, 32'sd958267, 32'sd2529467, 32'sd177353, 32'sd660894, 32'sd1260706, 32'sd1224561, -32'sd1123592, 32'sd311227, -32'sd1337252, 32'sd1945590, 32'sd692781, -32'sd1327587, -32'sd1825863, -32'sd1111864, -32'sd772512, 32'sd1624903, -32'sd1583900, -32'sd420444, 32'sd1365211, 32'sd1178432, 32'sd2938006, 32'sd1645727, 32'sd77368, -32'sd733715, -32'sd350763, 32'sd1767092, 32'sd389196, -32'sd89469, 32'sd468816, 32'sd196726, 32'sd418331, 32'sd2031746, -32'sd341291, 32'sd437745, 32'sd855482, -32'sd2186185, -32'sd782235, 32'sd83856, -32'sd1172173, -32'sd1735325, 32'sd84757, -32'sd1066859, 32'sd788362, -32'sd1386579, 32'sd363183, -32'sd868536, 32'sd436648, 32'sd947293, 32'sd689319, 32'sd830269, -32'sd84032, -32'sd2901459, -32'sd77449, 32'sd2081461, 32'sd197592, 32'sd1465970, 32'sd172513, 32'sd464066, 32'sd1793796, -32'sd371256, 32'sd681971, -32'sd817923, 32'sd265739, -32'sd1641373, 32'sd811281, -32'sd857132, 32'sd333991, -32'sd577506, 32'sd1114887, -32'sd930342, -32'sd1981963, -32'sd1360802, 32'sd84978, 32'sd313234, 32'sd64534, -32'sd1358025, 32'sd201782, -32'sd697348, -32'sd1823068, -32'sd2045791, -32'sd1987312, -32'sd262960, -32'sd2063624, 32'sd646850, -32'sd597676, 32'sd293323, 32'sd137519, 32'sd1540747, 32'sd1055683, 32'sd684606, -32'sd1034209, -32'sd559736, -32'sd632849, 32'sd86748, 32'sd1164037, -32'sd575655, 32'sd2043051, 32'sd1295613, -32'sd1135748, -32'sd2140025, -32'sd2888709, -32'sd2823312, 32'sd124843, -32'sd2138056, 32'sd1690485, 32'sd377876, 32'sd637595, 32'sd955083, -32'sd943052, -32'sd865952, -32'sd1689208, -32'sd1000272, -32'sd498794, -32'sd27270, -32'sd7138, 32'sd1419366, 32'sd1480843, -32'sd2344913, 32'sd156955, -32'sd125454, -32'sd328147, -32'sd641440, 32'sd469554, -32'sd92576, 32'sd1187508, 32'sd416281, -32'sd3249842, -32'sd2440322, -32'sd1411470, 32'sd1317954, -32'sd54237, -32'sd2302559, -32'sd70308, 32'sd471524, 32'sd1145229, 32'sd1465907, 32'sd1045091, -32'sd1229263, -32'sd2918679, -32'sd2793902, -32'sd2784741, -32'sd69971, 32'sd2355731, 32'sd1322940, 32'sd2297446, -32'sd844768, -32'sd359171, -32'sd1672146, 32'sd671196, -32'sd1284991, 32'sd155784, -32'sd74305, 32'sd817909, -32'sd351230, -32'sd1900648, -32'sd2811306, 32'sd530508, 32'sd1077557, 32'sd2400559, -32'sd981621, 32'sd721903, -32'sd2592040, 32'sd592355, -32'sd661684, -32'sd2217679, -32'sd858656, -32'sd4047069, -32'sd2900079, -32'sd2482387, -32'sd286879, 32'sd367907, -32'sd766310, -32'sd588938, -32'sd1262223, 32'sd358915, -32'sd1000566, 32'sd0, 32'sd489716, -32'sd812176, 32'sd1650547, 32'sd1194812, -32'sd1144919, -32'sd209976, 32'sd407256, 32'sd34207, 32'sd409106, -32'sd344373, 32'sd665785, -32'sd1765382, -32'sd2010677, -32'sd2646831, -32'sd100172, -32'sd2734543, 32'sd133850, -32'sd456802, -32'sd2226234, -32'sd1765593, 32'sd839533, -32'sd451763, -32'sd643130, 32'sd1279756, 32'sd873109, -32'sd54766, -32'sd1057211, -32'sd1102212, -32'sd1146645, 32'sd1062408, -32'sd657088, -32'sd1011778, 32'sd171307, -32'sd1451787, -32'sd526197, -32'sd53974, 32'sd369784, 32'sd860002, -32'sd707670, -32'sd1956136, -32'sd1834837, -32'sd1021277, 32'sd18574, -32'sd263615, -32'sd36948, 32'sd1188732, -32'sd1669327, -32'sd1229036, 32'sd932526, 32'sd713660, 32'sd911288, 32'sd1065050, -32'sd1615357, -32'sd777034, -32'sd1627875, -32'sd591097, 32'sd225307, 32'sd222643, -32'sd882199, -32'sd297535, 32'sd1822834, -32'sd1420551, 32'sd310947, 32'sd2126, 32'sd525240, 32'sd2639871, -32'sd218397, -32'sd694675, -32'sd1176398, 32'sd406867, -32'sd51862, 32'sd1451119, 32'sd1997699, -32'sd106919, 32'sd529472, -32'sd800690, 32'sd197280, 32'sd981979, -32'sd1351287, -32'sd73259, -32'sd389527, -32'sd45173, -32'sd1104801, 32'sd0, -32'sd1360853, -32'sd1397999, 32'sd246017, 32'sd333781, 32'sd894199, -32'sd1236495, -32'sd1049028, 32'sd2994440, 32'sd1976995, 32'sd1585663, -32'sd1062725, -32'sd1155369, 32'sd393573, -32'sd2303664, -32'sd2119232, -32'sd1106999, -32'sd114803, -32'sd286625, -32'sd337604, -32'sd2168501, -32'sd2234424, -32'sd227429, 32'sd689189, -32'sd44056, 32'sd1059945, -32'sd895447, -32'sd183559, -32'sd584223, -32'sd1237847, -32'sd1497302, -32'sd863383, 32'sd1802239, 32'sd1871345, 32'sd1154068, 32'sd1012645, 32'sd2308068, 32'sd1883968, 32'sd704880, 32'sd1287961, -32'sd1614453, 32'sd1112006, -32'sd320173, -32'sd770409, -32'sd2278675, -32'sd664668, -32'sd961645, -32'sd415108, -32'sd2480633, -32'sd2051629, 32'sd1095237, -32'sd723732, -32'sd1947286, -32'sd436945, 32'sd2448261, 32'sd128218, -32'sd716223, -32'sd1478153, 32'sd736112, 32'sd371983, 32'sd1672631, 32'sd708852, 32'sd294434, 32'sd1549947, 32'sd944798, -32'sd8109, 32'sd2247088, 32'sd1581587, 32'sd588431, 32'sd2591681, 32'sd970474, -32'sd520982, -32'sd613515, -32'sd680978, -32'sd579704, -32'sd1738454, -32'sd2349911, -32'sd2421343, -32'sd1928502, -32'sd1118153, 32'sd635351, 32'sd1252351, 32'sd1055630, 32'sd704977, 32'sd0, -32'sd389029, 32'sd345867, -32'sd660195, -32'sd212278, 32'sd1261931, 32'sd46732, 32'sd843110, 32'sd2778243, -32'sd984694, -32'sd1301812, 32'sd1557464, 32'sd35638, -32'sd844983, 32'sd1395810, -32'sd417101, 32'sd1138417, -32'sd41021, -32'sd1168411, -32'sd755993, -32'sd2868317, -32'sd1160188, -32'sd619765, 32'sd181156, 32'sd1017110, 32'sd1287219, -32'sd834894, 32'sd0, 32'sd0, 32'sd0, 32'sd370113, 32'sd397112, 32'sd74667, 32'sd1182193, 32'sd100545, -32'sd708777, 32'sd1502323, -32'sd572203, -32'sd1308229, -32'sd300394, -32'sd567266, 32'sd295123, -32'sd781198, 32'sd353869, -32'sd885093, -32'sd3625039, -32'sd2696681, -32'sd1370581, -32'sd524979, -32'sd417761, 32'sd805358, -32'sd171081, 32'sd867214, -32'sd659722, -32'sd741842, 32'sd0, 32'sd0, 32'sd0, 32'sd299211, -32'sd982691, -32'sd1338787, -32'sd236905, 32'sd456700, -32'sd422499, 32'sd570496, -32'sd1420143, 32'sd1205351, 32'sd459335, -32'sd265365, -32'sd2245933, -32'sd1390158, -32'sd130414, -32'sd1081366, -32'sd558966, 32'sd289858, -32'sd1446060, -32'sd1519903, -32'sd1909805, -32'sd477905, -32'sd2085783, -32'sd1359470, -32'sd1156246, -32'sd888929, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd487027, 32'sd314339, -32'sd289038, -32'sd570268, -32'sd350970, 32'sd1888486, 32'sd982541, 32'sd1149958, 32'sd1775978, 32'sd668564, 32'sd999731, 32'sd78415, -32'sd573927, -32'sd148137, -32'sd472565, -32'sd2165321, 32'sd13997, -32'sd1686414, -32'sd1297529, 32'sd1410539, -32'sd306089, 32'sd488176, 32'sd318716, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd963282, -32'sd808058, 32'sd121476, 32'sd182790, 32'sd1057902, -32'sd1234457, -32'sd59840, -32'sd93066, 32'sd228271, 32'sd629602, 32'sd1040598, -32'sd1542743, 32'sd915711, 32'sd729074, -32'sd1843761, 32'sd19472, -32'sd1024187, -32'sd809400, 32'sd479406, 32'sd31485, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1325080, 32'sd405879, 32'sd166969, -32'sd1350784, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd600612, -32'sd1284623, 32'sd1067325, 32'sd2162929, -32'sd867192, 32'sd371823, 32'sd32970, 32'sd1349560, 32'sd1276922, -32'sd1749724, -32'sd422112, -32'sd302523, 32'sd488714, 32'sd321385, 32'sd927131, -32'sd727777, 32'sd373515, -32'sd872350, 32'sd477770, -32'sd171424, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd734727, -32'sd1048186, 32'sd1008797, -32'sd965800, -32'sd375856, 32'sd367516, -32'sd594999, -32'sd1692775, -32'sd1245588, 32'sd1509266, 32'sd205345, 32'sd184845, -32'sd704043, -32'sd244108, -32'sd1381835, 32'sd373112, -32'sd245357, -32'sd1020968, -32'sd105855, -32'sd894953, 32'sd585046, 32'sd207131, -32'sd745411, -32'sd392494, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd467788, 32'sd773555, 32'sd1618566, 32'sd1109200, 32'sd1861845, -32'sd1171995, -32'sd973404, -32'sd518647, -32'sd784924, 32'sd30744, -32'sd1805588, 32'sd671578, -32'sd168277, -32'sd1419892, 32'sd675886, -32'sd98796, 32'sd2339981, 32'sd831115, -32'sd1133333, 32'sd1282055, -32'sd559617, -32'sd125568, -32'sd989922, -32'sd1585737, 32'sd82043, 32'sd0, 32'sd0, -32'sd499940, -32'sd230313, -32'sd762136, 32'sd861121, 32'sd425882, -32'sd211612, 32'sd583640, -32'sd431274, 32'sd1183552, -32'sd1483997, -32'sd487831, -32'sd805803, 32'sd450862, -32'sd798701, -32'sd243867, 32'sd1275969, -32'sd1086177, 32'sd1407269, 32'sd393324, -32'sd812749, 32'sd1580871, 32'sd2130620, -32'sd135079, -32'sd32783, 32'sd173192, -32'sd1024262, 32'sd1277756, 32'sd0, -32'sd513501, 32'sd517558, 32'sd739660, -32'sd830347, -32'sd1333333, 32'sd704145, 32'sd2132252, 32'sd1664743, 32'sd1857671, 32'sd1849953, -32'sd828896, -32'sd1784611, -32'sd343514, -32'sd895911, -32'sd936432, 32'sd2316552, 32'sd2305913, -32'sd445753, 32'sd301503, -32'sd714701, 32'sd2344700, 32'sd2732381, 32'sd637453, -32'sd1034501, -32'sd1367446, 32'sd127646, -32'sd1320484, 32'sd0, -32'sd73205, -32'sd142237, -32'sd1052920, 32'sd853716, 32'sd673986, 32'sd588701, 32'sd2113116, 32'sd761916, 32'sd2211699, 32'sd1177591, -32'sd158214, -32'sd20335, 32'sd1022804, 32'sd1089926, -32'sd208800, -32'sd1172337, 32'sd1360764, 32'sd1785674, 32'sd664020, -32'sd560805, 32'sd692120, 32'sd1861837, 32'sd1900139, -32'sd165082, 32'sd986041, -32'sd194564, 32'sd807850, 32'sd549105, 32'sd98056, 32'sd172627, 32'sd37785, -32'sd1464563, 32'sd1213012, 32'sd440579, 32'sd136610, 32'sd3378415, 32'sd1347221, 32'sd1894776, -32'sd126528, 32'sd74656, -32'sd1502155, -32'sd309893, 32'sd1147198, 32'sd361434, 32'sd1142820, 32'sd1470970, 32'sd306241, -32'sd727844, 32'sd2303169, 32'sd1457864, 32'sd1638044, -32'sd478492, -32'sd729715, -32'sd843675, -32'sd833617, -32'sd587141, -32'sd384178, 32'sd321284, 32'sd603611, 32'sd56504, 32'sd138286, 32'sd1496744, 32'sd195465, 32'sd1171292, 32'sd1955395, -32'sd1616073, 32'sd299002, 32'sd273732, -32'sd14363, -32'sd481386, -32'sd681579, -32'sd1012342, 32'sd257814, -32'sd1106508, -32'sd532097, 32'sd888707, 32'sd177690, 32'sd174812, 32'sd748502, -32'sd1153703, 32'sd905944, -32'sd1952650, 32'sd617200, -32'sd445384, -32'sd1379106, -32'sd454889, 32'sd715145, -32'sd848628, -32'sd858902, -32'sd1661711, 32'sd1570710, 32'sd2740130, 32'sd1986340, 32'sd1860358, 32'sd28957, 32'sd413469, -32'sd1948436, -32'sd3932394, -32'sd811995, -32'sd1832367, -32'sd676177, -32'sd819004, 32'sd1362295, -32'sd1460279, 32'sd595976, 32'sd226654, 32'sd1207112, 32'sd732738, -32'sd477972, 32'sd695071, -32'sd310856, 32'sd178818, 32'sd542003, -32'sd153227, -32'sd984925, 32'sd152556, 32'sd1957049, -32'sd369269, 32'sd785021, -32'sd121347, 32'sd1450427, 32'sd1451560, 32'sd489138, -32'sd1237710, -32'sd1930685, -32'sd2334477, -32'sd1987225, -32'sd2365167, -32'sd1952530, 32'sd500376, -32'sd67405, -32'sd960646, 32'sd2424279, 32'sd2059311, 32'sd1798838, 32'sd1139775, 32'sd381843, 32'sd182680, 32'sd948085, -32'sd272179, -32'sd894318, -32'sd223845, -32'sd1477439, 32'sd1679843, 32'sd925283, -32'sd1404605, -32'sd441934, -32'sd871654, -32'sd659610, 32'sd1541871, 32'sd2092655, 32'sd101004, 32'sd958874, -32'sd77489, -32'sd3207819, -32'sd3389686, -32'sd1841439, -32'sd4109960, 32'sd1195638, 32'sd291681, -32'sd1342340, -32'sd2065799, -32'sd3246990, 32'sd478463, -32'sd857367, 32'sd1589742, -32'sd1715870, 32'sd629836, -32'sd1288269, 32'sd330672, -32'sd490346, -32'sd597681, 32'sd1596020, 32'sd798665, 32'sd529028, 32'sd624307, 32'sd1261769, 32'sd1962647, 32'sd2252048, 32'sd2226965, -32'sd904035, -32'sd1531769, -32'sd5397975, -32'sd2311603, -32'sd2690559, -32'sd556939, -32'sd639112, -32'sd1568782, 32'sd251130, -32'sd2707838, -32'sd1766193, 32'sd1222855, 32'sd699983, 32'sd1533524, -32'sd660916, 32'sd864177, -32'sd170168, -32'sd1712444, 32'sd204885, -32'sd676257, 32'sd837685, 32'sd517233, 32'sd303013, 32'sd565772, 32'sd2373115, 32'sd135433, 32'sd1815334, 32'sd1422440, 32'sd364236, -32'sd3802275, -32'sd3346529, -32'sd2250361, -32'sd2034201, 32'sd604030, -32'sd686391, -32'sd1309811, -32'sd1482100, -32'sd806873, 32'sd681670, -32'sd213965, 32'sd806777, 32'sd409304, 32'sd555045, 32'sd2032088, 32'sd466490, -32'sd64491, 32'sd812981, 32'sd805790, -32'sd1348810, 32'sd191901, -32'sd180368, -32'sd142170, -32'sd315984, 32'sd900403, 32'sd2282324, 32'sd1708631, 32'sd1142228, -32'sd2687620, -32'sd3467110, 32'sd333776, -32'sd929580, -32'sd191584, -32'sd2576269, -32'sd1799251, -32'sd30587, 32'sd138360, 32'sd1226531, -32'sd550445, 32'sd203507, 32'sd579246, 32'sd748675, -32'sd447941, 32'sd343311, 32'sd704227, -32'sd1536230, -32'sd522075, -32'sd284782, -32'sd139149, 32'sd768598, -32'sd93545, 32'sd443693, -32'sd855883, 32'sd1511596, 32'sd3323083, 32'sd2006363, 32'sd1059535, 32'sd1159691, 32'sd88563, -32'sd1037754, -32'sd1767937, -32'sd3299503, -32'sd3263742, -32'sd1516040, -32'sd1970183, -32'sd105437, -32'sd153982, 32'sd34009, -32'sd142703, 32'sd1046108, 32'sd601804, -32'sd830991, 32'sd1876697, -32'sd943665, -32'sd979853, -32'sd1153591, -32'sd749106, -32'sd2678353, -32'sd2396358, -32'sd505525, 32'sd278145, 32'sd53863, 32'sd784231, 32'sd2280202, 32'sd1358550, -32'sd543502, -32'sd1531246, -32'sd828356, -32'sd2590495, 32'sd166991, -32'sd2145914, -32'sd1101552, -32'sd792560, 32'sd645197, 32'sd98181, 32'sd876995, -32'sd1041549, -32'sd703987, 32'sd0, -32'sd113699, 32'sd702234, -32'sd1363613, -32'sd618530, -32'sd1085653, -32'sd664299, -32'sd3222199, -32'sd1990043, -32'sd1399956, 32'sd783901, 32'sd629270, 32'sd3698003, 32'sd3276505, 32'sd1475670, 32'sd8576, -32'sd537412, -32'sd3487376, -32'sd1841533, -32'sd709351, -32'sd729906, 32'sd817396, 32'sd2964235, 32'sd1719411, -32'sd26671, -32'sd1712607, -32'sd1218617, 32'sd102671, -32'sd506655, -32'sd194504, 32'sd334096, -32'sd872373, 32'sd260281, -32'sd1349525, -32'sd557747, -32'sd2910776, -32'sd1969999, -32'sd1007593, -32'sd1030849, -32'sd1289250, 32'sd2775097, 32'sd565611, -32'sd588136, 32'sd140755, -32'sd2446448, -32'sd2996991, -32'sd2293135, -32'sd681397, 32'sd861397, 32'sd417837, 32'sd1243377, -32'sd289896, 32'sd861023, 32'sd511744, -32'sd1250036, -32'sd466703, -32'sd657974, 32'sd139522, 32'sd181633, 32'sd1342470, -32'sd1427679, -32'sd164851, -32'sd1627667, 32'sd572509, -32'sd1791852, -32'sd2533504, -32'sd996010, -32'sd2044004, 32'sd3080938, -32'sd1509732, -32'sd3661597, -32'sd2713729, -32'sd919059, 32'sd1522708, 32'sd787791, 32'sd297202, 32'sd1183099, 32'sd2146892, -32'sd325889, -32'sd85932, 32'sd1483065, 32'sd96499, -32'sd903164, 32'sd52476, 32'sd0, 32'sd1554923, 32'sd849572, 32'sd671064, 32'sd108679, -32'sd894609, 32'sd941046, 32'sd25040, 32'sd316584, -32'sd1307794, 32'sd1278908, 32'sd758183, 32'sd1087823, -32'sd2192108, -32'sd2212401, 32'sd968690, 32'sd733750, 32'sd1798977, 32'sd2228822, 32'sd1135753, 32'sd2078444, 32'sd134319, -32'sd1154434, 32'sd288067, 32'sd1321660, 32'sd372327, -32'sd257681, 32'sd85361, -32'sd416519, 32'sd901526, 32'sd226515, -32'sd595539, 32'sd810656, -32'sd500240, -32'sd277818, 32'sd820655, 32'sd383232, 32'sd277075, 32'sd1702966, -32'sd595240, -32'sd1049725, -32'sd975642, -32'sd284602, 32'sd863477, 32'sd316176, 32'sd2155039, 32'sd1506803, 32'sd2207877, 32'sd2334820, 32'sd1887143, 32'sd967577, 32'sd286545, -32'sd538969, -32'sd202899, 32'sd871395, -32'sd658088, 32'sd7477, -32'sd915942, 32'sd799198, 32'sd1364847, 32'sd470399, -32'sd674200, 32'sd29082, 32'sd451242, 32'sd75632, 32'sd601055, -32'sd1292274, 32'sd1775995, 32'sd914566, 32'sd702909, 32'sd410572, 32'sd2203909, 32'sd1859895, 32'sd3822414, 32'sd2836998, 32'sd555961, 32'sd1234649, 32'sd700758, 32'sd874856, 32'sd129114, 32'sd135494, 32'sd423650, 32'sd168189, 32'sd706372, 32'sd0, 32'sd780427, -32'sd251648, 32'sd2218604, 32'sd239004, -32'sd657402, -32'sd654977, 32'sd524985, 32'sd367777, -32'sd990026, -32'sd519399, -32'sd123513, 32'sd2490149, 32'sd1724323, 32'sd912793, 32'sd3238342, 32'sd3521950, 32'sd2266036, 32'sd2356402, 32'sd791195, 32'sd1404811, 32'sd629574, 32'sd1399251, 32'sd847360, -32'sd520719, 32'sd1589661, 32'sd1209987, 32'sd0, 32'sd0, 32'sd0, -32'sd334996, 32'sd1255880, 32'sd21617, -32'sd764851, -32'sd2343461, -32'sd921627, 32'sd1465978, 32'sd1569434, 32'sd1372857, 32'sd2588101, 32'sd2966929, 32'sd3363766, 32'sd3264075, 32'sd4017719, 32'sd2330632, 32'sd1816681, 32'sd1531907, 32'sd1669687, 32'sd1083464, 32'sd1123578, 32'sd116324, -32'sd1390734, -32'sd1937742, -32'sd1782972, -32'sd303428, 32'sd0, 32'sd0, 32'sd0, 32'sd72592, 32'sd217547, -32'sd783226, -32'sd1265727, 32'sd433460, 32'sd376513, 32'sd2053342, 32'sd469786, -32'sd366196, 32'sd1776467, 32'sd1239229, 32'sd1552713, 32'sd1544893, 32'sd1209490, 32'sd1013552, 32'sd1212307, 32'sd224350, -32'sd1047941, -32'sd211195, -32'sd340971, 32'sd1108355, -32'sd1043201, -32'sd1144174, 32'sd347724, -32'sd592933, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd235621, 32'sd324350, -32'sd1207672, -32'sd1158174, 32'sd55155, -32'sd663258, 32'sd282148, -32'sd260931, -32'sd14301, 32'sd1248846, 32'sd1659091, -32'sd1211834, 32'sd795320, 32'sd256135, -32'sd191871, -32'sd137901, -32'sd1047930, 32'sd1069486, -32'sd141190, -32'sd388592, -32'sd310059, -32'sd39603, -32'sd647174, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd421121, 32'sd49052, -32'sd765953, 32'sd1350648, 32'sd418040, 32'sd1083736, -32'sd91925, -32'sd425356, 32'sd666852, 32'sd390016, -32'sd198506, -32'sd730709, -32'sd522348, 32'sd534663, 32'sd647792, -32'sd484103, -32'sd319606, -32'sd410141, -32'sd888010, 32'sd29427, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd79639, 32'sd1392654, 32'sd888930, 32'sd1359272, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd944939, 32'sd463405, 32'sd1271067, 32'sd1609889, 32'sd974819, 32'sd1387276, 32'sd316121, -32'sd889897, 32'sd1066806, 32'sd1570883, 32'sd158683, 32'sd950806, -32'sd1256460, 32'sd963946, 32'sd43095, -32'sd341724, 32'sd233613, 32'sd282560, -32'sd604891, 32'sd52856, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd225348, -32'sd655835, 32'sd175952, -32'sd408356, 32'sd770461, 32'sd1948067, 32'sd1420121, 32'sd2250267, 32'sd857504, -32'sd345463, -32'sd1211182, -32'sd1233230, 32'sd1608644, -32'sd200913, -32'sd1047772, 32'sd546902, -32'sd1853648, -32'sd1551618, -32'sd8610, 32'sd300418, 32'sd163971, 32'sd1917613, 32'sd383000, 32'sd843724, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd272792, 32'sd78544, -32'sd567413, 32'sd1063456, 32'sd757565, 32'sd127676, -32'sd849413, -32'sd150211, 32'sd726023, -32'sd274451, 32'sd999809, -32'sd2112055, 32'sd1100980, 32'sd81392, 32'sd2124588, 32'sd472748, -32'sd1813157, 32'sd419414, 32'sd537076, 32'sd1796834, -32'sd170843, -32'sd879105, -32'sd1336851, 32'sd1524180, 32'sd103101, 32'sd0, 32'sd0, 32'sd706629, -32'sd602298, 32'sd191759, -32'sd99307, -32'sd156493, -32'sd557704, -32'sd755046, -32'sd2179302, -32'sd3027918, -32'sd2261594, -32'sd2001773, -32'sd1874200, 32'sd85494, 32'sd1625495, 32'sd1558951, 32'sd1620479, 32'sd1322591, -32'sd639207, -32'sd1357879, 32'sd2041099, 32'sd1231167, -32'sd147233, -32'sd622534, -32'sd1618154, -32'sd986, 32'sd261474, -32'sd157990, 32'sd0, -32'sd51164, 32'sd537881, -32'sd1011580, 32'sd904270, 32'sd545677, 32'sd1177287, -32'sd2894664, -32'sd2288516, -32'sd3434790, -32'sd1433871, -32'sd873432, -32'sd845302, 32'sd1002102, 32'sd1250480, 32'sd505801, 32'sd2131429, 32'sd2606522, 32'sd787006, 32'sd1156537, 32'sd258868, -32'sd1730953, -32'sd1174142, -32'sd2063988, -32'sd1580985, 32'sd486258, 32'sd226454, -32'sd644650, 32'sd0, 32'sd319784, 32'sd619197, -32'sd1367210, -32'sd797232, 32'sd93310, -32'sd865038, -32'sd1260912, -32'sd2420495, -32'sd2607399, -32'sd1469261, -32'sd1581967, -32'sd683605, -32'sd380008, 32'sd181003, -32'sd874811, -32'sd1287613, 32'sd452992, -32'sd2222813, 32'sd76175, -32'sd545142, -32'sd1970322, 32'sd200325, 32'sd1238036, 32'sd925233, -32'sd173179, -32'sd146658, -32'sd915912, 32'sd604445, 32'sd510295, 32'sd1207602, -32'sd596224, 32'sd340287, -32'sd861772, -32'sd1411788, -32'sd1600257, -32'sd771210, -32'sd2901902, -32'sd911468, 32'sd87387, -32'sd643726, -32'sd601461, 32'sd601542, -32'sd1866286, -32'sd1906770, -32'sd135745, -32'sd2499101, -32'sd846395, -32'sd908763, -32'sd649534, 32'sd754344, -32'sd586552, 32'sd847643, -32'sd185351, 32'sd389054, -32'sd1129047, 32'sd216157, 32'sd392100, 32'sd975304, -32'sd3506593, -32'sd1016340, -32'sd921261, 32'sd36594, -32'sd1607787, -32'sd336001, -32'sd1100722, -32'sd3088864, -32'sd46538, 32'sd1357908, 32'sd1474750, 32'sd648842, 32'sd305573, -32'sd398571, -32'sd2297346, -32'sd2024607, -32'sd1915192, -32'sd501477, -32'sd342135, -32'sd2371251, -32'sd578166, -32'sd919377, 32'sd1857316, 32'sd1842354, 32'sd707448, 32'sd851405, -32'sd156637, -32'sd715492, -32'sd1451958, -32'sd416931, 32'sd861728, -32'sd970796, 32'sd283833, -32'sd1377886, 32'sd662211, -32'sd2768892, -32'sd1663245, 32'sd1466157, 32'sd25108, -32'sd659616, -32'sd19791, -32'sd254826, -32'sd1652623, -32'sd2039488, -32'sd1195339, -32'sd1289502, -32'sd1012741, -32'sd2158909, -32'sd2376577, -32'sd1846693, -32'sd1419863, 32'sd541449, -32'sd830688, -32'sd507725, -32'sd1155878, -32'sd1080995, -32'sd1150848, -32'sd75274, 32'sd966791, -32'sd280584, 32'sd1680500, 32'sd1178464, -32'sd655140, -32'sd744117, -32'sd1386291, -32'sd1483302, -32'sd1579000, -32'sd1500948, -32'sd1736522, -32'sd599702, -32'sd924931, -32'sd82073, -32'sd129274, -32'sd1672597, -32'sd2355071, -32'sd1237420, -32'sd3398705, 32'sd584166, 32'sd1001327, 32'sd2171253, -32'sd463318, -32'sd231350, 32'sd948718, -32'sd469582, -32'sd1003939, -32'sd353826, -32'sd530976, 32'sd2637684, -32'sd77226, 32'sd2121708, -32'sd790609, -32'sd785841, -32'sd1317188, 32'sd527876, -32'sd1876176, -32'sd1368699, -32'sd886187, -32'sd671512, 32'sd55885, 32'sd1717659, 32'sd1774781, -32'sd1146753, -32'sd549450, -32'sd2587646, 32'sd37224, 32'sd333395, 32'sd1181398, -32'sd473712, -32'sd1118937, -32'sd124280, -32'sd948031, -32'sd2002789, -32'sd269263, -32'sd161393, 32'sd75443, 32'sd1276955, 32'sd932876, 32'sd497510, -32'sd1508772, -32'sd1669655, 32'sd158933, 32'sd2147223, -32'sd1402806, -32'sd1822961, -32'sd1391334, 32'sd1169498, -32'sd150174, -32'sd86331, 32'sd1494617, 32'sd808279, -32'sd717346, 32'sd542305, -32'sd1876894, 32'sd170892, -32'sd253594, 32'sd456740, -32'sd418312, 32'sd544418, -32'sd617638, -32'sd2778906, 32'sd302718, -32'sd388020, 32'sd1791967, 32'sd1630551, 32'sd3195885, 32'sd1628948, 32'sd2131820, 32'sd2179976, 32'sd1828134, 32'sd2769604, 32'sd100396, -32'sd443123, -32'sd360488, 32'sd453889, -32'sd1976492, 32'sd1157073, 32'sd333311, -32'sd1425675, -32'sd695861, -32'sd2098493, 32'sd122530, 32'sd1612279, 32'sd878691, -32'sd203703, -32'sd150603, -32'sd401421, 32'sd689635, -32'sd840118, -32'sd1367660, -32'sd996527, 32'sd1275490, 32'sd536978, 32'sd3691735, 32'sd1495793, 32'sd2087523, 32'sd2034944, -32'sd113548, 32'sd1467652, -32'sd1160154, -32'sd660474, 32'sd1822095, 32'sd2090351, 32'sd136260, 32'sd830666, 32'sd291239, -32'sd2325727, 32'sd858338, 32'sd62777, 32'sd417923, 32'sd668695, 32'sd1620018, -32'sd215973, 32'sd1045400, -32'sd401005, -32'sd138184, 32'sd1589287, -32'sd1173736, 32'sd1042096, 32'sd1117676, 32'sd2997473, 32'sd2048791, 32'sd2991086, 32'sd1943787, 32'sd2396556, 32'sd243795, 32'sd1971649, -32'sd429040, 32'sd113849, 32'sd1260966, 32'sd1875021, 32'sd2945232, 32'sd2970555, 32'sd2290092, 32'sd392983, 32'sd454413, 32'sd446346, -32'sd140827, 32'sd426303, 32'sd2368943, 32'sd370959, 32'sd1632847, -32'sd499909, -32'sd558764, 32'sd38672, 32'sd1602103, -32'sd296367, -32'sd1737480, 32'sd355673, 32'sd495162, 32'sd2491216, 32'sd283348, -32'sd169619, 32'sd1155918, 32'sd1775089, -32'sd113163, 32'sd1124763, 32'sd4170073, 32'sd4173156, 32'sd2902626, 32'sd896601, 32'sd2385790, 32'sd1812022, 32'sd939533, 32'sd2097439, -32'sd211128, -32'sd503428, 32'sd1016260, 32'sd862436, 32'sd356214, 32'sd0, -32'sd341743, 32'sd1477706, -32'sd8976, 32'sd196110, 32'sd2009806, 32'sd430388, 32'sd64659, -32'sd125442, 32'sd788935, 32'sd2139951, 32'sd4172879, 32'sd2081641, 32'sd2663463, 32'sd2139329, 32'sd3990078, 32'sd1805195, -32'sd493941, 32'sd692650, -32'sd899047, 32'sd2498573, 32'sd2467675, 32'sd2854341, 32'sd354908, -32'sd1207759, 32'sd806346, 32'sd790553, -32'sd248545, -32'sd158971, -32'sd354057, -32'sd835913, 32'sd1931071, 32'sd1253519, 32'sd482884, -32'sd377205, 32'sd789520, 32'sd785783, 32'sd1199776, -32'sd128429, 32'sd3304347, 32'sd4776402, 32'sd1954753, 32'sd1057029, 32'sd1312999, 32'sd1859322, 32'sd1066657, -32'sd724405, 32'sd974013, 32'sd2653761, 32'sd2989493, 32'sd1007853, 32'sd1386665, 32'sd935201, 32'sd1182385, -32'sd515893, 32'sd364147, -32'sd250242, -32'sd1342055, 32'sd100992, 32'sd1499291, 32'sd2954359, 32'sd795466, 32'sd941941, 32'sd474981, -32'sd845850, 32'sd239506, 32'sd72237, 32'sd831165, 32'sd2674112, -32'sd161933, 32'sd202173, 32'sd890249, 32'sd2137328, 32'sd668893, 32'sd1263785, 32'sd733232, 32'sd1835211, 32'sd2515799, 32'sd1554866, 32'sd2791972, 32'sd2664558, 32'sd1134452, 32'sd1435145, -32'sd44371, 32'sd0, 32'sd753002, 32'sd1083716, 32'sd1282233, 32'sd522209, 32'sd394753, -32'sd671537, -32'sd478839, -32'sd1359167, -32'sd651690, -32'sd1420192, 32'sd329796, -32'sd225758, 32'sd437899, -32'sd1616660, -32'sd1233004, -32'sd383139, 32'sd1063708, 32'sd496291, -32'sd70131, 32'sd1881439, 32'sd2452086, 32'sd990788, 32'sd1625175, 32'sd1216104, 32'sd581839, 32'sd633598, 32'sd177049, 32'sd146751, 32'sd574780, -32'sd1705927, -32'sd1961917, 32'sd1069348, -32'sd228000, -32'sd65528, 32'sd479470, 32'sd278394, -32'sd281251, -32'sd1112787, -32'sd1803665, -32'sd732141, -32'sd1442498, -32'sd1592536, -32'sd2047179, 32'sd711858, -32'sd971664, -32'sd1744728, -32'sd1146930, 32'sd452804, -32'sd679681, 32'sd2586023, 32'sd1727806, 32'sd1218838, 32'sd1174091, -32'sd998847, 32'sd17103, -32'sd624408, -32'sd1407930, 32'sd786538, -32'sd2139166, 32'sd615393, -32'sd1363452, -32'sd163682, 32'sd68376, -32'sd354079, -32'sd1309317, -32'sd1872363, -32'sd269515, -32'sd1560199, -32'sd1926496, -32'sd1546274, -32'sd890809, 32'sd187431, -32'sd743498, -32'sd824210, -32'sd697921, 32'sd989822, -32'sd1290439, 32'sd569796, 32'sd73499, 32'sd1493950, -32'sd503220, 32'sd1270071, -32'sd383337, 32'sd0, -32'sd271152, -32'sd91397, 32'sd1761869, 32'sd2000324, -32'sd2427144, -32'sd1647561, -32'sd1647901, -32'sd2703684, -32'sd3118664, -32'sd2593236, -32'sd1776159, -32'sd2700538, -32'sd418468, -32'sd863383, -32'sd2385219, -32'sd1566909, -32'sd1053562, -32'sd799025, -32'sd955678, 32'sd99248, -32'sd846304, -32'sd344816, -32'sd796038, -32'sd257244, -32'sd318966, 32'sd352402, 32'sd0, 32'sd0, 32'sd0, 32'sd70891, 32'sd348803, 32'sd2517309, 32'sd1378956, -32'sd155850, -32'sd697547, -32'sd1506725, -32'sd426186, -32'sd1206183, 32'sd404062, -32'sd1117046, -32'sd174727, -32'sd115921, -32'sd771056, -32'sd253458, -32'sd1488154, 32'sd450773, 32'sd132092, -32'sd295957, 32'sd635098, -32'sd740281, 32'sd1098473, -32'sd806199, 32'sd179432, -32'sd444191, 32'sd0, 32'sd0, 32'sd0, 32'sd248136, -32'sd398402, -32'sd1281678, -32'sd732386, 32'sd255801, 32'sd256831, -32'sd284142, 32'sd542106, 32'sd669423, 32'sd553837, -32'sd1019119, -32'sd1934554, -32'sd616969, -32'sd1014932, 32'sd673048, -32'sd1116256, 32'sd516042, -32'sd660409, -32'sd904768, -32'sd1150620, -32'sd816492, 32'sd1430597, -32'sd362665, -32'sd27663, 32'sd889666, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd329231, 32'sd181140, -32'sd593252, -32'sd1393698, -32'sd1167186, 32'sd656136, -32'sd1406012, -32'sd1160218, -32'sd295774, 32'sd131301, -32'sd753319, -32'sd240866, 32'sd780814, -32'sd1223654, 32'sd1352893, 32'sd548978, 32'sd284558, -32'sd596367, 32'sd272562, -32'sd2114339, -32'sd771602, 32'sd4043, 32'sd371979, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd17642, 32'sd657798, 32'sd1236188, 32'sd354168, -32'sd211331, 32'sd378254, 32'sd12819, 32'sd1039515, -32'sd833700, 32'sd778321, -32'sd479572, 32'sd750546, 32'sd171194, 32'sd225109, -32'sd262435, 32'sd907668, 32'sd1214153, 32'sd1191576, -32'sd370014, 32'sd143742, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd78694, 32'sd328372, 32'sd915533, 32'sd1301460, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd280325, -32'sd489785, -32'sd1421387, 32'sd251240, 32'sd195571, -32'sd228273, 32'sd43905, 32'sd684262, -32'sd1299943, -32'sd33569, 32'sd522345, 32'sd731851, 32'sd545855, -32'sd1325726, 32'sd86831, -32'sd712347, -32'sd323300, 32'sd488221, -32'sd252171, 32'sd1046939, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd649813, 32'sd804934, 32'sd531851, 32'sd1433528, 32'sd529495, 32'sd193437, -32'sd1376559, -32'sd1177171, 32'sd792045, -32'sd1726362, 32'sd393411, 32'sd417288, -32'sd1264473, 32'sd247344, -32'sd101058, 32'sd1194037, 32'sd701358, 32'sd1328901, -32'sd869376, 32'sd860965, -32'sd602037, -32'sd1166816, 32'sd745147, 32'sd236563, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd660284, -32'sd853748, -32'sd197797, -32'sd1649953, 32'sd491372, 32'sd708802, -32'sd389942, 32'sd118403, 32'sd573089, -32'sd901712, -32'sd2546461, -32'sd1557922, 32'sd506055, 32'sd491677, 32'sd566183, 32'sd1021410, -32'sd87315, -32'sd569955, -32'sd596466, -32'sd971943, -32'sd469810, -32'sd183394, 32'sd720798, 32'sd436544, -32'sd2658672, 32'sd0, 32'sd0, 32'sd19046, 32'sd582087, 32'sd733081, 32'sd1840507, -32'sd172535, -32'sd771177, -32'sd1462254, -32'sd135153, 32'sd1261650, 32'sd2260648, 32'sd21852, 32'sd862173, 32'sd633482, -32'sd886709, -32'sd381001, -32'sd474993, -32'sd777132, 32'sd217612, 32'sd1575425, 32'sd2235821, -32'sd67312, 32'sd1867359, 32'sd433087, 32'sd849183, -32'sd151715, -32'sd467696, -32'sd651064, 32'sd0, 32'sd844533, -32'sd23410, -32'sd805182, -32'sd292452, 32'sd205878, 32'sd1365915, 32'sd56681, -32'sd384755, 32'sd1083198, 32'sd1560735, 32'sd839048, -32'sd392093, -32'sd3261798, -32'sd942534, -32'sd1039083, -32'sd1640348, -32'sd1125682, 32'sd329415, 32'sd1381274, 32'sd767995, 32'sd481250, 32'sd2627198, 32'sd484356, 32'sd1198502, 32'sd2079379, 32'sd129156, 32'sd724268, 32'sd0, 32'sd768119, -32'sd399625, -32'sd457700, 32'sd440813, 32'sd162135, 32'sd1092756, -32'sd631614, -32'sd555302, -32'sd1189674, -32'sd1234207, 32'sd146208, 32'sd732569, -32'sd825792, -32'sd595157, -32'sd3760587, -32'sd5150447, -32'sd1076776, -32'sd279796, -32'sd222016, 32'sd406019, -32'sd589018, 32'sd696539, 32'sd2104156, 32'sd2468682, -32'sd1047450, -32'sd439191, -32'sd114844, 32'sd178393, -32'sd226354, 32'sd865419, 32'sd298676, 32'sd3109946, 32'sd2107301, 32'sd865996, -32'sd630367, -32'sd2492097, 32'sd1289377, -32'sd512297, 32'sd2008752, 32'sd3211656, 32'sd3639355, -32'sd588182, -32'sd4239285, -32'sd3332453, 32'sd593199, 32'sd2335354, 32'sd946758, -32'sd1008859, 32'sd1005430, 32'sd1059308, 32'sd2886762, 32'sd2146711, -32'sd1022008, -32'sd102608, -32'sd2771001, 32'sd398292, -32'sd6698, 32'sd1112735, 32'sd503101, 32'sd415985, -32'sd2205962, 32'sd391811, 32'sd1722520, -32'sd1963814, -32'sd1302733, 32'sd470287, 32'sd161398, 32'sd2066871, 32'sd3055052, -32'sd2349538, -32'sd3886756, -32'sd2753632, 32'sd286634, 32'sd1325699, -32'sd650759, 32'sd310622, 32'sd1213233, -32'sd264320, -32'sd589981, 32'sd417426, -32'sd302415, -32'sd1811139, -32'sd203248, 32'sd1918651, -32'sd185421, 32'sd650915, 32'sd749017, -32'sd1462390, 32'sd412810, -32'sd978763, 32'sd785406, -32'sd1490600, -32'sd175316, -32'sd693361, 32'sd1572668, 32'sd1541336, 32'sd267248, -32'sd830059, -32'sd5129496, -32'sd4127521, -32'sd969252, 32'sd3251518, 32'sd2304821, 32'sd1334728, 32'sd3126296, -32'sd1485009, -32'sd831243, 32'sd481198, -32'sd1503022, 32'sd86690, 32'sd55383, -32'sd354770, 32'sd311812, -32'sd2244023, 32'sd468161, -32'sd337361, -32'sd302405, 32'sd7354, -32'sd622107, -32'sd1423708, -32'sd190847, -32'sd12392, 32'sd1755519, 32'sd2163479, 32'sd207415, -32'sd4523835, -32'sd7559432, -32'sd3216568, 32'sd1501854, 32'sd2404403, 32'sd1278825, -32'sd420801, 32'sd1678842, -32'sd236094, 32'sd404477, 32'sd258908, -32'sd967215, -32'sd1590738, -32'sd1835526, 32'sd267423, -32'sd123058, -32'sd654739, -32'sd260095, 32'sd604086, 32'sd196211, -32'sd297184, 32'sd895876, -32'sd313296, -32'sd396978, 32'sd551457, -32'sd507168, 32'sd1197822, -32'sd1712907, -32'sd3823373, -32'sd6757157, -32'sd935562, 32'sd2179022, 32'sd2162892, 32'sd1078371, 32'sd904353, 32'sd874823, 32'sd352959, -32'sd1689959, -32'sd669132, -32'sd2287383, 32'sd246749, 32'sd280235, 32'sd505997, 32'sd25884, -32'sd318599, -32'sd30012, -32'sd1212167, -32'sd859915, -32'sd748422, -32'sd1653861, -32'sd302283, 32'sd1486168, -32'sd15116, 32'sd230395, 32'sd762055, -32'sd235715, -32'sd2175141, -32'sd4890677, -32'sd490878, 32'sd2352454, 32'sd472618, 32'sd659999, 32'sd364262, 32'sd1236630, 32'sd2554064, -32'sd1948035, -32'sd82333, 32'sd267972, 32'sd571910, -32'sd788610, -32'sd57495, 32'sd483814, -32'sd1212376, -32'sd559622, 32'sd939227, -32'sd422033, 32'sd233603, -32'sd794736, 32'sd511915, 32'sd2416029, -32'sd470659, 32'sd1548727, 32'sd1359159, -32'sd1984713, -32'sd3074197, -32'sd3304781, 32'sd576813, 32'sd2458842, 32'sd1845090, 32'sd1422616, -32'sd581358, 32'sd2115952, 32'sd686941, -32'sd238607, -32'sd400148, -32'sd2244168, -32'sd587502, 32'sd1221636, -32'sd30323, 32'sd446113, -32'sd207388, -32'sd870299, -32'sd921898, 32'sd860298, -32'sd6651, 32'sd2485069, 32'sd565027, 32'sd1713008, 32'sd549268, 32'sd457541, 32'sd126214, -32'sd2362335, -32'sd2024846, -32'sd3368529, -32'sd8634, 32'sd2886669, -32'sd1465748, 32'sd626621, -32'sd158322, 32'sd2061318, -32'sd129066, -32'sd397141, 32'sd144230, 32'sd691098, -32'sd2078422, 32'sd1035008, -32'sd258402, 32'sd2338398, 32'sd1972026, -32'sd921480, 32'sd305151, -32'sd968340, -32'sd713782, 32'sd2715452, 32'sd1600491, 32'sd36352, 32'sd511637, 32'sd2131789, 32'sd1464013, -32'sd1255591, -32'sd662504, -32'sd662853, 32'sd801778, 32'sd1694832, -32'sd309691, 32'sd678406, -32'sd308342, -32'sd2056185, -32'sd59871, -32'sd1983775, 32'sd503909, 32'sd752706, -32'sd257457, 32'sd1035097, 32'sd812654, -32'sd393288, 32'sd473507, 32'sd566302, 32'sd823080, -32'sd1626295, 32'sd443422, -32'sd699061, -32'sd106872, -32'sd562433, -32'sd366092, -32'sd1692215, -32'sd1257465, -32'sd86646, -32'sd151264, 32'sd417066, -32'sd1077606, 32'sd885960, 32'sd141852, -32'sd212440, -32'sd1383496, -32'sd652317, -32'sd546309, -32'sd2243117, -32'sd1227882, -32'sd72320, -32'sd195101, -32'sd264427, 32'sd0, -32'sd388838, -32'sd748674, 32'sd800638, 32'sd1755036, -32'sd630896, 32'sd74372, 32'sd318320, 32'sd645463, -32'sd1510265, -32'sd845585, 32'sd105337, 32'sd677498, 32'sd3209484, -32'sd376270, 32'sd294056, -32'sd581086, 32'sd1302739, 32'sd130178, 32'sd1531111, -32'sd579323, -32'sd193121, 32'sd1436236, -32'sd659142, -32'sd2849831, 32'sd813958, 32'sd313110, 32'sd284269, -32'sd185448, -32'sd656386, -32'sd1204994, 32'sd354792, -32'sd111275, 32'sd136369, -32'sd246758, 32'sd420093, -32'sd310773, 32'sd1189190, 32'sd73666, 32'sd34277, 32'sd2202824, 32'sd737959, 32'sd1182659, -32'sd229905, 32'sd674429, -32'sd355114, 32'sd899953, 32'sd1512178, 32'sd33737, -32'sd534093, -32'sd1271357, -32'sd1748902, -32'sd807635, -32'sd107864, 32'sd1384431, 32'sd854858, 32'sd348528, 32'sd537906, 32'sd199947, 32'sd72984, 32'sd360360, 32'sd361016, -32'sd1001950, 32'sd223343, 32'sd811820, -32'sd11864, -32'sd630205, 32'sd245703, 32'sd1462865, 32'sd868275, 32'sd64490, 32'sd574318, 32'sd522243, 32'sd382283, 32'sd810034, -32'sd687539, 32'sd54098, 32'sd2314850, 32'sd245384, 32'sd254953, 32'sd378602, 32'sd182799, 32'sd26890, 32'sd2103612, 32'sd0, 32'sd472624, -32'sd542984, -32'sd1224259, -32'sd1739390, 32'sd183703, -32'sd199394, 32'sd185625, -32'sd1374413, -32'sd651221, 32'sd378167, 32'sd1782965, 32'sd280174, 32'sd1495686, 32'sd235773, -32'sd1229090, 32'sd1901033, 32'sd632352, 32'sd549831, 32'sd2218011, 32'sd256443, 32'sd2227860, 32'sd1474567, 32'sd890270, -32'sd971807, -32'sd219036, -32'sd391661, -32'sd388869, -32'sd338660, -32'sd127073, 32'sd1487868, -32'sd31779, -32'sd2105878, -32'sd420176, -32'sd521915, -32'sd838732, -32'sd307926, -32'sd588317, -32'sd537238, 32'sd1152432, 32'sd533622, 32'sd908286, -32'sd1225513, -32'sd1145864, 32'sd575163, 32'sd654163, 32'sd614792, 32'sd1403058, 32'sd2103216, -32'sd1376684, -32'sd505177, 32'sd477736, 32'sd437108, -32'sd941237, -32'sd230675, 32'sd1372875, 32'sd320591, 32'sd1250105, -32'sd83281, 32'sd1153305, -32'sd52342, -32'sd722026, -32'sd36852, -32'sd730792, 32'sd47280, -32'sd1494127, -32'sd1569830, 32'sd689061, 32'sd1886898, 32'sd198504, 32'sd208648, -32'sd746408, 32'sd641762, -32'sd1854233, -32'sd1884116, 32'sd901224, 32'sd1466375, 32'sd1755331, -32'sd541497, 32'sd1966847, 32'sd1537561, 32'sd374485, 32'sd968611, 32'sd467290, 32'sd0, -32'sd21199, -32'sd726560, -32'sd119689, -32'sd405829, -32'sd2355991, 32'sd175538, 32'sd1878085, -32'sd1728, -32'sd800062, -32'sd688638, 32'sd1358731, 32'sd1539066, 32'sd1011152, 32'sd897819, 32'sd1191454, 32'sd895733, -32'sd1056474, -32'sd2162723, -32'sd2258284, -32'sd24887, -32'sd283927, -32'sd177731, 32'sd1013752, 32'sd1879908, 32'sd1325162, -32'sd654452, 32'sd0, 32'sd0, 32'sd0, -32'sd117315, -32'sd201, -32'sd917036, -32'sd528781, -32'sd982018, 32'sd1043621, 32'sd1337826, -32'sd894041, -32'sd172335, 32'sd823279, 32'sd2779174, 32'sd940736, 32'sd1483354, -32'sd564332, 32'sd1770766, -32'sd1181961, -32'sd1951845, -32'sd1237950, -32'sd1247444, -32'sd905952, 32'sd492720, -32'sd443940, 32'sd481839, 32'sd122020, -32'sd378136, 32'sd0, 32'sd0, 32'sd0, -32'sd402746, -32'sd675498, 32'sd83244, -32'sd1888181, 32'sd2207627, -32'sd745034, 32'sd472159, -32'sd605930, 32'sd1330367, 32'sd26074, 32'sd1353102, -32'sd1690640, -32'sd17231, 32'sd36465, 32'sd858929, -32'sd782877, -32'sd1565774, -32'sd191291, -32'sd317017, -32'sd801205, -32'sd371366, 32'sd1004516, -32'sd1942799, 32'sd562530, 32'sd1438312, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd639099, -32'sd332208, -32'sd1191540, -32'sd263474, -32'sd1002808, 32'sd313371, -32'sd1404564, -32'sd1463775, -32'sd1246323, -32'sd1000151, 32'sd139215, -32'sd1565483, 32'sd670747, -32'sd1363235, 32'sd1166886, 32'sd919505, -32'sd1944537, -32'sd1534845, -32'sd475745, 32'sd637172, 32'sd125150, 32'sd1579412, 32'sd793593, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd359592, 32'sd685272, 32'sd411202, 32'sd655415, -32'sd1141738, 32'sd1010010, 32'sd288255, 32'sd231100, -32'sd224259, 32'sd346474, 32'sd157349, -32'sd523223, -32'sd1731144, -32'sd280116, 32'sd233443, 32'sd877945, -32'sd398121, 32'sd864453, -32'sd973008, 32'sd227264, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd412298, -32'sd845594, -32'sd523236, -32'sd80830, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1287517, -32'sd1404415, -32'sd788765, 32'sd545747, 32'sd332022, -32'sd121055, -32'sd560759, -32'sd413265, -32'sd1734443, 32'sd444794, -32'sd317080, -32'sd2364159, -32'sd1190745, 32'sd1732558, 32'sd1714950, 32'sd1067708, 32'sd486555, -32'sd645791, -32'sd1400438, -32'sd162799, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1131134, -32'sd458999, 32'sd1034495, -32'sd451020, 32'sd928999, 32'sd112770, 32'sd353661, 32'sd1250371, 32'sd712822, -32'sd2180547, -32'sd199618, 32'sd781490, -32'sd2019303, -32'sd131622, -32'sd445702, -32'sd1277814, 32'sd38783, 32'sd296188, -32'sd108890, 32'sd381037, 32'sd1177748, 32'sd1192924, -32'sd1008881, -32'sd1180661, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1294179, -32'sd809581, 32'sd1466005, -32'sd679646, 32'sd182124, 32'sd1027934, -32'sd1296305, 32'sd156399, 32'sd1194190, -32'sd350514, -32'sd773263, 32'sd1253286, 32'sd4227, -32'sd614033, 32'sd18565, -32'sd126902, 32'sd2253201, 32'sd457829, -32'sd2148714, 32'sd1673033, 32'sd801706, -32'sd568920, -32'sd934625, -32'sd603767, -32'sd860347, 32'sd0, 32'sd0, -32'sd618911, -32'sd973237, -32'sd1317839, 32'sd646618, -32'sd1477795, 32'sd568776, 32'sd1060074, -32'sd1166678, -32'sd740157, -32'sd1003154, -32'sd1078556, 32'sd919918, 32'sd218316, 32'sd810175, 32'sd1843195, -32'sd399683, -32'sd1312405, 32'sd1405394, 32'sd1160661, 32'sd1187065, 32'sd1863755, -32'sd521017, -32'sd1464074, -32'sd2420830, -32'sd1047245, -32'sd71890, -32'sd800846, 32'sd0, -32'sd872709, -32'sd1016035, 32'sd72917, 32'sd752968, -32'sd401941, -32'sd73484, 32'sd94281, 32'sd89835, 32'sd62407, 32'sd54193, 32'sd719091, -32'sd732904, 32'sd2560128, 32'sd1366726, 32'sd1969027, 32'sd291194, -32'sd162517, -32'sd496599, 32'sd1454196, 32'sd1304522, 32'sd175010, -32'sd777028, -32'sd2603969, -32'sd1300612, -32'sd1559059, -32'sd450963, -32'sd1464519, 32'sd0, 32'sd911330, -32'sd861331, -32'sd401836, 32'sd76808, -32'sd940885, -32'sd1645804, 32'sd1550450, 32'sd580618, -32'sd1392800, -32'sd767118, -32'sd288495, -32'sd1052848, -32'sd493361, -32'sd82129, -32'sd755667, 32'sd145890, 32'sd646549, 32'sd1748711, 32'sd1180641, 32'sd1323100, -32'sd493286, 32'sd1557632, -32'sd391129, -32'sd460610, -32'sd50574, -32'sd128466, 32'sd112711, -32'sd562798, -32'sd940290, -32'sd330875, -32'sd1050129, 32'sd1000937, -32'sd1506434, -32'sd1535508, -32'sd2902327, 32'sd248532, -32'sd360467, -32'sd717453, -32'sd826933, -32'sd2497596, -32'sd2333950, -32'sd1607610, 32'sd1069109, 32'sd41549, 32'sd2392093, 32'sd2112435, 32'sd482384, 32'sd1221523, 32'sd178675, 32'sd1311836, -32'sd140773, -32'sd1633311, 32'sd93261, -32'sd547403, -32'sd515984, 32'sd1407481, -32'sd1624009, -32'sd1307236, -32'sd781559, -32'sd542723, -32'sd2106182, 32'sd120592, -32'sd1078891, -32'sd1042338, -32'sd1764905, -32'sd716468, 32'sd1349289, 32'sd451040, -32'sd274835, 32'sd1229353, -32'sd921971, 32'sd1133911, 32'sd2077220, 32'sd816313, 32'sd2147671, 32'sd1304012, 32'sd141632, -32'sd407111, 32'sd1084431, 32'sd638518, 32'sd1001662, 32'sd318746, 32'sd397267, -32'sd4747, -32'sd504926, 32'sd768700, 32'sd254148, -32'sd676424, -32'sd2287027, -32'sd1047766, -32'sd523150, -32'sd1599430, -32'sd765269, 32'sd473730, 32'sd2785118, 32'sd1904209, 32'sd2511586, 32'sd1816212, -32'sd171326, -32'sd2199737, -32'sd1794394, -32'sd2731659, 32'sd312189, 32'sd2160820, 32'sd1898035, -32'sd541111, 32'sd300762, 32'sd551453, 32'sd2117352, 32'sd904664, -32'sd1586592, 32'sd173222, 32'sd30105, 32'sd113715, -32'sd834832, 32'sd408012, -32'sd597278, -32'sd1376670, -32'sd1975442, -32'sd2119245, 32'sd2083847, 32'sd2062237, -32'sd481631, 32'sd127558, 32'sd2787341, 32'sd2677643, -32'sd432806, -32'sd543305, -32'sd199607, -32'sd166660, -32'sd815680, 32'sd1375611, 32'sd406093, 32'sd723014, 32'sd22707, 32'sd1015672, 32'sd901718, 32'sd950552, -32'sd495918, 32'sd751005, 32'sd405672, 32'sd1508535, -32'sd142263, -32'sd507372, 32'sd191435, -32'sd133188, 32'sd1587477, 32'sd309765, 32'sd897586, 32'sd2430378, 32'sd1997800, 32'sd1073395, 32'sd1562048, 32'sd2677063, 32'sd1106700, 32'sd1310744, -32'sd736649, -32'sd2335479, -32'sd693134, 32'sd1435664, 32'sd2935298, 32'sd1387292, 32'sd1133813, 32'sd11613, 32'sd1527601, -32'sd1071060, -32'sd1263787, 32'sd182642, -32'sd1425784, -32'sd1057857, 32'sd100365, 32'sd113932, -32'sd1127306, 32'sd1267765, 32'sd1363135, 32'sd591961, 32'sd2375166, 32'sd1434696, 32'sd1679346, 32'sd867492, 32'sd3702404, 32'sd1851656, 32'sd1162624, 32'sd2026374, 32'sd1201682, 32'sd9978, 32'sd681018, 32'sd638701, 32'sd1119882, 32'sd249855, 32'sd1736054, -32'sd784109, 32'sd172638, -32'sd173344, 32'sd666877, 32'sd865779, -32'sd1491566, -32'sd1859519, -32'sd768133, -32'sd2751669, -32'sd270691, 32'sd1042712, 32'sd1750003, 32'sd852543, 32'sd2226262, -32'sd358820, 32'sd1300688, 32'sd1259557, 32'sd1701594, 32'sd993323, 32'sd1235480, 32'sd2452512, 32'sd624814, 32'sd507506, -32'sd708561, -32'sd415543, -32'sd451678, -32'sd353009, -32'sd1136955, -32'sd961236, 32'sd1048791, -32'sd958217, -32'sd466684, -32'sd994702, -32'sd1360484, -32'sd930132, 32'sd636251, 32'sd311763, -32'sd173733, -32'sd524521, 32'sd1580231, 32'sd2240617, -32'sd277919, 32'sd792186, 32'sd1457030, 32'sd629441, 32'sd900112, 32'sd62764, 32'sd495682, 32'sd657518, 32'sd1972587, 32'sd530944, -32'sd1570645, -32'sd1982213, -32'sd892419, -32'sd524602, 32'sd283921, -32'sd2062362, -32'sd1182187, 32'sd693717, 32'sd130016, -32'sd1409520, -32'sd900788, -32'sd1197912, -32'sd855809, 32'sd233030, 32'sd385340, -32'sd60111, 32'sd2174566, 32'sd412063, 32'sd1865583, -32'sd531877, 32'sd1350328, 32'sd2168942, 32'sd1226013, -32'sd1014978, -32'sd1152451, -32'sd499562, -32'sd693244, -32'sd1809956, -32'sd1379488, -32'sd1792160, -32'sd533858, -32'sd1161427, 32'sd73284, -32'sd1409231, -32'sd578320, -32'sd456501, -32'sd49990, 32'sd904275, -32'sd1567781, -32'sd331847, -32'sd2245710, -32'sd2575629, 32'sd287935, 32'sd469953, 32'sd2729341, 32'sd2671513, 32'sd3590681, 32'sd3252928, 32'sd2398577, 32'sd572971, -32'sd1189703, -32'sd4163122, -32'sd3000364, -32'sd2006313, -32'sd724834, -32'sd3077895, -32'sd1438651, -32'sd826105, -32'sd996095, 32'sd289733, -32'sd343341, 32'sd106537, -32'sd573068, -32'sd873296, -32'sd624825, 32'sd0, 32'sd793238, -32'sd249655, -32'sd2557734, -32'sd352296, -32'sd1084872, -32'sd271094, 32'sd2051815, 32'sd2022851, 32'sd2829580, 32'sd4977337, 32'sd552243, -32'sd1418858, -32'sd4688162, -32'sd3813355, -32'sd2716442, -32'sd564763, -32'sd2347162, -32'sd1789645, -32'sd453697, 32'sd964220, -32'sd1009644, 32'sd103264, 32'sd65164, -32'sd162431, -32'sd2444181, -32'sd1815468, -32'sd1325604, -32'sd746184, -32'sd1118590, 32'sd649694, -32'sd1381170, 32'sd415787, -32'sd638465, 32'sd85226, 32'sd2002202, 32'sd618102, 32'sd3019523, 32'sd2897431, 32'sd109078, -32'sd3361834, -32'sd3031804, -32'sd2240082, -32'sd709920, -32'sd606091, -32'sd1862907, -32'sd1699066, 32'sd45844, -32'sd1216936, -32'sd610126, -32'sd2328653, -32'sd1518749, -32'sd355921, -32'sd1317045, -32'sd775628, -32'sd1580999, -32'sd540393, -32'sd1044131, -32'sd30403, 32'sd75449, -32'sd726985, 32'sd1205105, -32'sd1229740, 32'sd1055403, 32'sd1485867, 32'sd1207373, 32'sd2255040, 32'sd599263, -32'sd4443560, -32'sd3369607, -32'sd1988174, 32'sd848586, -32'sd10827, -32'sd1436872, -32'sd1438448, -32'sd1277608, -32'sd880562, 32'sd1458592, 32'sd929698, 32'sd84185, 32'sd217081, -32'sd842515, -32'sd2047239, -32'sd1321909, 32'sd0, 32'sd716300, -32'sd1039572, 32'sd595999, -32'sd317499, 32'sd2281616, 32'sd362017, 32'sd745800, 32'sd1400897, 32'sd1467920, 32'sd641438, 32'sd1205541, -32'sd3067309, -32'sd2720452, -32'sd617860, -32'sd1091678, -32'sd1491309, -32'sd2641454, -32'sd810808, 32'sd463098, 32'sd769021, 32'sd180250, -32'sd849973, -32'sd1775471, -32'sd457752, -32'sd207266, -32'sd1721979, -32'sd956219, -32'sd325944, 32'sd355794, -32'sd1454665, 32'sd1319627, -32'sd861018, -32'sd501114, 32'sd2351858, 32'sd2046990, 32'sd738562, 32'sd1271773, 32'sd2377675, 32'sd647745, -32'sd740227, -32'sd1734837, -32'sd163520, -32'sd111634, -32'sd380055, 32'sd430460, -32'sd65852, 32'sd455252, 32'sd1543839, -32'sd58233, 32'sd1007413, -32'sd1657729, 32'sd262600, 32'sd453623, 32'sd149043, 32'sd693802, -32'sd999304, -32'sd1265368, -32'sd1690892, 32'sd1013365, -32'sd568531, 32'sd263043, 32'sd622978, 32'sd632897, 32'sd1559768, -32'sd100574, 32'sd1799970, 32'sd2724378, 32'sd1654543, 32'sd431252, 32'sd673921, 32'sd881116, -32'sd1294721, 32'sd147402, -32'sd591535, -32'sd931832, 32'sd283851, 32'sd592124, 32'sd1290713, -32'sd901190, -32'sd2338763, -32'sd287359, -32'sd1130181, 32'sd789634, 32'sd0, -32'sd1105141, -32'sd8376, -32'sd487240, -32'sd601926, -32'sd734302, 32'sd48113, 32'sd1131719, 32'sd519808, 32'sd1663224, -32'sd1004015, -32'sd281359, 32'sd1907586, 32'sd1255906, 32'sd1383537, 32'sd672890, -32'sd1694982, 32'sd854487, -32'sd935687, 32'sd330726, -32'sd2269762, -32'sd992833, 32'sd1258848, -32'sd2005933, -32'sd1108046, -32'sd828019, -32'sd1532570, 32'sd0, 32'sd0, 32'sd0, -32'sd155324, -32'sd389211, -32'sd1927573, -32'sd558770, 32'sd254564, 32'sd72682, -32'sd504131, -32'sd179299, 32'sd856319, 32'sd2604894, 32'sd3937711, 32'sd1455975, -32'sd810410, -32'sd674200, -32'sd416415, 32'sd1009642, -32'sd560179, -32'sd1582673, -32'sd2439658, -32'sd1122351, 32'sd381187, -32'sd873718, -32'sd1076231, -32'sd1428786, -32'sd1248384, 32'sd0, 32'sd0, 32'sd0, 32'sd277585, 32'sd36250, -32'sd685693, -32'sd599026, 32'sd1857084, -32'sd817639, 32'sd1126407, 32'sd931744, 32'sd1282010, 32'sd1514838, 32'sd1100637, 32'sd1138609, 32'sd353838, -32'sd1233493, 32'sd865246, -32'sd319928, -32'sd606237, 32'sd365470, 32'sd604101, -32'sd921361, -32'sd1062998, -32'sd1335223, -32'sd1851202, -32'sd1420036, -32'sd1174358, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd806155, -32'sd1249454, -32'sd253546, -32'sd1135964, -32'sd698575, 32'sd35710, 32'sd529989, -32'sd96924, 32'sd849519, 32'sd422221, 32'sd1081714, 32'sd1763208, -32'sd2320626, -32'sd1907769, -32'sd301858, -32'sd200287, 32'sd224046, -32'sd1374234, -32'sd1480500, -32'sd183141, -32'sd1637580, -32'sd1164757, -32'sd1296193, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd135100, -32'sd1286983, -32'sd657445, -32'sd1036785, -32'sd1301049, -32'sd629276, 32'sd694694, 32'sd1025766, 32'sd780669, 32'sd1560191, -32'sd253921, 32'sd1374994, 32'sd1004939, 32'sd759934, -32'sd1428070, 32'sd195747, -32'sd1291410, -32'sd1131582, -32'sd346150, -32'sd1027331, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd870875, -32'sd525359, -32'sd200896, -32'sd309480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd559557, -32'sd48502, -32'sd614032, -32'sd347697, 32'sd151384, -32'sd78681, -32'sd87544, 32'sd460955, 32'sd138891, 32'sd766732, -32'sd72043, -32'sd686263, 32'sd491724, -32'sd1076693, 32'sd998884, -32'sd1003961, 32'sd125631, 32'sd270375, -32'sd634951, -32'sd327342, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd324473, -32'sd14568, 32'sd413761, -32'sd1043445, -32'sd232681, 32'sd435361, 32'sd1650540, 32'sd783585, -32'sd1026250, -32'sd269604, -32'sd658899, 32'sd436965, -32'sd246292, -32'sd384504, -32'sd652220, 32'sd70854, 32'sd1862674, 32'sd1643079, 32'sd1181267, -32'sd779286, 32'sd224035, 32'sd576541, 32'sd1040399, 32'sd290167, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd892312, 32'sd336782, 32'sd917158, -32'sd545490, -32'sd724248, 32'sd1024029, -32'sd238412, -32'sd1157110, -32'sd116856, 32'sd2360812, 32'sd440383, 32'sd790517, 32'sd228916, -32'sd746041, -32'sd1643831, 32'sd416824, 32'sd104162, -32'sd1838653, -32'sd707982, 32'sd392167, -32'sd65180, -32'sd351373, 32'sd1070028, 32'sd210820, 32'sd8248, 32'sd0, 32'sd0, -32'sd43365, 32'sd27936, -32'sd1257363, -32'sd1025248, -32'sd6548, -32'sd1228866, -32'sd1269435, -32'sd1984193, -32'sd294340, -32'sd622074, -32'sd849749, -32'sd1723405, 32'sd1161075, -32'sd123482, 32'sd1069723, -32'sd989032, 32'sd532595, 32'sd1698845, -32'sd582051, 32'sd68678, 32'sd138828, 32'sd2556531, 32'sd1412863, -32'sd1013750, -32'sd1360614, -32'sd977217, -32'sd309644, 32'sd0, 32'sd203969, -32'sd70627, -32'sd343373, 32'sd1127150, 32'sd1502744, 32'sd844222, 32'sd18539, 32'sd674210, -32'sd200229, -32'sd780556, 32'sd353977, -32'sd126008, 32'sd2630580, 32'sd2621560, -32'sd1562247, 32'sd98861, 32'sd2201960, 32'sd316379, 32'sd163626, 32'sd943748, 32'sd1043220, 32'sd571394, 32'sd97261, -32'sd1979806, 32'sd395319, -32'sd1137668, 32'sd961175, 32'sd0, -32'sd93596, -32'sd257845, -32'sd263578, -32'sd75316, -32'sd649933, -32'sd1863257, -32'sd732394, -32'sd2302633, -32'sd246887, -32'sd53088, -32'sd106628, 32'sd1155941, 32'sd2308337, 32'sd1366704, 32'sd3124746, 32'sd2093571, 32'sd4125002, 32'sd2712390, 32'sd1321854, -32'sd89742, -32'sd570108, -32'sd633835, -32'sd2186945, -32'sd1515222, -32'sd1971510, -32'sd1139387, 32'sd1075743, 32'sd37048, -32'sd806397, -32'sd28007, -32'sd579446, 32'sd1036565, -32'sd1202928, 32'sd587593, 32'sd1195273, 32'sd1533047, 32'sd1862856, 32'sd537018, 32'sd448921, 32'sd1694890, 32'sd1017403, 32'sd738414, 32'sd1333352, 32'sd2717619, 32'sd807385, 32'sd2231238, 32'sd1869125, 32'sd1715199, -32'sd630242, -32'sd1234080, -32'sd642567, 32'sd111133, -32'sd189169, 32'sd537260, 32'sd1760962, -32'sd59422, 32'sd350058, 32'sd367359, 32'sd439720, -32'sd890994, 32'sd607347, -32'sd175688, 32'sd240744, -32'sd480686, 32'sd543847, 32'sd1110546, 32'sd1235438, 32'sd679983, 32'sd324508, -32'sd90454, -32'sd125302, -32'sd722792, -32'sd955596, 32'sd72549, -32'sd989351, 32'sd513656, -32'sd118326, -32'sd1834742, -32'sd1978225, -32'sd2340852, -32'sd570661, 32'sd243561, -32'sd610677, -32'sd59715, -32'sd678326, 32'sd843419, -32'sd916810, 32'sd477472, -32'sd162980, -32'sd1088356, -32'sd670975, -32'sd1111228, -32'sd811957, 32'sd1126171, -32'sd808304, -32'sd1640530, -32'sd2367783, -32'sd1110128, -32'sd782937, -32'sd1136512, -32'sd750531, -32'sd732919, 32'sd131817, -32'sd55672, -32'sd1853769, -32'sd2418070, -32'sd3190909, -32'sd815569, -32'sd1230640, -32'sd89446, -32'sd989839, -32'sd692177, 32'sd370836, 32'sd1293198, -32'sd2080320, -32'sd459595, -32'sd13833, -32'sd169549, -32'sd303323, 32'sd729947, -32'sd1245317, 32'sd718469, 32'sd565347, -32'sd3022459, -32'sd1726843, -32'sd1639051, -32'sd1675793, -32'sd1313959, -32'sd947107, 32'sd1879297, 32'sd179998, -32'sd590746, -32'sd1893200, -32'sd680268, -32'sd657095, 32'sd53382, -32'sd1090942, -32'sd160898, -32'sd604773, 32'sd814774, -32'sd957447, -32'sd2119408, 32'sd28262, -32'sd1259066, -32'sd583183, 32'sd16095, 32'sd1223407, 32'sd2128524, 32'sd584349, -32'sd1078957, 32'sd441868, -32'sd938165, -32'sd84218, -32'sd1346386, -32'sd1786037, 32'sd300338, 32'sd559084, 32'sd1227714, -32'sd550614, -32'sd366034, -32'sd1048313, 32'sd455147, 32'sd1507668, 32'sd1001672, -32'sd285153, 32'sd992482, 32'sd1050995, -32'sd517477, 32'sd319618, 32'sd1217227, -32'sd993770, 32'sd992025, 32'sd68435, -32'sd976783, 32'sd1887532, 32'sd1037560, -32'sd540865, 32'sd1563163, 32'sd1333774, -32'sd117664, -32'sd593849, -32'sd1877336, -32'sd1116547, -32'sd147951, -32'sd1491774, -32'sd1104540, -32'sd1324015, -32'sd540015, -32'sd500648, -32'sd55852, 32'sd224321, -32'sd1962052, -32'sd2517246, -32'sd1394847, -32'sd167841, -32'sd529399, 32'sd46458, 32'sd1387647, 32'sd234729, 32'sd89567, 32'sd2436316, -32'sd202544, 32'sd92153, 32'sd692448, -32'sd30617, 32'sd120615, -32'sd789109, -32'sd117551, -32'sd710319, -32'sd2317448, -32'sd1372654, -32'sd655612, -32'sd1897088, 32'sd242781, 32'sd233030, -32'sd645250, -32'sd1542100, -32'sd2436406, -32'sd1079315, 32'sd254118, 32'sd423680, -32'sd1429425, 32'sd289098, 32'sd783844, 32'sd1196082, -32'sd386707, -32'sd1424755, 32'sd268437, 32'sd641442, -32'sd220681, -32'sd2013639, -32'sd760679, 32'sd514355, 32'sd2772847, 32'sd1121186, -32'sd363226, 32'sd1256788, 32'sd391155, -32'sd2213645, -32'sd1504615, -32'sd697170, -32'sd78375, -32'sd1472699, 32'sd325027, 32'sd798877, 32'sd1076052, 32'sd572290, -32'sd915201, 32'sd1362192, -32'sd1133220, -32'sd1286057, 32'sd1560077, -32'sd806850, -32'sd1182211, -32'sd593019, -32'sd2080018, -32'sd1258347, -32'sd2659227, -32'sd1000470, -32'sd1899602, 32'sd774150, 32'sd846116, 32'sd1044629, -32'sd203026, 32'sd2001511, -32'sd329523, 32'sd1708793, 32'sd427230, -32'sd551988, 32'sd428783, -32'sd2319250, -32'sd1149254, 32'sd1973295, 32'sd1114787, 32'sd735103, 32'sd67348, 32'sd106751, 32'sd1105881, -32'sd755306, 32'sd66044, -32'sd25915, -32'sd2449423, -32'sd1248524, -32'sd980503, -32'sd1517927, -32'sd1190139, -32'sd2486487, -32'sd404605, 32'sd704953, 32'sd562004, 32'sd950834, 32'sd91288, 32'sd819975, 32'sd1585877, 32'sd529209, 32'sd529236, -32'sd337493, -32'sd2519789, -32'sd2075432, 32'sd99782, 32'sd930922, -32'sd667969, -32'sd2192359, -32'sd2652357, -32'sd207814, 32'sd361025, -32'sd404040, 32'sd0, 32'sd87742, -32'sd4016, -32'sd701683, -32'sd272970, -32'sd1466004, -32'sd1648516, -32'sd1017464, -32'sd3003819, -32'sd1348429, -32'sd2031242, -32'sd1032896, -32'sd377866, 32'sd1862775, 32'sd980330, -32'sd171831, 32'sd265249, 32'sd822105, 32'sd952812, -32'sd1503904, -32'sd1029038, 32'sd206349, 32'sd232393, -32'sd1673017, 32'sd788294, 32'sd1036410, 32'sd590468, -32'sd688372, -32'sd502360, -32'sd58890, -32'sd1713446, -32'sd130891, 32'sd1405754, -32'sd2392370, -32'sd1659842, -32'sd2464585, -32'sd2884812, -32'sd3957859, -32'sd563931, -32'sd420285, 32'sd1712055, -32'sd640454, 32'sd188628, 32'sd87179, 32'sd2766603, 32'sd1842860, 32'sd559277, -32'sd1782108, -32'sd2108727, 32'sd722124, -32'sd852357, -32'sd1245144, -32'sd714963, 32'sd624194, 32'sd1119506, -32'sd784392, -32'sd554596, -32'sd1183436, 32'sd1075660, -32'sd954488, 32'sd877282, -32'sd1341393, -32'sd1824281, -32'sd2896214, -32'sd2958348, -32'sd3340570, -32'sd3981853, -32'sd1875230, 32'sd7538, -32'sd1243898, 32'sd473507, 32'sd261401, -32'sd782377, 32'sd1312970, -32'sd344987, -32'sd167272, -32'sd1844860, 32'sd464100, -32'sd2253, -32'sd556777, 32'sd1696727, -32'sd98462, -32'sd559558, 32'sd381095, 32'sd0, -32'sd329469, 32'sd1620208, 32'sd1901117, -32'sd63261, -32'sd1691680, -32'sd857788, -32'sd608703, -32'sd273402, -32'sd4294855, -32'sd2551276, -32'sd1602577, -32'sd230308, -32'sd1748048, -32'sd1603856, -32'sd1034322, -32'sd1573290, -32'sd548038, -32'sd2244693, -32'sd1975804, 32'sd251660, -32'sd150050, 32'sd670686, -32'sd520493, 32'sd558266, -32'sd688742, -32'sd486847, -32'sd329939, -32'sd375923, -32'sd252229, 32'sd34126, 32'sd1543506, 32'sd959234, 32'sd84854, -32'sd959566, 32'sd781923, -32'sd492098, -32'sd1240122, 32'sd1543157, -32'sd145240, -32'sd671363, 32'sd95321, -32'sd411727, 32'sd390517, 32'sd126777, -32'sd1221798, -32'sd390051, -32'sd1719999, -32'sd2980410, 32'sd946884, -32'sd163271, -32'sd811826, -32'sd993968, -32'sd999023, 32'sd1141229, 32'sd615419, 32'sd185537, -32'sd407815, 32'sd701540, 32'sd1502192, -32'sd1169422, -32'sd77236, 32'sd944269, 32'sd588219, 32'sd390935, 32'sd510148, 32'sd1497107, 32'sd407646, 32'sd2331692, 32'sd546339, 32'sd1532121, -32'sd549725, -32'sd2960179, 32'sd930939, -32'sd1393445, -32'sd2597595, -32'sd234665, 32'sd184085, -32'sd812144, -32'sd1848661, -32'sd737003, -32'sd677202, -32'sd961813, 32'sd164685, 32'sd0, -32'sd33156, -32'sd993546, 32'sd144978, 32'sd285094, 32'sd1398871, 32'sd2465392, 32'sd618831, 32'sd174074, -32'sd286757, 32'sd1693067, 32'sd2266681, 32'sd94130, 32'sd2450776, 32'sd1074632, -32'sd726954, -32'sd2923485, -32'sd3247280, -32'sd1190134, -32'sd2421142, -32'sd1498824, -32'sd659882, 32'sd741899, 32'sd490370, 32'sd336059, 32'sd844431, -32'sd769691, 32'sd0, 32'sd0, 32'sd0, 32'sd679094, -32'sd1031910, 32'sd495729, -32'sd363233, 32'sd1248647, 32'sd232451, 32'sd1030767, 32'sd964579, 32'sd1938160, 32'sd282558, 32'sd719218, -32'sd187373, 32'sd744039, 32'sd796513, -32'sd3461240, -32'sd3933545, -32'sd2833374, -32'sd2947955, -32'sd98258, -32'sd186566, -32'sd777928, -32'sd188886, -32'sd356908, -32'sd2020373, -32'sd250603, 32'sd0, 32'sd0, 32'sd0, 32'sd924939, -32'sd48583, 32'sd516825, -32'sd495632, -32'sd2134718, 32'sd1486024, -32'sd238146, -32'sd1054079, 32'sd170283, 32'sd1595101, 32'sd1891038, 32'sd2240676, -32'sd813214, -32'sd1334976, 32'sd457092, -32'sd848705, 32'sd892104, -32'sd652401, -32'sd636642, 32'sd1409412, 32'sd823583, 32'sd847285, -32'sd934191, -32'sd698383, -32'sd395310, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd455722, -32'sd168753, -32'sd97846, 32'sd637879, -32'sd1312677, -32'sd740, 32'sd1713726, 32'sd2516646, 32'sd2595938, 32'sd836550, 32'sd2798633, 32'sd1041147, -32'sd698121, -32'sd1508362, 32'sd1133062, -32'sd18262, -32'sd517588, 32'sd78500, 32'sd1072053, -32'sd352210, -32'sd740758, 32'sd679912, -32'sd458086, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd343030, 32'sd156424, 32'sd321084, 32'sd533954, 32'sd412551, 32'sd75796, 32'sd958654, 32'sd1700926, -32'sd233091, 32'sd521786, 32'sd1820318, 32'sd1472867, 32'sd1246428, 32'sd562173, 32'sd1403072, 32'sd1558261, 32'sd2017568, -32'sd920441, -32'sd1469156, 32'sd136721, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1078878, 32'sd914671, 32'sd573895, 32'sd206360, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd100756, 32'sd792275, -32'sd61703, 32'sd466841, 32'sd1856553, -32'sd449817, 32'sd1308221, 32'sd826398, 32'sd722827, -32'sd1041321, -32'sd606090, -32'sd720104, 32'sd295567, 32'sd1071518, 32'sd236092, 32'sd428845, 32'sd594115, 32'sd480987, 32'sd672552, 32'sd1408577, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1719097, 32'sd505476, -32'sd164455, 32'sd1134127, 32'sd1468497, 32'sd1704817, -32'sd687698, -32'sd239407, 32'sd915931, 32'sd550781, 32'sd1773803, 32'sd792625, -32'sd1310664, 32'sd530865, -32'sd862593, 32'sd1176534, 32'sd1595181, 32'sd245998, 32'sd1721107, 32'sd252023, 32'sd1747837, -32'sd50328, 32'sd43722, 32'sd1440967, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1653748, 32'sd481678, -32'sd662417, 32'sd2204120, 32'sd507485, -32'sd2381917, -32'sd197095, 32'sd152286, 32'sd1246265, -32'sd609883, 32'sd1998225, 32'sd1838108, 32'sd51184, -32'sd2848129, 32'sd564637, 32'sd1701608, -32'sd507107, -32'sd652531, -32'sd484353, -32'sd208732, -32'sd384307, -32'sd596737, 32'sd314724, -32'sd1179348, 32'sd321059, 32'sd0, 32'sd0, 32'sd1243644, 32'sd1379870, -32'sd74834, 32'sd1447266, -32'sd763541, -32'sd71257, 32'sd597061, -32'sd530586, -32'sd234809, 32'sd1679135, 32'sd76243, 32'sd718458, 32'sd378610, 32'sd1694107, 32'sd1014765, -32'sd478335, 32'sd455395, 32'sd528306, 32'sd94243, 32'sd1072937, -32'sd713408, -32'sd1549697, 32'sd752333, -32'sd1254833, 32'sd776272, 32'sd845438, -32'sd596159, 32'sd0, 32'sd396793, 32'sd399397, 32'sd876063, 32'sd798650, 32'sd489681, -32'sd1560765, 32'sd183571, 32'sd724256, -32'sd900131, -32'sd37073, -32'sd70129, 32'sd1240253, 32'sd2441813, 32'sd1235421, 32'sd132410, 32'sd1343484, 32'sd1589083, -32'sd899223, -32'sd1058177, -32'sd1362701, 32'sd726891, 32'sd196798, 32'sd815633, 32'sd603651, 32'sd852740, -32'sd769009, 32'sd1492736, 32'sd0, 32'sd1185192, -32'sd317597, 32'sd592359, -32'sd165655, 32'sd1096459, -32'sd772007, -32'sd2459309, 32'sd575955, -32'sd1256230, -32'sd815953, -32'sd715031, -32'sd404217, 32'sd1982493, 32'sd527201, -32'sd88952, -32'sd317238, -32'sd1820110, -32'sd853632, -32'sd1301607, -32'sd338007, 32'sd2166334, 32'sd246862, 32'sd1603846, 32'sd475876, 32'sd13514, 32'sd549501, 32'sd32697, 32'sd1424340, 32'sd452565, 32'sd1528680, 32'sd220872, 32'sd403506, 32'sd1072140, 32'sd756497, 32'sd434757, -32'sd1741881, -32'sd547589, 32'sd612966, -32'sd382979, 32'sd952724, -32'sd503900, 32'sd709600, 32'sd1536324, 32'sd1808766, 32'sd1713390, 32'sd184978, -32'sd314958, 32'sd1941311, 32'sd2538911, 32'sd758681, -32'sd321347, 32'sd1757184, 32'sd1270112, -32'sd1051886, 32'sd906470, 32'sd1451763, -32'sd308400, 32'sd1089380, 32'sd1012055, 32'sd1102843, 32'sd1370403, 32'sd1384366, 32'sd2319972, 32'sd997305, 32'sd1029297, 32'sd438459, -32'sd943284, 32'sd592127, -32'sd10103, -32'sd164692, 32'sd2265141, 32'sd1306856, 32'sd41202, 32'sd112168, 32'sd529848, 32'sd1234989, 32'sd1610505, -32'sd889377, -32'sd1156596, 32'sd372412, 32'sd609156, 32'sd1777792, 32'sd1466535, 32'sd531223, 32'sd1505624, 32'sd1463899, 32'sd261063, -32'sd526507, 32'sd790082, 32'sd220368, 32'sd943317, -32'sd1665563, -32'sd394820, -32'sd711453, -32'sd1064160, -32'sd18024, 32'sd1300978, -32'sd2380103, -32'sd2270027, -32'sd1433929, -32'sd827722, -32'sd1087501, -32'sd299842, 32'sd1605307, 32'sd342331, -32'sd564869, -32'sd365091, 32'sd595528, 32'sd816024, 32'sd85166, -32'sd1682606, -32'sd58273, 32'sd321458, 32'sd163120, 32'sd2323564, -32'sd545272, -32'sd124704, -32'sd200518, -32'sd1989585, -32'sd1649967, -32'sd935066, 32'sd342201, 32'sd671930, 32'sd1326929, -32'sd990629, -32'sd1257350, -32'sd3362082, -32'sd2638808, -32'sd2603316, -32'sd1184239, -32'sd2006820, 32'sd243016, 32'sd2711840, -32'sd453078, 32'sd636499, 32'sd270930, 32'sd1341587, 32'sd2096665, 32'sd85898, -32'sd205805, 32'sd784770, 32'sd638865, 32'sd1084199, 32'sd496488, -32'sd820298, -32'sd147980, -32'sd234033, 32'sd757852, 32'sd993798, -32'sd409098, -32'sd391404, -32'sd1914652, -32'sd1774520, -32'sd1178459, -32'sd1628019, -32'sd929732, -32'sd2036978, -32'sd2325985, -32'sd459037, -32'sd1729360, -32'sd1456155, 32'sd1382889, 32'sd3756270, 32'sd603657, 32'sd1205946, 32'sd326752, -32'sd15317, 32'sd616715, -32'sd539357, -32'sd927748, 32'sd531492, 32'sd1215596, -32'sd503176, -32'sd196541, 32'sd978421, 32'sd2234123, -32'sd91645, -32'sd27662, 32'sd613649, 32'sd457694, -32'sd716800, 32'sd588637, -32'sd1421143, 32'sd355381, -32'sd18412, -32'sd379129, -32'sd2245064, -32'sd1684161, -32'sd1223083, 32'sd99133, 32'sd1231949, -32'sd125286, -32'sd476561, 32'sd708027, -32'sd587642, 32'sd772679, -32'sd158498, 32'sd795247, 32'sd192576, -32'sd711850, 32'sd1270967, 32'sd1154388, 32'sd1787072, 32'sd1855359, -32'sd64380, 32'sd2756093, 32'sd1615488, 32'sd1704015, 32'sd2711509, 32'sd1851209, -32'sd212379, 32'sd708081, -32'sd1767752, 32'sd721768, -32'sd2523480, 32'sd244342, -32'sd1173685, -32'sd404022, 32'sd1173655, -32'sd447470, -32'sd206376, 32'sd587570, -32'sd229402, 32'sd2469492, -32'sd588090, -32'sd243579, -32'sd1479496, 32'sd289989, 32'sd304079, 32'sd85074, 32'sd2183587, 32'sd2131895, 32'sd1044611, 32'sd2231462, 32'sd1979835, 32'sd351133, 32'sd3665047, 32'sd4115266, 32'sd2888200, 32'sd907511, -32'sd1079292, 32'sd5057, -32'sd497360, 32'sd1075223, 32'sd323838, -32'sd212864, -32'sd1921017, -32'sd1134781, -32'sd1324855, 32'sd1226916, 32'sd555064, 32'sd1874411, 32'sd555141, -32'sd998728, -32'sd1665646, -32'sd808648, 32'sd1026006, 32'sd1001725, 32'sd329703, -32'sd1240303, 32'sd790321, 32'sd1850521, 32'sd3767973, 32'sd2780592, 32'sd4447888, 32'sd3719559, 32'sd2528917, 32'sd1238421, 32'sd602587, 32'sd1698144, -32'sd1741803, -32'sd561700, 32'sd1387275, 32'sd2251441, -32'sd1688752, -32'sd2099502, -32'sd298584, 32'sd1487072, 32'sd238347, 32'sd1003369, 32'sd1231261, 32'sd1165760, -32'sd574049, 32'sd472065, -32'sd253174, -32'sd705636, -32'sd2277547, -32'sd5122579, -32'sd2311832, -32'sd878570, 32'sd846209, 32'sd3719302, 32'sd814570, 32'sd1120200, 32'sd670000, 32'sd1157159, 32'sd347471, 32'sd2816361, 32'sd468507, 32'sd522498, 32'sd188624, 32'sd1100538, -32'sd2102940, -32'sd1069732, 32'sd1866991, 32'sd2241569, 32'sd1495087, 32'sd0, 32'sd769489, -32'sd996093, -32'sd802232, -32'sd1401683, -32'sd2003901, 32'sd251031, -32'sd1638627, -32'sd2474559, -32'sd2023265, -32'sd2564408, -32'sd4008149, -32'sd2288508, -32'sd2863781, -32'sd2668571, 32'sd1730980, 32'sd2919413, 32'sd1583045, 32'sd1147312, 32'sd1847964, 32'sd1546917, 32'sd2051969, 32'sd1789743, -32'sd1463946, 32'sd1381690, -32'sd383260, 32'sd958182, 32'sd547635, 32'sd243985, 32'sd1408687, 32'sd243047, -32'sd2527176, -32'sd327232, -32'sd488541, -32'sd1575224, -32'sd2602455, -32'sd2701664, -32'sd5397722, -32'sd3166272, -32'sd4032116, -32'sd3915076, -32'sd6044921, -32'sd2397158, -32'sd873889, 32'sd344031, 32'sd2027482, -32'sd243634, 32'sd705766, 32'sd951755, 32'sd1354000, -32'sd334997, -32'sd1402905, 32'sd781568, -32'sd537675, -32'sd49655, -32'sd1073548, 32'sd738965, 32'sd515630, -32'sd675650, 32'sd471689, 32'sd656007, -32'sd1438412, -32'sd1441293, -32'sd2165898, -32'sd4612171, -32'sd2975082, -32'sd4246474, -32'sd3970651, -32'sd2286513, -32'sd4511594, -32'sd2447317, -32'sd2095401, 32'sd181942, 32'sd538821, 32'sd2213414, -32'sd1598793, 32'sd913353, 32'sd1654810, -32'sd126421, -32'sd2196466, -32'sd1192342, 32'sd1702046, 32'sd1766089, -32'sd558673, 32'sd0, -32'sd255834, 32'sd1188490, 32'sd112042, 32'sd262505, -32'sd1614980, -32'sd636120, -32'sd1051122, -32'sd1405572, -32'sd1478016, -32'sd662257, -32'sd534409, -32'sd915499, -32'sd273494, 32'sd898548, -32'sd1610162, 32'sd1251608, 32'sd2234135, 32'sd3093929, 32'sd894337, 32'sd1561098, 32'sd1335408, 32'sd539902, -32'sd2228045, -32'sd23485, -32'sd424896, -32'sd353925, 32'sd604539, 32'sd547899, 32'sd653951, 32'sd1486591, -32'sd376218, 32'sd3544379, 32'sd801895, 32'sd2303581, 32'sd1315631, 32'sd1009224, -32'sd1446615, 32'sd1934353, 32'sd1501649, 32'sd1356428, 32'sd2287444, 32'sd1704933, 32'sd174693, 32'sd652568, 32'sd79263, -32'sd361588, 32'sd556363, 32'sd2197138, -32'sd419640, -32'sd868893, -32'sd1381730, -32'sd1940981, 32'sd1420237, -32'sd1603021, 32'sd1200337, 32'sd883406, -32'sd484423, -32'sd163355, -32'sd813133, 32'sd2079633, 32'sd2263989, 32'sd916784, 32'sd2348798, 32'sd1125345, -32'sd894168, 32'sd1398499, 32'sd2303106, 32'sd2243730, 32'sd1667447, -32'sd822076, 32'sd1546685, 32'sd248308, -32'sd657692, -32'sd1705068, 32'sd493558, 32'sd631884, -32'sd436273, -32'sd3478583, -32'sd261086, -32'sd1129618, 32'sd62020, 32'sd823128, 32'sd770777, 32'sd0, 32'sd1315773, 32'sd796512, 32'sd1714929, 32'sd542588, 32'sd1231055, -32'sd2114002, -32'sd1809207, 32'sd1659663, 32'sd1033762, 32'sd3009838, 32'sd3392476, 32'sd2055374, 32'sd1998839, 32'sd147876, 32'sd141294, -32'sd200843, -32'sd1290810, -32'sd687816, 32'sd665735, 32'sd218368, -32'sd2375552, -32'sd47381, 32'sd59869, -32'sd541534, 32'sd528767, 32'sd65781, 32'sd0, 32'sd0, 32'sd0, 32'sd184566, 32'sd1550097, 32'sd147535, -32'sd137196, 32'sd440327, -32'sd1581643, -32'sd400499, 32'sd223624, 32'sd1241442, 32'sd2210639, 32'sd2079334, 32'sd880688, 32'sd400088, 32'sd1449473, 32'sd695649, 32'sd390393, -32'sd686900, -32'sd269518, -32'sd151676, -32'sd404513, -32'sd437574, -32'sd1499145, 32'sd812901, 32'sd601147, -32'sd310410, 32'sd0, 32'sd0, 32'sd0, 32'sd418770, -32'sd163617, 32'sd456319, 32'sd1114095, 32'sd1001102, -32'sd1146503, 32'sd99132, 32'sd1834453, 32'sd1875616, 32'sd1028580, 32'sd1880699, 32'sd471706, 32'sd1442628, 32'sd1079319, -32'sd1399186, -32'sd3624391, -32'sd21259, 32'sd1608356, 32'sd445854, 32'sd285229, 32'sd1713720, 32'sd1421797, 32'sd540437, 32'sd1536469, 32'sd630896, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd612032, 32'sd561303, 32'sd1145960, 32'sd897054, -32'sd519761, 32'sd44841, 32'sd867461, 32'sd711645, 32'sd268105, -32'sd727929, 32'sd443488, 32'sd1723037, 32'sd530675, 32'sd891436, -32'sd1148951, -32'sd821050, 32'sd202626, 32'sd451247, 32'sd1155487, 32'sd1208698, 32'sd1425771, 32'sd1827441, 32'sd466913, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1770955, 32'sd1217651, -32'sd199763, 32'sd812818, 32'sd221455, 32'sd572833, -32'sd647490, -32'sd46784, 32'sd368313, 32'sd1572555, 32'sd941504, -32'sd144598, -32'sd1099174, 32'sd1271755, 32'sd1011948, -32'sd492063, -32'sd577159, -32'sd699353, -32'sd1843688, -32'sd198204, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd405951, 32'sd1910791, -32'sd426935, 32'sd749284, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd300935, 32'sd314832, 32'sd1063898, 32'sd418366, 32'sd1301204, 32'sd474241, 32'sd573195, 32'sd1405982, 32'sd1650533, 32'sd949699, 32'sd1330248, 32'sd112415, 32'sd1083648, 32'sd1314660, 32'sd499791, -32'sd49812, 32'sd946303, 32'sd1686831, 32'sd178430, 32'sd960467, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd186506, -32'sd788960, 32'sd71162, -32'sd1309585, 32'sd572265, 32'sd1445678, -32'sd1526243, -32'sd1642774, 32'sd474814, -32'sd1019371, -32'sd1020684, -32'sd680633, 32'sd1209569, 32'sd771526, 32'sd1969910, 32'sd2343056, 32'sd135247, 32'sd156862, -32'sd548807, -32'sd1628549, 32'sd242848, 32'sd116860, 32'sd296536, 32'sd947861, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd341976, 32'sd1430851, 32'sd1266266, -32'sd1750892, -32'sd369401, -32'sd488844, -32'sd3717133, -32'sd2190875, -32'sd1635721, 32'sd655256, 32'sd66312, 32'sd1399364, 32'sd2309911, 32'sd1327622, 32'sd1752903, 32'sd958301, 32'sd214032, -32'sd1284875, -32'sd1905071, -32'sd1877008, 32'sd37866, -32'sd54157, -32'sd494033, -32'sd956605, 32'sd1599829, 32'sd0, 32'sd0, 32'sd517104, 32'sd799067, -32'sd1144659, -32'sd454830, -32'sd965350, -32'sd217781, -32'sd370479, -32'sd741943, 32'sd1507922, -32'sd939065, -32'sd2233707, -32'sd1236440, 32'sd2516778, 32'sd1504776, 32'sd968093, 32'sd1465715, 32'sd2715116, 32'sd1388421, 32'sd1874450, -32'sd368018, -32'sd2606950, -32'sd1289601, -32'sd1656928, -32'sd786301, -32'sd123032, 32'sd591140, 32'sd877544, 32'sd0, 32'sd379195, -32'sd850548, 32'sd1152325, -32'sd1394684, 32'sd1568074, -32'sd75585, -32'sd70556, 32'sd1396275, 32'sd1623548, 32'sd186331, 32'sd544385, -32'sd1075704, -32'sd2129419, -32'sd2917231, -32'sd795457, 32'sd59339, 32'sd99089, 32'sd1678600, 32'sd1521564, 32'sd1444343, -32'sd666310, -32'sd1562241, 32'sd1837846, 32'sd712772, 32'sd917907, -32'sd184742, -32'sd1105082, 32'sd0, 32'sd271346, 32'sd81911, 32'sd672854, 32'sd342931, 32'sd897084, 32'sd139283, -32'sd405601, 32'sd1736434, 32'sd1560957, -32'sd1951524, -32'sd1676328, 32'sd178984, -32'sd1505502, -32'sd1803168, -32'sd2534410, -32'sd3305944, 32'sd1167094, 32'sd2736227, 32'sd2302288, 32'sd1051854, 32'sd1494936, 32'sd539762, 32'sd244749, 32'sd670306, 32'sd874432, -32'sd1031574, 32'sd755708, 32'sd194478, 32'sd423803, 32'sd1507937, 32'sd1255579, 32'sd1982158, 32'sd1551829, 32'sd290129, 32'sd455995, 32'sd1153502, -32'sd11640, -32'sd956981, 32'sd1143014, 32'sd2221739, -32'sd758851, -32'sd2519871, -32'sd3060132, -32'sd2920420, -32'sd1284898, 32'sd1672648, 32'sd2595576, 32'sd368309, -32'sd168038, 32'sd1048461, -32'sd1164068, -32'sd585413, -32'sd809531, -32'sd1561910, -32'sd1393552, 32'sd233716, 32'sd535419, 32'sd913786, 32'sd1262810, 32'sd547518, 32'sd1291311, 32'sd150316, 32'sd1724131, -32'sd473419, 32'sd1213793, 32'sd1072659, 32'sd1710934, 32'sd964487, -32'sd1070100, -32'sd4028435, -32'sd5199862, -32'sd3030330, 32'sd1736178, 32'sd4424881, 32'sd2618330, 32'sd664107, 32'sd1267184, -32'sd56835, -32'sd267712, -32'sd2966555, -32'sd1717039, -32'sd1032116, 32'sd24269, -32'sd725351, 32'sd594003, -32'sd586857, 32'sd89450, 32'sd2458801, -32'sd87233, -32'sd1036297, 32'sd1908062, 32'sd1871358, 32'sd278795, 32'sd148374, 32'sd1793115, 32'sd1094351, -32'sd1094036, -32'sd2178248, -32'sd5629066, -32'sd3094731, 32'sd2840485, 32'sd4771067, 32'sd2970133, 32'sd2771282, 32'sd1039640, -32'sd1948833, -32'sd1130363, -32'sd1832604, 32'sd118521, -32'sd821235, 32'sd894643, 32'sd884454, -32'sd778517, 32'sd1342053, 32'sd1686133, 32'sd313459, -32'sd955673, -32'sd871721, 32'sd1213372, 32'sd542780, 32'sd59312, 32'sd833987, 32'sd537963, -32'sd842749, -32'sd2983625, -32'sd2282177, -32'sd2117873, 32'sd93091, 32'sd2765991, 32'sd3265653, 32'sd1892163, 32'sd890678, 32'sd1189853, -32'sd1595164, -32'sd2682353, -32'sd2624287, -32'sd226297, -32'sd1362764, -32'sd101364, -32'sd569977, 32'sd915044, 32'sd712787, 32'sd1127596, 32'sd430298, -32'sd1253675, -32'sd412349, 32'sd733482, 32'sd2227448, -32'sd1358629, 32'sd1472132, 32'sd65791, -32'sd520353, -32'sd847333, -32'sd1408632, 32'sd320739, 32'sd462089, 32'sd2749784, 32'sd2640194, -32'sd1522347, 32'sd988598, -32'sd886446, -32'sd694074, -32'sd1372388, 32'sd498810, -32'sd45604, -32'sd516971, 32'sd20280, 32'sd222051, 32'sd1086217, -32'sd1115837, -32'sd536372, -32'sd904084, 32'sd1663820, -32'sd12906, 32'sd86810, -32'sd982584, 32'sd1650197, 32'sd1117613, 32'sd915491, -32'sd692708, -32'sd276566, 32'sd157715, -32'sd1768232, 32'sd1946596, 32'sd1594636, 32'sd176656, -32'sd296892, -32'sd802795, -32'sd1321296, -32'sd339129, -32'sd1113037, 32'sd1916600, -32'sd1123570, -32'sd1179184, 32'sd483625, -32'sd139862, -32'sd186265, 32'sd1252209, 32'sd369936, -32'sd1118589, 32'sd109767, 32'sd580748, 32'sd687112, 32'sd728804, 32'sd1429577, -32'sd877652, 32'sd1301881, -32'sd1789723, -32'sd1519114, -32'sd439536, -32'sd360902, 32'sd68982, 32'sd2133499, 32'sd668478, -32'sd1263505, 32'sd606713, 32'sd160948, -32'sd14743, -32'sd1355596, -32'sd1610193, -32'sd1292050, -32'sd130955, 32'sd493221, -32'sd682316, 32'sd961386, -32'sd689155, -32'sd2370517, 32'sd1014105, 32'sd1329774, 32'sd369227, -32'sd1302976, -32'sd835385, 32'sd2166230, 32'sd1843680, 32'sd969606, 32'sd287954, 32'sd490126, 32'sd883125, -32'sd597746, -32'sd1984634, 32'sd654072, 32'sd832966, -32'sd39558, 32'sd38372, 32'sd1507958, 32'sd1487408, -32'sd538761, 32'sd640278, -32'sd47750, 32'sd616793, 32'sd1176837, -32'sd252591, 32'sd393185, 32'sd73714, 32'sd1288344, 32'sd430592, -32'sd1847641, -32'sd1159334, 32'sd276200, 32'sd2393982, 32'sd1559408, 32'sd2204698, 32'sd686093, -32'sd909301, 32'sd1675536, 32'sd1467115, -32'sd339748, -32'sd1620034, -32'sd1229176, 32'sd229581, 32'sd2094046, -32'sd587190, -32'sd158680, 32'sd677231, -32'sd1718490, 32'sd1561609, -32'sd1277287, -32'sd2010371, 32'sd28335, 32'sd130160, -32'sd508316, 32'sd99419, -32'sd875848, -32'sd144588, -32'sd1836744, -32'sd2919775, 32'sd702271, 32'sd1669390, 32'sd1999116, 32'sd1204825, 32'sd310128, -32'sd901586, 32'sd1310204, 32'sd2258875, 32'sd353767, 32'sd31348, -32'sd1619306, -32'sd1114001, 32'sd1228734, -32'sd929303, 32'sd20328, -32'sd774492, -32'sd920727, -32'sd395451, -32'sd837246, -32'sd529856, 32'sd378962, 32'sd0, 32'sd654766, 32'sd411028, 32'sd1194463, -32'sd75602, -32'sd729626, -32'sd1190760, 32'sd2808295, 32'sd2169837, 32'sd369466, 32'sd582549, -32'sd994687, 32'sd125668, 32'sd166922, 32'sd1491294, 32'sd748274, -32'sd922851, 32'sd697299, 32'sd516151, -32'sd586029, -32'sd1167119, -32'sd1051758, 32'sd174152, -32'sd1707216, -32'sd1242199, -32'sd1257456, -32'sd823712, 32'sd1601803, -32'sd129420, 32'sd934469, 32'sd553022, 32'sd2037645, -32'sd104410, -32'sd745380, -32'sd982016, 32'sd2324218, 32'sd2286012, 32'sd886789, 32'sd347650, -32'sd1021276, -32'sd2888221, -32'sd2112632, -32'sd753683, 32'sd213637, -32'sd146493, -32'sd1137781, 32'sd1260903, 32'sd249178, 32'sd557497, 32'sd80041, -32'sd622485, -32'sd2851059, -32'sd805175, 32'sd1385064, -32'sd1247016, -32'sd60568, 32'sd362654, -32'sd474966, -32'sd876058, 32'sd2393542, -32'sd1250810, -32'sd586490, -32'sd2125649, 32'sd1093960, 32'sd316939, 32'sd552110, 32'sd2416531, 32'sd680942, -32'sd4196184, -32'sd1684928, -32'sd476588, 32'sd2320173, 32'sd1884210, 32'sd111831, -32'sd1134977, -32'sd874987, -32'sd1052083, -32'sd866134, -32'sd465520, -32'sd1631666, -32'sd762949, -32'sd304598, -32'sd1803800, -32'sd269380, 32'sd0, 32'sd772164, 32'sd502240, 32'sd1171074, 32'sd330514, -32'sd46112, -32'sd877133, -32'sd431999, 32'sd1411618, 32'sd561392, 32'sd1759188, -32'sd449662, -32'sd1097070, -32'sd836173, -32'sd1321831, 32'sd1637376, 32'sd194436, -32'sd1063328, -32'sd544650, 32'sd383280, 32'sd964503, 32'sd827975, -32'sd1948152, 32'sd772606, -32'sd349224, -32'sd422087, 32'sd937597, -32'sd685061, -32'sd349267, 32'sd731610, 32'sd1502045, 32'sd857410, -32'sd254656, -32'sd843392, 32'sd594460, 32'sd436563, 32'sd623089, 32'sd1649626, 32'sd1070914, -32'sd554385, 32'sd137423, 32'sd451797, 32'sd104546, 32'sd1669639, -32'sd289096, -32'sd308256, -32'sd889808, -32'sd142028, 32'sd214541, 32'sd558966, 32'sd499179, 32'sd627524, -32'sd1270812, 32'sd1195565, 32'sd1596153, 32'sd466830, -32'sd78735, -32'sd1026023, 32'sd653940, 32'sd1104505, 32'sd719719, 32'sd226024, 32'sd262430, -32'sd75766, 32'sd2351840, 32'sd764668, 32'sd274781, 32'sd562384, 32'sd977476, 32'sd1088027, -32'sd807769, 32'sd1496270, 32'sd661983, -32'sd626085, -32'sd490084, 32'sd144356, 32'sd65538, -32'sd257873, -32'sd1645589, -32'sd2056728, -32'sd175681, -32'sd60915, 32'sd110015, -32'sd303552, 32'sd0, -32'sd43624, 32'sd538055, 32'sd874185, 32'sd538581, 32'sd1214153, 32'sd1150284, 32'sd1640295, 32'sd2670741, -32'sd62210, -32'sd323282, 32'sd996198, -32'sd1103424, -32'sd1877594, -32'sd376012, -32'sd102635, -32'sd487578, -32'sd1832517, -32'sd125851, -32'sd337278, -32'sd856560, 32'sd732607, -32'sd659268, 32'sd1207046, 32'sd834087, -32'sd1615592, 32'sd375159, 32'sd0, 32'sd0, 32'sd0, 32'sd434415, -32'sd573539, 32'sd1287344, 32'sd1644987, -32'sd1377394, -32'sd308129, -32'sd594843, 32'sd164084, 32'sd592223, 32'sd662032, -32'sd1494256, -32'sd1189438, -32'sd532448, -32'sd1734004, -32'sd502400, -32'sd855838, -32'sd1317814, 32'sd746518, 32'sd1132124, 32'sd617066, -32'sd961193, -32'sd778277, -32'sd1240451, -32'sd203341, 32'sd756441, 32'sd0, 32'sd0, 32'sd0, -32'sd307287, 32'sd950399, -32'sd62115, -32'sd83021, -32'sd1117558, -32'sd1643949, -32'sd541362, 32'sd141452, 32'sd749025, -32'sd793528, -32'sd2094366, -32'sd1469604, -32'sd2178836, -32'sd1748162, -32'sd912142, 32'sd502235, 32'sd288659, -32'sd2315801, -32'sd343751, -32'sd718970, -32'sd981137, 32'sd1358076, -32'sd443564, -32'sd162129, -32'sd285219, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd384846, 32'sd57348, -32'sd1735083, 32'sd856997, -32'sd4384, 32'sd1910197, 32'sd878250, -32'sd719273, -32'sd2579582, 32'sd1590774, -32'sd26801, -32'sd1170065, -32'sd955586, -32'sd563797, 32'sd2227960, -32'sd977839, -32'sd2181708, -32'sd1507090, -32'sd2379596, -32'sd2329929, 32'sd921040, 32'sd1343977, 32'sd744164, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd908721, 32'sd543860, 32'sd629200, -32'sd811061, -32'sd405446, 32'sd255947, -32'sd684905, -32'sd733081, 32'sd918387, -32'sd268044, -32'sd820430, 32'sd273176, -32'sd758495, -32'sd120627, -32'sd49423, 32'sd325639, 32'sd1077126, -32'sd210048, -32'sd417877, -32'sd188947, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd198910, -32'sd196652, -32'sd304937, 32'sd38511, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd531534, 32'sd1076875, -32'sd1060786, 32'sd455995, 32'sd889780, -32'sd1013357, 32'sd1428580, 32'sd258498, 32'sd245846, -32'sd981312, 32'sd1253573, 32'sd383230, -32'sd1041635, 32'sd1047603, 32'sd345738, 32'sd69105, 32'sd1155272, 32'sd1421948, 32'sd989201, 32'sd1022581, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1442975, 32'sd1482895, 32'sd546808, 32'sd170440, 32'sd72443, -32'sd948121, -32'sd218601, -32'sd354071, 32'sd1757536, 32'sd647998, 32'sd133481, -32'sd328305, -32'sd2994082, -32'sd2879495, -32'sd1980951, 32'sd870788, 32'sd465929, 32'sd1311663, -32'sd300928, 32'sd70910, 32'sd1614340, -32'sd76820, 32'sd334805, 32'sd227990, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1864336, 32'sd1778655, -32'sd604464, 32'sd1384091, 32'sd254531, 32'sd1320515, 32'sd957310, -32'sd2089781, -32'sd805284, -32'sd735275, 32'sd511844, -32'sd2248829, -32'sd1759955, -32'sd602053, -32'sd1314015, 32'sd552639, -32'sd2054315, 32'sd798008, -32'sd293607, -32'sd553521, 32'sd216807, -32'sd669450, -32'sd314666, -32'sd1159953, -32'sd258485, 32'sd0, 32'sd0, 32'sd337182, 32'sd273021, 32'sd658374, -32'sd1025605, 32'sd528658, -32'sd1539025, 32'sd267804, -32'sd481139, -32'sd1505136, -32'sd1220684, -32'sd449614, -32'sd1617460, -32'sd2414010, -32'sd699693, -32'sd1155991, 32'sd486293, -32'sd577270, 32'sd39226, -32'sd588891, -32'sd609714, 32'sd953431, -32'sd211799, -32'sd1217852, -32'sd715338, 32'sd1145531, 32'sd1015751, -32'sd845821, 32'sd0, 32'sd936097, 32'sd836473, -32'sd1674251, -32'sd1124954, 32'sd555402, -32'sd364666, -32'sd418856, 32'sd704033, 32'sd59306, -32'sd563654, -32'sd2393271, -32'sd1205750, -32'sd1425558, 32'sd980145, 32'sd974919, 32'sd1132938, 32'sd95408, -32'sd1940041, -32'sd2619041, -32'sd612640, -32'sd1460983, 32'sd285526, 32'sd2351702, -32'sd34329, 32'sd427156, 32'sd933301, -32'sd20737, 32'sd0, 32'sd375557, 32'sd990891, 32'sd754888, 32'sd1168625, 32'sd82957, -32'sd286459, -32'sd834247, 32'sd1269473, -32'sd504283, 32'sd1866935, 32'sd1149318, -32'sd1457976, -32'sd2093011, -32'sd978136, -32'sd988918, -32'sd606571, -32'sd1598853, -32'sd33171, 32'sd908454, 32'sd743082, -32'sd266146, 32'sd4421, 32'sd1306844, 32'sd1889481, -32'sd953130, -32'sd157355, 32'sd1305954, 32'sd500128, 32'sd245116, 32'sd221464, 32'sd406258, -32'sd5010, -32'sd180967, -32'sd609477, 32'sd506881, -32'sd583483, 32'sd1756275, 32'sd848605, 32'sd739037, -32'sd1594219, -32'sd2206719, -32'sd239308, 32'sd774740, 32'sd476705, 32'sd1920787, -32'sd1071682, 32'sd1700044, 32'sd3005354, 32'sd491289, 32'sd2553592, 32'sd235101, 32'sd445064, -32'sd717839, -32'sd722425, -32'sd926661, 32'sd889411, 32'sd384125, -32'sd1179379, -32'sd118056, -32'sd1662087, -32'sd24172, -32'sd194980, -32'sd228328, -32'sd324228, 32'sd1003114, -32'sd792096, -32'sd1799941, 32'sd218869, 32'sd1367626, 32'sd242092, 32'sd788348, 32'sd1399812, 32'sd1960549, 32'sd2521033, 32'sd2596058, 32'sd1529987, 32'sd1611474, 32'sd919108, 32'sd1577406, 32'sd1629394, 32'sd574754, 32'sd253467, 32'sd681579, 32'sd1787672, -32'sd274998, 32'sd1342962, -32'sd1484138, -32'sd438625, -32'sd1096033, -32'sd932852, -32'sd654597, -32'sd1379856, -32'sd681669, -32'sd395354, 32'sd600378, -32'sd974069, -32'sd747492, -32'sd2545360, -32'sd2135615, 32'sd1866162, 32'sd228410, 32'sd2805623, -32'sd903123, 32'sd475495, 32'sd926474, 32'sd891903, 32'sd568307, 32'sd2276017, 32'sd1193298, 32'sd440186, -32'sd637587, 32'sd560431, 32'sd999115, 32'sd1626757, 32'sd1795301, 32'sd203340, 32'sd143343, -32'sd851559, -32'sd2184274, -32'sd926625, 32'sd750698, -32'sd102699, -32'sd1676494, -32'sd2394841, -32'sd2643361, -32'sd3215681, -32'sd941551, -32'sd968391, -32'sd615990, -32'sd1470711, -32'sd3224251, 32'sd101296, 32'sd683188, 32'sd2143352, 32'sd423628, 32'sd828547, 32'sd1522226, 32'sd945150, -32'sd257676, 32'sd1540238, 32'sd397316, 32'sd267484, -32'sd880947, -32'sd1615610, 32'sd1680629, 32'sd212284, -32'sd1294477, -32'sd1542011, -32'sd398619, -32'sd580259, -32'sd1021642, -32'sd3429132, -32'sd2525520, 32'sd163502, -32'sd1946910, -32'sd3305932, -32'sd2502190, -32'sd2661418, -32'sd4069231, -32'sd1678524, -32'sd914501, -32'sd2179033, -32'sd951751, -32'sd307303, 32'sd378806, -32'sd648512, 32'sd926484, 32'sd420714, 32'sd238246, -32'sd331439, -32'sd1268232, -32'sd717263, -32'sd281728, -32'sd700326, -32'sd500794, -32'sd1652286, -32'sd633267, -32'sd903071, -32'sd499403, -32'sd1651191, -32'sd593571, 32'sd2237037, -32'sd752479, -32'sd3086944, -32'sd3570978, -32'sd1254250, -32'sd3423299, -32'sd2412006, -32'sd2327272, -32'sd241788, 32'sd562836, -32'sd957247, -32'sd3218831, -32'sd2445213, 32'sd680832, 32'sd658931, 32'sd514380, -32'sd430591, -32'sd1369174, -32'sd394843, 32'sd485045, 32'sd574620, 32'sd128799, -32'sd1306038, 32'sd997960, -32'sd478202, -32'sd1436346, -32'sd227877, -32'sd1467665, 32'sd1836391, -32'sd307125, -32'sd1337460, -32'sd2100096, -32'sd1183881, -32'sd2524215, -32'sd1759581, -32'sd1375179, -32'sd1305018, 32'sd1562165, -32'sd400963, 32'sd409423, -32'sd2578460, 32'sd334922, 32'sd1188009, -32'sd239761, -32'sd626783, -32'sd72818, 32'sd2172336, -32'sd1190079, -32'sd1214632, 32'sd879500, 32'sd2018912, 32'sd589155, -32'sd450956, -32'sd1670080, -32'sd2584711, -32'sd1462392, 32'sd1567722, -32'sd682839, -32'sd1653995, -32'sd1057773, -32'sd1217183, -32'sd2592572, -32'sd1930287, -32'sd1577934, 32'sd169297, 32'sd2634690, 32'sd3966969, -32'sd204188, -32'sd1367505, 32'sd170296, 32'sd2208697, 32'sd145487, -32'sd1880987, -32'sd1013724, 32'sd1229266, -32'sd568871, -32'sd76655, 32'sd840148, 32'sd388192, 32'sd2284875, 32'sd100449, -32'sd44904, -32'sd652, 32'sd497927, -32'sd856955, -32'sd792096, -32'sd1055270, -32'sd935747, -32'sd1699089, -32'sd3437152, -32'sd3109953, -32'sd870353, -32'sd1107637, 32'sd1585359, 32'sd2946228, -32'sd1232057, -32'sd2000028, 32'sd465586, 32'sd440511, -32'sd484645, -32'sd573629, -32'sd1743138, -32'sd1143502, -32'sd111226, -32'sd1391215, -32'sd1181864, -32'sd1626985, 32'sd596145, 32'sd1764776, 32'sd548901, 32'sd583303, 32'sd1964580, 32'sd443262, -32'sd1211099, -32'sd2013010, -32'sd1719935, -32'sd469597, 32'sd234207, -32'sd3217922, 32'sd715261, 32'sd1575229, 32'sd1376685, 32'sd3254937, 32'sd755611, -32'sd1217634, 32'sd1218904, 32'sd0, -32'sd238138, -32'sd351545, -32'sd1456730, -32'sd628793, -32'sd1095577, -32'sd1217964, -32'sd1768514, -32'sd607069, -32'sd1326609, -32'sd2582454, -32'sd559096, -32'sd1521250, -32'sd50550, -32'sd2509489, -32'sd2713965, -32'sd1723730, -32'sd938976, -32'sd999275, 32'sd420094, 32'sd1685226, 32'sd726509, 32'sd1686975, 32'sd2281718, 32'sd2795852, -32'sd87959, 32'sd1105229, -32'sd865174, 32'sd441580, -32'sd275031, 32'sd95441, 32'sd42409, 32'sd825268, 32'sd102170, -32'sd2758512, -32'sd2477356, -32'sd1509500, -32'sd4018278, -32'sd2305561, -32'sd2415985, -32'sd1689839, -32'sd11452, -32'sd3517467, -32'sd4763553, -32'sd262460, -32'sd938846, -32'sd297284, 32'sd345396, 32'sd1517245, -32'sd831971, 32'sd416347, 32'sd394277, -32'sd1461066, 32'sd810082, 32'sd784636, -32'sd944303, 32'sd944743, 32'sd778688, -32'sd1111679, 32'sd269234, -32'sd1681548, -32'sd286943, -32'sd919194, -32'sd1504450, -32'sd2395279, -32'sd3117938, -32'sd4019807, -32'sd4356521, -32'sd3659134, -32'sd720514, -32'sd1232351, -32'sd2971297, -32'sd1817909, -32'sd1129561, 32'sd1178908, 32'sd1110052, 32'sd2870047, -32'sd574890, -32'sd531587, 32'sd981679, 32'sd661717, -32'sd58671, 32'sd966494, -32'sd726549, 32'sd0, 32'sd311802, -32'sd131810, -32'sd952107, 32'sd1301217, 32'sd123406, 32'sd47221, -32'sd1137093, -32'sd58064, -32'sd2101906, -32'sd2068059, -32'sd3372989, -32'sd3151832, -32'sd1219317, -32'sd1050242, -32'sd2317358, 32'sd318307, 32'sd777661, 32'sd438181, 32'sd2112138, 32'sd2297695, -32'sd80385, -32'sd227173, 32'sd161622, 32'sd2246205, -32'sd488133, 32'sd550438, 32'sd1239090, 32'sd706000, 32'sd960151, 32'sd1352680, 32'sd168108, 32'sd890200, 32'sd1059095, -32'sd1011381, 32'sd403414, 32'sd2011124, 32'sd1075407, -32'sd1628282, 32'sd1945923, -32'sd76239, 32'sd318523, -32'sd291060, 32'sd1103697, 32'sd1379867, -32'sd1358167, 32'sd1865753, 32'sd640219, 32'sd1024719, -32'sd436934, 32'sd352111, -32'sd241495, 32'sd599597, -32'sd1864576, 32'sd1231774, 32'sd380237, 32'sd1543516, 32'sd1119068, 32'sd1280298, 32'sd1500939, -32'sd707737, 32'sd2338376, 32'sd1372311, 32'sd839610, 32'sd654141, 32'sd101507, 32'sd813109, 32'sd2176862, -32'sd792280, 32'sd856981, -32'sd563365, 32'sd213078, -32'sd431534, 32'sd883486, 32'sd546359, 32'sd1478438, 32'sd1778984, 32'sd218609, 32'sd554008, 32'sd302612, -32'sd2033938, -32'sd2493238, -32'sd359124, 32'sd1084944, 32'sd0, 32'sd475428, -32'sd1091137, -32'sd29970, 32'sd198661, 32'sd1429432, -32'sd461489, 32'sd484349, -32'sd766520, 32'sd2065486, 32'sd1305800, 32'sd307727, -32'sd727139, -32'sd322968, 32'sd760067, 32'sd890108, 32'sd2608627, 32'sd1358560, -32'sd2350614, -32'sd2170411, -32'sd1025945, 32'sd338616, 32'sd513519, -32'sd1030992, -32'sd345342, 32'sd593258, -32'sd1392471, 32'sd0, 32'sd0, 32'sd0, -32'sd181068, 32'sd673172, 32'sd365842, 32'sd321108, 32'sd398519, -32'sd16860, -32'sd277142, 32'sd701938, -32'sd1197676, -32'sd262838, -32'sd960327, 32'sd13473, 32'sd435962, 32'sd337834, -32'sd889673, 32'sd1447579, -32'sd703581, -32'sd2682202, -32'sd817988, 32'sd744375, -32'sd1003896, -32'sd1734486, 32'sd17969, 32'sd1202004, 32'sd167414, 32'sd0, 32'sd0, 32'sd0, 32'sd964777, -32'sd332335, 32'sd556224, -32'sd642815, -32'sd649952, 32'sd56093, 32'sd1479966, 32'sd523125, -32'sd221721, -32'sd165390, 32'sd139666, 32'sd919796, 32'sd719115, 32'sd1216856, -32'sd771188, -32'sd506408, 32'sd314443, 32'sd1098106, 32'sd970945, 32'sd664325, 32'sd97374, -32'sd2504984, -32'sd220807, 32'sd549690, 32'sd472095, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1376507, -32'sd1214871, -32'sd297748, -32'sd979627, -32'sd357391, -32'sd2284420, -32'sd907814, 32'sd334911, 32'sd659283, -32'sd1301281, -32'sd774127, -32'sd138320, -32'sd28823, -32'sd1875324, 32'sd485838, 32'sd861818, 32'sd418299, -32'sd980909, 32'sd457977, -32'sd1855264, -32'sd88486, 32'sd436813, 32'sd913929, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1537478, 32'sd1183412, 32'sd527150, 32'sd219210, -32'sd29631, 32'sd399064, 32'sd132080, 32'sd908723, 32'sd886824, 32'sd2390, -32'sd1268668, 32'sd964331, -32'sd77668, -32'sd281631, 32'sd128749, -32'sd691833, 32'sd483379, -32'sd420513, -32'sd1723799, 32'sd1237016, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd169833, -32'sd1199568, -32'sd234296, -32'sd385996, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd799526, 32'sd1074801, 32'sd639485, 32'sd180031, 32'sd1648275, 32'sd1098076, -32'sd539690, 32'sd1380239, 32'sd375283, -32'sd642472, 32'sd554836, 32'sd1357209, 32'sd422534, -32'sd183002, 32'sd952197, 32'sd400198, 32'sd1153999, 32'sd1109231, -32'sd423870, 32'sd338706, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd182117, -32'sd252889, 32'sd191857, -32'sd259847, 32'sd424127, 32'sd123785, -32'sd673231, -32'sd1720403, 32'sd130868, -32'sd711063, 32'sd816042, 32'sd237226, 32'sd634764, -32'sd816521, -32'sd2082522, -32'sd473524, 32'sd175041, 32'sd385552, -32'sd967059, 32'sd2091487, -32'sd194260, 32'sd1667548, 32'sd506871, -32'sd294612, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd350207, -32'sd685268, -32'sd1408549, 32'sd307042, -32'sd378349, -32'sd1917039, 32'sd1088196, -32'sd69619, -32'sd1088866, 32'sd163139, -32'sd532589, 32'sd885854, -32'sd353500, -32'sd291603, 32'sd68699, -32'sd2125813, -32'sd2742259, -32'sd2060784, -32'sd3190407, -32'sd671762, -32'sd983646, 32'sd1095109, -32'sd522183, -32'sd79428, -32'sd164082, 32'sd0, 32'sd0, 32'sd137643, -32'sd28367, -32'sd1399913, 32'sd446509, -32'sd815306, 32'sd362123, -32'sd92473, -32'sd879263, -32'sd1020416, 32'sd1442148, -32'sd81368, 32'sd1840946, 32'sd2033069, 32'sd2010817, -32'sd679598, -32'sd1345751, -32'sd1345095, -32'sd833528, 32'sd435556, 32'sd1908962, -32'sd753914, 32'sd59409, -32'sd2030842, 32'sd754818, 32'sd468228, 32'sd957630, -32'sd194963, 32'sd0, -32'sd356934, 32'sd716727, -32'sd618752, 32'sd356474, 32'sd214484, 32'sd1151261, 32'sd981538, 32'sd230540, -32'sd1383174, -32'sd196544, -32'sd1287695, 32'sd1798948, 32'sd1202498, -32'sd1728282, -32'sd148899, 32'sd109973, -32'sd981904, -32'sd1387263, -32'sd931884, -32'sd2021860, -32'sd973921, -32'sd13894, 32'sd577461, -32'sd1762013, -32'sd629837, 32'sd52550, -32'sd93003, 32'sd0, 32'sd545927, -32'sd35328, -32'sd2085030, -32'sd20684, -32'sd894967, 32'sd530411, 32'sd1420161, 32'sd223667, -32'sd1030910, -32'sd1558980, -32'sd959372, -32'sd949303, -32'sd907006, 32'sd733334, 32'sd923368, 32'sd893849, -32'sd776082, -32'sd366655, -32'sd123267, 32'sd145386, 32'sd222546, 32'sd572478, -32'sd1283823, -32'sd2864328, -32'sd2486426, 32'sd1727144, -32'sd28692, 32'sd351191, 32'sd267844, -32'sd1463035, 32'sd1226504, 32'sd314183, -32'sd1070198, -32'sd232278, -32'sd1300265, -32'sd462573, -32'sd1457958, -32'sd1805784, -32'sd349876, -32'sd1549451, -32'sd927599, 32'sd1119437, 32'sd2613767, 32'sd702472, -32'sd352724, -32'sd459516, -32'sd1895668, -32'sd1290977, 32'sd702948, -32'sd198381, -32'sd1510497, -32'sd2838460, -32'sd2195596, -32'sd640498, -32'sd371328, -32'sd352310, 32'sd942674, -32'sd573428, -32'sd1221529, 32'sd1484639, -32'sd1432682, -32'sd995718, -32'sd915117, -32'sd1016797, -32'sd1347355, -32'sd2179052, -32'sd1489974, -32'sd1202009, -32'sd2160979, -32'sd544913, -32'sd1048871, -32'sd1858457, -32'sd604928, 32'sd1046982, -32'sd734154, -32'sd550034, 32'sd1050665, -32'sd774237, -32'sd2830169, -32'sd3180459, -32'sd600259, 32'sd656296, -32'sd35770, 32'sd1579995, -32'sd256208, -32'sd1626802, -32'sd206222, -32'sd880297, -32'sd2797455, -32'sd1144207, -32'sd1187112, -32'sd257498, 32'sd211856, 32'sd713413, -32'sd355434, -32'sd1379845, -32'sd1012346, -32'sd1530394, -32'sd844602, 32'sd1213744, 32'sd1867803, -32'sd1718946, -32'sd417390, -32'sd1072493, -32'sd193301, -32'sd2164579, 32'sd17073, 32'sd667058, -32'sd904655, -32'sd828146, -32'sd413020, -32'sd218852, -32'sd21977, -32'sd537232, 32'sd300254, -32'sd403582, -32'sd3101365, -32'sd3845177, 32'sd129135, -32'sd283661, 32'sd2248095, 32'sd1094166, 32'sd755866, 32'sd511913, -32'sd1719492, 32'sd574028, -32'sd2858626, -32'sd772962, 32'sd1113208, 32'sd1887405, -32'sd229533, -32'sd2172522, -32'sd3983522, -32'sd1458972, -32'sd2226234, -32'sd155947, -32'sd2949368, -32'sd701242, -32'sd280368, 32'sd650929, 32'sd1224627, 32'sd549313, -32'sd842729, -32'sd1491256, -32'sd2640148, -32'sd2244495, 32'sd1086516, 32'sd1494115, 32'sd792744, 32'sd471189, 32'sd1705748, -32'sd448926, 32'sd1134374, 32'sd235560, -32'sd2990058, -32'sd594269, 32'sd1788674, 32'sd3287252, 32'sd1738552, 32'sd9424, -32'sd1130653, -32'sd1210398, -32'sd1854350, -32'sd2823402, -32'sd475367, 32'sd84816, 32'sd1258352, -32'sd337682, -32'sd1614936, -32'sd325743, -32'sd1315604, 32'sd68439, -32'sd1019375, -32'sd1784944, -32'sd700832, 32'sd883309, 32'sd1561545, -32'sd856464, 32'sd100084, -32'sd2307700, -32'sd1776191, -32'sd209507, 32'sd119662, 32'sd1369502, 32'sd1610412, 32'sd3198804, 32'sd1017067, 32'sd677896, -32'sd632687, -32'sd1033397, -32'sd2040735, -32'sd351460, 32'sd100388, 32'sd183100, 32'sd1254565, -32'sd334174, -32'sd186641, 32'sd222232, -32'sd409895, -32'sd168836, -32'sd2050761, 32'sd535077, -32'sd121481, 32'sd622633, 32'sd833391, -32'sd641302, -32'sd720012, -32'sd2569382, -32'sd499462, 32'sd1348441, 32'sd587499, 32'sd607649, 32'sd2034654, 32'sd2496144, 32'sd1967096, -32'sd204346, -32'sd579790, -32'sd1772653, -32'sd3998, -32'sd1863819, -32'sd1737862, -32'sd969903, 32'sd1153763, 32'sd85920, -32'sd460687, -32'sd865719, 32'sd641022, -32'sd1231657, -32'sd2257003, -32'sd2952717, -32'sd954240, 32'sd1312133, -32'sd407682, -32'sd520603, -32'sd1820759, 32'sd677235, 32'sd1437855, 32'sd144664, 32'sd1190819, 32'sd1696696, -32'sd147135, -32'sd597960, 32'sd2737521, 32'sd1037025, -32'sd2119684, -32'sd2149100, -32'sd1886538, 32'sd41185, -32'sd810573, 32'sd794839, 32'sd389774, -32'sd331354, -32'sd993949, 32'sd239114, -32'sd69588, -32'sd1472463, -32'sd1163778, -32'sd3264268, 32'sd1407758, 32'sd1437401, -32'sd2281698, -32'sd728218, -32'sd768896, 32'sd2018666, 32'sd1246428, 32'sd559313, -32'sd1275113, -32'sd245577, 32'sd760605, 32'sd318011, 32'sd776681, -32'sd1221353, -32'sd1756342, -32'sd1600662, -32'sd2271839, 32'sd199102, -32'sd1222476, -32'sd477651, -32'sd619590, 32'sd192982, 32'sd558706, -32'sd62050, -32'sd1020706, -32'sd224897, -32'sd864577, -32'sd3729303, 32'sd139585, -32'sd538607, -32'sd1997799, -32'sd548567, 32'sd1026782, 32'sd1313317, 32'sd85566, 32'sd749641, -32'sd1330319, 32'sd1620956, 32'sd1674429, -32'sd1181901, -32'sd1644008, -32'sd1191106, -32'sd3168987, -32'sd3096065, -32'sd1581143, 32'sd796322, -32'sd885876, -32'sd202571, 32'sd543087, 32'sd0, -32'sd223696, -32'sd143948, -32'sd455214, -32'sd1292353, -32'sd1969712, -32'sd1816655, -32'sd1572157, -32'sd2673049, -32'sd2768824, 32'sd427072, 32'sd1813426, 32'sd1165992, 32'sd294618, -32'sd1776549, 32'sd348194, 32'sd799109, 32'sd283677, -32'sd83473, -32'sd1680488, -32'sd399979, -32'sd683600, -32'sd597061, -32'sd586149, 32'sd657803, -32'sd1470914, 32'sd919786, 32'sd387033, -32'sd391325, 32'sd326684, -32'sd1513925, -32'sd1299480, -32'sd1199105, -32'sd3801009, -32'sd2918313, -32'sd2257100, -32'sd769006, 32'sd277047, 32'sd2886201, 32'sd1582160, 32'sd620955, 32'sd1080167, -32'sd549340, 32'sd1034383, -32'sd631582, -32'sd822469, -32'sd1613363, -32'sd626760, 32'sd110337, -32'sd1532713, -32'sd1954201, -32'sd1112974, 32'sd544436, -32'sd1643119, -32'sd490667, 32'sd1151817, -32'sd185374, 32'sd1002947, 32'sd408690, -32'sd216772, -32'sd1592323, -32'sd2600129, -32'sd3161908, -32'sd2977696, -32'sd309083, 32'sd1067131, 32'sd1370267, 32'sd357302, 32'sd1949808, 32'sd182651, -32'sd688633, 32'sd1222683, -32'sd79986, -32'sd591223, -32'sd2219115, -32'sd432627, -32'sd1526643, -32'sd1578610, -32'sd547124, -32'sd708392, -32'sd360336, 32'sd130197, 32'sd631573, -32'sd761991, 32'sd0, -32'sd431915, -32'sd2164076, -32'sd49538, -32'sd2592710, -32'sd1384412, -32'sd2362056, -32'sd932038, -32'sd2332610, 32'sd2015131, 32'sd3041212, 32'sd411421, -32'sd1957749, -32'sd2289304, -32'sd380979, -32'sd699415, 32'sd343516, -32'sd855702, -32'sd632549, 32'sd208781, 32'sd428492, 32'sd752465, -32'sd2397072, -32'sd49528, 32'sd41466, -32'sd1362758, -32'sd452692, 32'sd547441, -32'sd150611, -32'sd190690, -32'sd1645185, -32'sd72574, -32'sd1375833, 32'sd302388, -32'sd2280821, -32'sd1413717, -32'sd244655, 32'sd694742, 32'sd1654932, -32'sd1815003, -32'sd196526, 32'sd1097447, 32'sd1283164, 32'sd31988, -32'sd137427, 32'sd1024603, -32'sd998322, 32'sd1025293, -32'sd1936444, -32'sd2301976, -32'sd1291183, -32'sd800732, 32'sd1739856, 32'sd1523045, 32'sd1481259, 32'sd651970, -32'sd8321, -32'sd871220, 32'sd777624, -32'sd767152, -32'sd112669, -32'sd1626566, -32'sd1990819, -32'sd2522328, -32'sd1095730, -32'sd1377425, -32'sd106309, -32'sd513148, 32'sd460567, 32'sd508038, 32'sd2488484, -32'sd884575, 32'sd856322, 32'sd1056036, -32'sd807169, 32'sd541447, -32'sd2270838, -32'sd3020806, -32'sd1462907, -32'sd1211920, 32'sd485299, 32'sd930432, 32'sd1863785, 32'sd354840, 32'sd0, -32'sd310486, -32'sd342141, 32'sd616931, -32'sd839334, -32'sd1020924, -32'sd1299164, -32'sd2097381, -32'sd657358, 32'sd719733, -32'sd1595541, -32'sd639724, 32'sd1452899, 32'sd1643375, 32'sd1191144, -32'sd2227110, -32'sd277773, 32'sd52085, 32'sd734164, 32'sd561258, -32'sd316288, -32'sd41763, -32'sd143151, -32'sd2836196, -32'sd1083550, -32'sd1123479, -32'sd1189359, 32'sd0, 32'sd0, 32'sd0, 32'sd59570, 32'sd194737, 32'sd529550, 32'sd271888, -32'sd748382, -32'sd1172120, -32'sd1465197, -32'sd1145439, 32'sd39155, -32'sd923901, -32'sd1206829, -32'sd1526315, -32'sd1125162, -32'sd1941546, 32'sd915246, -32'sd952600, -32'sd45366, -32'sd1002384, -32'sd824106, -32'sd731031, 32'sd743431, -32'sd795786, -32'sd301718, 32'sd319083, -32'sd233557, 32'sd0, 32'sd0, 32'sd0, -32'sd486677, -32'sd15236, -32'sd2388228, 32'sd578662, 32'sd1681364, 32'sd1322728, 32'sd473947, 32'sd457754, -32'sd1687183, -32'sd1054333, -32'sd198010, 32'sd1157439, 32'sd2371885, 32'sd326719, 32'sd1949460, 32'sd1129306, 32'sd841572, 32'sd573279, 32'sd1069154, -32'sd133811, -32'sd82324, -32'sd280388, -32'sd519006, 32'sd568565, -32'sd236672, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd67386, -32'sd1439936, 32'sd400896, -32'sd92472, 32'sd1628285, 32'sd463300, 32'sd729684, -32'sd595703, -32'sd335974, 32'sd614161, -32'sd1041754, -32'sd367071, 32'sd557303, 32'sd310700, 32'sd1910352, 32'sd2307967, -32'sd90646, 32'sd334764, 32'sd87916, 32'sd41619, -32'sd1258086, 32'sd903987, 32'sd60976, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd136210, -32'sd480261, -32'sd501929, 32'sd932806, 32'sd2045191, 32'sd981934, 32'sd1498148, -32'sd344397, 32'sd1324406, 32'sd615589, 32'sd1478664, 32'sd1196752, 32'sd1300158, 32'sd1349895, -32'sd789433, -32'sd1322849, 32'sd409426, -32'sd185349, -32'sd245838, 32'sd790605, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd397405, 32'sd1270446, -32'sd116922, 32'sd1360388, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd31838, -32'sd498233, 32'sd43679, 32'sd1145555, -32'sd66471, -32'sd241404, 32'sd1480988, 32'sd684464, 32'sd188152, -32'sd825270, -32'sd1406143, -32'sd525524, -32'sd2120327, -32'sd31043, -32'sd1796961, 32'sd1192543, -32'sd352215, 32'sd38742, -32'sd200673, -32'sd338270, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd717789, -32'sd520921, 32'sd99096, 32'sd982081, 32'sd1163685, 32'sd723781, 32'sd302079, 32'sd1262344, 32'sd155517, 32'sd888073, 32'sd1625876, 32'sd1678513, -32'sd403559, 32'sd895078, 32'sd930490, 32'sd759359, -32'sd306803, 32'sd135272, 32'sd100996, 32'sd66853, 32'sd1303358, 32'sd1011276, 32'sd584275, -32'sd389254, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd906696, -32'sd527287, 32'sd905674, 32'sd169847, -32'sd1295361, 32'sd1039194, -32'sd180935, 32'sd1150223, 32'sd106471, 32'sd3741592, 32'sd2905636, 32'sd1610164, 32'sd537881, 32'sd1772706, 32'sd2041953, 32'sd822086, 32'sd1446017, -32'sd44938, -32'sd1735635, 32'sd961362, -32'sd72713, -32'sd1041302, 32'sd574849, -32'sd326793, -32'sd506019, 32'sd0, 32'sd0, -32'sd72469, 32'sd475949, -32'sd2046730, 32'sd188580, 32'sd2517005, -32'sd1088755, 32'sd251658, 32'sd139959, 32'sd554370, 32'sd2262844, 32'sd2313238, -32'sd296780, 32'sd2071483, 32'sd956636, -32'sd228651, -32'sd191865, -32'sd644368, -32'sd1085821, 32'sd1352949, 32'sd644954, -32'sd773521, -32'sd72691, 32'sd741561, 32'sd820988, -32'sd330486, -32'sd1588170, -32'sd743635, 32'sd0, 32'sd32354, -32'sd1125071, 32'sd186653, -32'sd704498, 32'sd2464499, 32'sd641837, 32'sd1680956, -32'sd984133, 32'sd1538562, 32'sd1572815, -32'sd957814, -32'sd3379784, -32'sd2212308, -32'sd1731954, 32'sd368317, -32'sd743049, -32'sd2291228, 32'sd67061, -32'sd74545, 32'sd1625867, 32'sd673488, 32'sd982359, 32'sd813477, -32'sd390178, 32'sd204839, -32'sd2137544, -32'sd53295, 32'sd0, -32'sd709851, 32'sd590202, -32'sd675546, -32'sd249770, 32'sd65473, -32'sd750843, -32'sd1367794, 32'sd1420442, -32'sd438901, 32'sd490515, -32'sd1161722, -32'sd3872860, -32'sd3515940, -32'sd613410, -32'sd1279596, 32'sd106111, -32'sd1605711, -32'sd2286751, -32'sd248740, 32'sd419284, -32'sd239687, 32'sd16117, -32'sd1631603, 32'sd1891204, 32'sd2064313, -32'sd848900, 32'sd795089, 32'sd415100, -32'sd134183, -32'sd725870, 32'sd747421, -32'sd984228, -32'sd1924604, -32'sd2139052, 32'sd833080, 32'sd725072, 32'sd2395468, -32'sd424974, -32'sd776784, -32'sd2898512, -32'sd3127757, -32'sd2960868, -32'sd2394402, -32'sd1394668, -32'sd1453725, -32'sd484702, -32'sd1861392, -32'sd170928, -32'sd804341, 32'sd78917, -32'sd1451605, -32'sd21049, -32'sd1309352, 32'sd1645478, -32'sd1565559, 32'sd94246, -32'sd556550, 32'sd642179, 32'sd1273285, -32'sd1836876, -32'sd2592776, -32'sd1347004, -32'sd947331, 32'sd2314268, 32'sd1046989, 32'sd726754, 32'sd74052, -32'sd1916851, -32'sd2260962, -32'sd1630475, 32'sd402546, -32'sd288508, 32'sd630626, -32'sd1387955, -32'sd829623, 32'sd878001, -32'sd1175953, -32'sd755958, 32'sd823603, -32'sd1234816, -32'sd376304, 32'sd1608653, -32'sd165765, -32'sd20843, -32'sd589139, 32'sd665969, 32'sd918678, 32'sd915946, 32'sd1602458, -32'sd2097318, -32'sd849781, -32'sd1697869, -32'sd449875, -32'sd311959, -32'sd1131608, 32'sd117894, -32'sd1102904, -32'sd1701616, 32'sd124650, 32'sd2315444, 32'sd1235298, 32'sd942283, -32'sd548267, 32'sd990683, -32'sd1130029, -32'sd521893, -32'sd3100602, -32'sd1742591, 32'sd378315, 32'sd724931, 32'sd519921, -32'sd118221, -32'sd1114935, -32'sd377207, 32'sd907827, 32'sd1876425, 32'sd1867835, -32'sd887861, -32'sd2032328, -32'sd1734531, -32'sd830100, -32'sd403786, -32'sd346590, -32'sd3244747, -32'sd2477250, -32'sd1602588, -32'sd454217, 32'sd1272375, 32'sd1280179, 32'sd28003, -32'sd298227, 32'sd307021, 32'sd1443859, -32'sd1982796, 32'sd471871, 32'sd1742529, -32'sd352075, 32'sd233023, -32'sd1363112, 32'sd939792, 32'sd820572, -32'sd578019, 32'sd583937, 32'sd1877354, 32'sd1920739, -32'sd743005, -32'sd695229, -32'sd2051297, -32'sd273426, -32'sd2259983, -32'sd2034669, -32'sd242859, -32'sd3714797, -32'sd4130853, -32'sd1194930, -32'sd2058385, -32'sd1263626, -32'sd3023495, -32'sd1286841, -32'sd1459316, 32'sd942469, -32'sd1042155, 32'sd451381, -32'sd1076563, -32'sd773024, 32'sd332847, -32'sd1195509, -32'sd488600, -32'sd821767, 32'sd663748, -32'sd968117, -32'sd808775, -32'sd86838, -32'sd531885, -32'sd369775, -32'sd1551390, -32'sd2209354, -32'sd277271, 32'sd924226, -32'sd412706, -32'sd414978, -32'sd698834, -32'sd1876830, -32'sd679763, -32'sd2450646, -32'sd2345058, -32'sd4353131, -32'sd2020643, -32'sd179523, 32'sd1894873, -32'sd1657109, 32'sd438849, -32'sd265209, 32'sd768724, -32'sd1189214, -32'sd178565, 32'sd508714, -32'sd1029297, -32'sd838685, -32'sd833966, -32'sd938887, -32'sd793085, -32'sd1023624, -32'sd2072258, -32'sd189627, 32'sd1780299, 32'sd1948169, -32'sd463835, 32'sd1657304, 32'sd330613, -32'sd2094956, -32'sd519761, -32'sd1684447, -32'sd1750684, -32'sd2337083, -32'sd365166, -32'sd464269, -32'sd1204904, -32'sd340477, 32'sd653168, -32'sd645272, 32'sd169762, -32'sd798069, 32'sd127300, 32'sd100758, 32'sd55230, -32'sd573235, -32'sd1848534, 32'sd260236, 32'sd1359941, -32'sd1901427, -32'sd2712704, 32'sd10501, 32'sd2113502, 32'sd1742394, 32'sd2435025, 32'sd1643623, 32'sd942700, -32'sd834040, -32'sd324655, -32'sd2561812, -32'sd650329, -32'sd1698685, -32'sd2483917, 32'sd228734, -32'sd196460, 32'sd817118, 32'sd3110948, 32'sd1225107, 32'sd640231, 32'sd306153, 32'sd1287331, 32'sd619231, -32'sd1199531, -32'sd410607, 32'sd491448, 32'sd2657847, 32'sd336221, 32'sd361455, 32'sd319275, 32'sd1438025, 32'sd738839, 32'sd2229961, 32'sd3678920, 32'sd3171339, 32'sd1652734, -32'sd1397701, -32'sd1057072, 32'sd936300, 32'sd997955, -32'sd478977, -32'sd2007301, -32'sd920971, 32'sd1091573, 32'sd536755, 32'sd2418377, 32'sd183785, -32'sd853651, -32'sd809161, -32'sd458922, -32'sd428226, -32'sd1408627, 32'sd1406727, 32'sd712647, 32'sd1264979, 32'sd1425118, 32'sd36028, -32'sd1208116, 32'sd2215491, 32'sd1736680, 32'sd1708696, 32'sd4192580, 32'sd2782951, 32'sd1642777, 32'sd785334, 32'sd1530936, 32'sd1627293, 32'sd1147712, 32'sd166286, -32'sd1721053, -32'sd30393, 32'sd1390617, 32'sd2729354, 32'sd2211587, -32'sd1149952, -32'sd876086, -32'sd928785, 32'sd0, -32'sd782258, -32'sd965876, 32'sd641582, -32'sd199476, -32'sd70700, 32'sd1445929, 32'sd988998, 32'sd1025326, 32'sd1040083, 32'sd449997, 32'sd2286210, 32'sd1090242, 32'sd226651, 32'sd160696, -32'sd1090021, 32'sd1693842, -32'sd57779, 32'sd1135589, 32'sd95988, 32'sd326702, 32'sd294385, 32'sd1631892, 32'sd582829, -32'sd840035, -32'sd412767, -32'sd2151377, 32'sd498245, -32'sd27578, 32'sd72919, 32'sd1610313, -32'sd752094, -32'sd865755, 32'sd1273546, 32'sd1452790, 32'sd355551, 32'sd1461512, 32'sd376415, 32'sd1591718, 32'sd1681801, 32'sd1430897, 32'sd1314062, 32'sd991068, 32'sd1781019, -32'sd349140, 32'sd2261042, 32'sd2070419, 32'sd667191, -32'sd542633, 32'sd102291, -32'sd698852, -32'sd1714570, -32'sd765472, 32'sd1658577, -32'sd1522982, -32'sd237012, 32'sd569147, -32'sd111481, 32'sd262180, -32'sd2659607, 32'sd407401, -32'sd754624, -32'sd328429, -32'sd1178305, -32'sd670773, 32'sd36086, 32'sd2668001, 32'sd984723, 32'sd1449470, 32'sd1123723, 32'sd1479469, 32'sd1161191, 32'sd273836, 32'sd1348007, 32'sd3175423, 32'sd139071, 32'sd1500994, 32'sd2584801, 32'sd920980, 32'sd946174, -32'sd3976187, 32'sd445987, -32'sd26300, -32'sd1056904, 32'sd0, -32'sd1259938, -32'sd271162, -32'sd2843446, 32'sd2430916, -32'sd1714855, -32'sd604689, 32'sd272392, 32'sd1404158, 32'sd3414624, 32'sd2829574, 32'sd2035517, 32'sd231241, -32'sd173734, 32'sd503123, -32'sd1324751, -32'sd1786955, 32'sd625200, 32'sd2707044, 32'sd180412, 32'sd1046468, 32'sd2409372, 32'sd1092866, 32'sd297482, -32'sd2236309, 32'sd76519, 32'sd1147553, -32'sd931607, -32'sd893498, 32'sd1377112, 32'sd986777, -32'sd743954, 32'sd1662221, 32'sd766741, -32'sd336508, 32'sd509051, 32'sd105617, 32'sd2332200, 32'sd1573767, 32'sd58947, 32'sd1311174, 32'sd1542075, -32'sd623947, -32'sd1306751, 32'sd279031, -32'sd511072, 32'sd1384819, 32'sd2163060, 32'sd2195501, 32'sd1656269, 32'sd462136, 32'sd87499, -32'sd2140912, -32'sd1667929, 32'sd1285860, -32'sd326764, -32'sd69266, -32'sd938165, -32'sd1181198, 32'sd132738, -32'sd1689923, -32'sd93667, -32'sd831315, -32'sd1515377, -32'sd1203354, 32'sd241628, 32'sd259195, -32'sd1408464, -32'sd759752, -32'sd503983, -32'sd734608, -32'sd364349, 32'sd312789, -32'sd2387783, -32'sd128805, 32'sd1045774, 32'sd1033813, -32'sd664657, -32'sd598421, -32'sd1166102, 32'sd46909, -32'sd278252, -32'sd256996, -32'sd140099, 32'sd0, -32'sd56559, 32'sd2632513, 32'sd534617, 32'sd81273, -32'sd824196, -32'sd156895, -32'sd1266388, -32'sd1369293, -32'sd295912, -32'sd464574, -32'sd2335952, -32'sd133422, -32'sd1725668, -32'sd513856, -32'sd772504, -32'sd3158870, -32'sd2362803, 32'sd634935, -32'sd325626, -32'sd817004, 32'sd606439, -32'sd567523, -32'sd2279178, -32'sd1264643, 32'sd646108, 32'sd695481, 32'sd0, 32'sd0, 32'sd0, 32'sd567765, -32'sd2053106, 32'sd500297, -32'sd1716285, -32'sd1169001, -32'sd2233706, -32'sd3859062, -32'sd2654863, -32'sd2669844, -32'sd3745572, -32'sd2220471, -32'sd350273, -32'sd2365561, -32'sd789370, 32'sd732554, 32'sd272938, -32'sd1005122, -32'sd1727718, -32'sd1886249, -32'sd67127, -32'sd954754, 32'sd185787, -32'sd104827, -32'sd224652, 32'sd457954, 32'sd0, 32'sd0, 32'sd0, -32'sd728249, -32'sd466087, -32'sd1206470, -32'sd641926, -32'sd912011, -32'sd837660, -32'sd1125324, -32'sd707711, -32'sd2479466, -32'sd1244931, 32'sd27308, -32'sd3354699, -32'sd807701, 32'sd556924, 32'sd1123216, -32'sd1487845, 32'sd693147, -32'sd2553020, -32'sd8834, -32'sd2194241, -32'sd910328, -32'sd1114591, 32'sd481007, 32'sd528882, 32'sd1248650, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd438081, 32'sd199557, 32'sd102470, -32'sd16052, -32'sd1072314, -32'sd1045215, 32'sd580327, 32'sd599156, 32'sd452631, -32'sd1155487, 32'sd1230603, 32'sd76209, -32'sd82762, 32'sd944540, -32'sd549304, -32'sd1993969, -32'sd736896, -32'sd902840, -32'sd774687, 32'sd33128, -32'sd1478792, 32'sd470488, -32'sd582897, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd731926, -32'sd774890, -32'sd545262, 32'sd268335, -32'sd978569, -32'sd754467, 32'sd58759, 32'sd1120515, 32'sd392404, -32'sd214168, 32'sd993246, 32'sd683067, -32'sd474817, -32'sd903818, -32'sd714075, -32'sd363813, 32'sd574310, -32'sd1562053, -32'sd40422, 32'sd223640, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd188671, 32'sd219479, -32'sd652772, -32'sd842628, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd74643, -32'sd1586999, -32'sd97414, -32'sd1689143, -32'sd1295350, -32'sd1839601, -32'sd2161872, -32'sd298660, 32'sd518316, -32'sd989343, -32'sd655447, 32'sd152669, -32'sd1253488, -32'sd2035877, -32'sd435213, -32'sd758447, 32'sd392934, -32'sd1209676, 32'sd153371, -32'sd274449, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd772563, -32'sd192730, -32'sd1355302, -32'sd1615048, -32'sd893708, -32'sd1142338, -32'sd765860, -32'sd1644311, -32'sd1022296, -32'sd2489010, -32'sd2091137, -32'sd2179511, -32'sd1847668, -32'sd1892808, -32'sd586681, -32'sd1492791, 32'sd471869, 32'sd258494, 32'sd284077, -32'sd1137335, 32'sd604344, -32'sd1410606, -32'sd1410473, -32'sd1374971, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd191938, -32'sd606979, -32'sd1401977, 32'sd563144, -32'sd129631, -32'sd1674953, -32'sd599466, -32'sd2419050, -32'sd797776, -32'sd2746156, -32'sd1655133, -32'sd4447744, -32'sd1830011, -32'sd347884, 32'sd524130, -32'sd2648619, -32'sd559435, -32'sd2045865, -32'sd2106574, 32'sd939587, 32'sd1202407, 32'sd540323, -32'sd736789, -32'sd749570, -32'sd927239, 32'sd0, 32'sd0, 32'sd495084, -32'sd1773445, -32'sd521528, -32'sd1334664, -32'sd398913, -32'sd602793, -32'sd776380, -32'sd1993501, -32'sd4321511, -32'sd724660, -32'sd1159754, -32'sd1981007, -32'sd4116140, -32'sd3056413, 32'sd640714, -32'sd612168, -32'sd739438, 32'sd66209, -32'sd2743462, -32'sd173756, 32'sd82097, -32'sd165909, -32'sd286271, -32'sd1119783, -32'sd1115170, -32'sd17878, -32'sd380580, 32'sd0, -32'sd155799, -32'sd2042773, -32'sd2661680, -32'sd1405495, 32'sd1074294, 32'sd864127, 32'sd143410, 32'sd596948, 32'sd433768, 32'sd445640, 32'sd1681252, 32'sd469564, -32'sd1700907, -32'sd163617, 32'sd1041014, -32'sd802319, -32'sd149895, 32'sd9942, 32'sd450736, -32'sd2500394, -32'sd1796577, -32'sd1810573, -32'sd3003276, -32'sd803159, -32'sd1841134, -32'sd87327, -32'sd1795662, 32'sd0, 32'sd198421, 32'sd1575304, 32'sd1108194, 32'sd1411015, 32'sd1842208, -32'sd392265, -32'sd370484, 32'sd1379002, 32'sd2813930, 32'sd2026983, 32'sd872249, 32'sd386213, -32'sd711637, -32'sd1754819, 32'sd983256, 32'sd1938254, 32'sd2753121, 32'sd2234774, 32'sd1156307, 32'sd37310, 32'sd979322, -32'sd351094, -32'sd3042419, -32'sd2273180, -32'sd1237324, -32'sd2333749, -32'sd1884988, -32'sd778171, 32'sd666427, 32'sd911130, 32'sd406673, 32'sd3261335, -32'sd633525, 32'sd1653054, 32'sd2345457, 32'sd406973, 32'sd1112010, -32'sd428108, -32'sd559307, -32'sd2459700, -32'sd2061807, -32'sd631516, -32'sd612834, 32'sd386649, -32'sd603619, 32'sd1107684, 32'sd363045, 32'sd776071, 32'sd1249658, -32'sd408165, -32'sd318840, 32'sd320264, -32'sd828388, -32'sd3512851, -32'sd927560, 32'sd127597, 32'sd1161425, 32'sd1154224, -32'sd745591, -32'sd300744, -32'sd355482, -32'sd196286, 32'sd1359844, 32'sd1273120, 32'sd912622, 32'sd1457733, -32'sd218997, -32'sd1185718, -32'sd2915096, 32'sd164067, 32'sd716172, 32'sd337342, -32'sd1693582, 32'sd1117290, -32'sd250817, -32'sd1028897, 32'sd20085, -32'sd2467549, -32'sd1273054, 32'sd866732, -32'sd654154, -32'sd1566977, -32'sd1724927, -32'sd96898, -32'sd691697, -32'sd170635, -32'sd530018, 32'sd1801002, -32'sd585407, 32'sd324093, -32'sd122283, 32'sd1054809, 32'sd2334749, 32'sd1573586, 32'sd1568833, 32'sd1775959, -32'sd1471571, 32'sd2014317, -32'sd660966, -32'sd2424390, -32'sd639930, -32'sd874999, -32'sd477488, -32'sd951969, -32'sd1058211, -32'sd2278480, -32'sd2697452, 32'sd773659, 32'sd4043, -32'sd438355, 32'sd647255, -32'sd17504, 32'sd283008, 32'sd874613, -32'sd747864, 32'sd1929404, -32'sd676348, -32'sd338209, -32'sd1740214, 32'sd2054701, 32'sd3672621, 32'sd692048, 32'sd788793, -32'sd1059139, 32'sd1026413, 32'sd1917673, -32'sd1836124, -32'sd2074530, -32'sd2293166, -32'sd1560304, 32'sd174353, -32'sd746548, -32'sd1498839, -32'sd3125104, -32'sd2066888, 32'sd112702, 32'sd324546, -32'sd231866, -32'sd1135105, -32'sd865916, -32'sd872058, 32'sd1919641, 32'sd1127923, -32'sd687723, -32'sd2934891, -32'sd1763518, -32'sd520335, 32'sd2185357, 32'sd2424876, 32'sd479359, 32'sd1024617, -32'sd1330830, -32'sd1176842, 32'sd610498, 32'sd973864, -32'sd1783551, -32'sd107652, 32'sd449299, 32'sd2365310, 32'sd1456303, -32'sd594893, 32'sd344470, -32'sd354304, 32'sd89209, -32'sd450975, -32'sd18461, -32'sd343864, -32'sd1062669, -32'sd1148882, 32'sd1407407, -32'sd880491, 32'sd1914136, -32'sd75510, 32'sd1366609, 32'sd1288100, 32'sd2020289, 32'sd484854, 32'sd1614638, -32'sd227528, -32'sd2785300, -32'sd1309498, -32'sd2027431, -32'sd979436, -32'sd418081, -32'sd684120, 32'sd2102311, 32'sd2143366, -32'sd558739, 32'sd626640, 32'sd507306, -32'sd1247105, -32'sd942185, 32'sd571164, -32'sd362299, 32'sd695573, -32'sd820505, -32'sd598852, -32'sd790930, -32'sd1127918, -32'sd219177, -32'sd664473, 32'sd1656321, 32'sd1195620, 32'sd1312763, -32'sd488787, 32'sd1424205, 32'sd1304926, -32'sd1499215, 32'sd1241262, -32'sd899182, 32'sd1242403, 32'sd256215, 32'sd22088, 32'sd2229945, 32'sd729393, 32'sd735067, 32'sd436715, -32'sd710451, -32'sd1545318, -32'sd1438253, -32'sd975459, -32'sd47085, -32'sd846582, -32'sd909131, -32'sd1059333, -32'sd1351709, -32'sd1053531, -32'sd382746, 32'sd340594, 32'sd888868, 32'sd894856, 32'sd60678, 32'sd1059301, 32'sd1487635, 32'sd1909026, 32'sd520703, 32'sd2022242, 32'sd2435719, 32'sd2139877, 32'sd125134, 32'sd2473371, 32'sd3904672, 32'sd3116500, -32'sd58156, -32'sd618916, -32'sd3005269, -32'sd2910662, -32'sd1844971, 32'sd386697, -32'sd2369663, -32'sd688988, -32'sd1257737, -32'sd1062631, -32'sd1037656, -32'sd1048994, 32'sd136727, -32'sd179105, -32'sd476685, 32'sd1853424, -32'sd600298, 32'sd1247090, 32'sd1333528, 32'sd292149, 32'sd483964, 32'sd663622, 32'sd1977962, 32'sd1920650, 32'sd1507101, 32'sd3980427, 32'sd3013254, 32'sd284805, 32'sd52096, -32'sd512878, -32'sd398973, -32'sd2118141, -32'sd1738960, -32'sd1695748, -32'sd1032664, 32'sd839352, 32'sd439978, -32'sd374327, -32'sd435819, -32'sd133841, -32'sd1454186, -32'sd2233316, 32'sd727173, 32'sd1160922, 32'sd491768, 32'sd657529, 32'sd955569, 32'sd987545, 32'sd837922, 32'sd1910946, 32'sd1073070, 32'sd1710148, 32'sd1044190, 32'sd924314, -32'sd455134, 32'sd121759, -32'sd476667, 32'sd36633, -32'sd162992, -32'sd2742420, -32'sd2321873, -32'sd2176963, -32'sd2675402, -32'sd874363, 32'sd0, -32'sd1883684, 32'sd201108, -32'sd2165803, -32'sd2260463, -32'sd598019, 32'sd1396331, 32'sd1775969, 32'sd115707, 32'sd1720377, -32'sd117166, 32'sd949629, -32'sd364029, 32'sd251674, 32'sd1068945, 32'sd590351, 32'sd1046622, 32'sd955359, 32'sd568121, -32'sd2812, -32'sd2144416, -32'sd941454, 32'sd287347, 32'sd67669, -32'sd837742, 32'sd974595, -32'sd2863827, -32'sd893973, -32'sd1303780, -32'sd166809, 32'sd734851, -32'sd2126909, -32'sd325716, -32'sd2914179, -32'sd779240, 32'sd1937550, 32'sd1892196, 32'sd560210, 32'sd646328, -32'sd406113, 32'sd448806, 32'sd1025416, 32'sd355897, 32'sd1961751, -32'sd904129, 32'sd875742, -32'sd1240726, -32'sd875466, -32'sd2573097, -32'sd834509, 32'sd1961851, 32'sd1410590, -32'sd1866711, -32'sd600215, -32'sd155507, -32'sd2009677, -32'sd661655, -32'sd23350, -32'sd254142, -32'sd948725, -32'sd1441607, -32'sd2056269, -32'sd3319550, -32'sd935340, 32'sd836430, -32'sd77814, 32'sd25700, 32'sd379121, -32'sd1084033, -32'sd1973126, 32'sd2513100, 32'sd1301455, 32'sd429987, 32'sd487774, -32'sd1007509, -32'sd1510512, -32'sd2654958, -32'sd1791558, -32'sd258200, -32'sd774265, 32'sd427779, 32'sd572140, 32'sd29786, -32'sd1160210, 32'sd0, -32'sd60723, -32'sd1368930, -32'sd828212, -32'sd2882548, -32'sd4265087, -32'sd4484801, 32'sd117836, -32'sd2174663, -32'sd1112494, 32'sd535889, -32'sd1819284, -32'sd2131865, -32'sd1350589, 32'sd1648076, 32'sd436784, 32'sd659168, 32'sd156435, -32'sd2349129, -32'sd2927399, -32'sd3365051, -32'sd477494, -32'sd198607, 32'sd556485, -32'sd212666, 32'sd816531, -32'sd1001060, -32'sd51596, -32'sd231004, -32'sd1920840, -32'sd681781, -32'sd357769, -32'sd425184, -32'sd2681325, -32'sd1668545, -32'sd2320554, -32'sd1873154, -32'sd555493, 32'sd136246, -32'sd400452, -32'sd1804001, -32'sd2231845, -32'sd2407068, -32'sd1718357, 32'sd1765760, 32'sd590536, -32'sd2515608, -32'sd2369460, -32'sd3074256, -32'sd972392, -32'sd2629390, -32'sd278809, -32'sd1027782, -32'sd14610, 32'sd917449, 32'sd288873, -32'sd1404695, -32'sd1620905, -32'sd722103, -32'sd964707, 32'sd17315, -32'sd114947, -32'sd724826, -32'sd2746985, -32'sd3457824, -32'sd1198119, 32'sd640294, -32'sd1676383, 32'sd244105, -32'sd1636836, -32'sd1149367, -32'sd2976237, -32'sd392646, -32'sd1975846, -32'sd819981, -32'sd2370805, -32'sd1558669, -32'sd4116713, -32'sd813868, -32'sd1789245, -32'sd1078648, 32'sd588336, -32'sd3996, 32'sd351546, 32'sd0, -32'sd669374, -32'sd2075171, -32'sd962552, -32'sd801211, -32'sd288870, -32'sd107812, -32'sd489160, -32'sd1892320, -32'sd1673852, -32'sd1690909, -32'sd2425313, -32'sd1425209, 32'sd1003423, 32'sd470178, -32'sd1609387, -32'sd304412, -32'sd2021275, 32'sd165036, -32'sd804981, -32'sd1979549, -32'sd2943919, -32'sd804801, -32'sd1916631, -32'sd2216692, 32'sd243552, 32'sd716007, 32'sd0, 32'sd0, 32'sd0, 32'sd41847, -32'sd1144855, 32'sd1912967, 32'sd1262660, -32'sd495490, -32'sd65534, 32'sd216294, -32'sd1101570, -32'sd198864, -32'sd246765, -32'sd240439, 32'sd684472, -32'sd1033378, -32'sd794678, 32'sd568909, 32'sd729411, 32'sd374447, -32'sd351774, -32'sd1123244, -32'sd3364796, -32'sd1008940, -32'sd1086076, -32'sd977842, -32'sd1498361, -32'sd790929, 32'sd0, 32'sd0, 32'sd0, 32'sd423775, 32'sd283891, 32'sd577400, 32'sd705753, 32'sd1022031, -32'sd591833, -32'sd556601, -32'sd973500, 32'sd1178498, 32'sd160311, 32'sd50528, -32'sd433608, -32'sd1722624, 32'sd417893, 32'sd2950890, 32'sd2037160, 32'sd744042, -32'sd887062, -32'sd665519, -32'sd3377875, -32'sd371126, 32'sd36139, -32'sd147825, 32'sd379157, -32'sd333749, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd690448, -32'sd1047060, -32'sd1540447, 32'sd701280, 32'sd3206260, 32'sd555750, 32'sd403826, -32'sd243400, -32'sd1094751, -32'sd997915, 32'sd2802700, 32'sd210807, -32'sd770591, 32'sd867891, 32'sd1260406, -32'sd167750, -32'sd28923, -32'sd383311, -32'sd1506228, 32'sd1126746, 32'sd667399, -32'sd385384, -32'sd66427, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1472418, 32'sd428123, 32'sd111425, -32'sd1290640, -32'sd1882398, -32'sd660987, 32'sd181936, 32'sd1508865, -32'sd468639, 32'sd488607, 32'sd92349, -32'sd436113, 32'sd221272, -32'sd834198, 32'sd1384578, -32'sd1150276, -32'sd1305001, -32'sd758432, -32'sd510064, -32'sd1448868, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd924579, 32'sd739858, 32'sd500307, -32'sd641398, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd530252, 32'sd81442, 32'sd623418, -32'sd328497, -32'sd1207495, 32'sd1254704, 32'sd914427, -32'sd493861, -32'sd492881, -32'sd2120501, -32'sd492108, 32'sd46806, 32'sd409301, 32'sd496698, -32'sd137060, -32'sd17354, -32'sd280261, 32'sd596312, 32'sd1472555, 32'sd406174, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1021565, 32'sd796183, 32'sd199946, 32'sd2753, 32'sd404167, -32'sd196861, 32'sd85810, -32'sd1516620, -32'sd843793, 32'sd659978, 32'sd1031962, 32'sd375495, -32'sd997402, -32'sd538762, 32'sd318062, 32'sd247013, -32'sd298828, 32'sd1911906, -32'sd58272, -32'sd1154697, -32'sd1107212, 32'sd151458, 32'sd332340, 32'sd1450480, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1074386, 32'sd1114624, -32'sd626943, -32'sd243874, -32'sd2061904, -32'sd2208126, -32'sd1987068, -32'sd1567369, -32'sd118126, -32'sd539639, 32'sd1405487, -32'sd2018164, 32'sd1395220, -32'sd2307896, -32'sd918042, -32'sd341960, -32'sd2451268, -32'sd1057586, 32'sd385511, 32'sd209925, -32'sd86826, -32'sd1264237, -32'sd1125629, -32'sd1952891, -32'sd216566, 32'sd0, 32'sd0, 32'sd1094035, 32'sd731918, 32'sd210044, 32'sd749735, 32'sd1190110, -32'sd476550, -32'sd1544936, -32'sd505350, -32'sd1344754, -32'sd906049, -32'sd1885330, -32'sd625676, 32'sd348786, -32'sd1078826, -32'sd48596, -32'sd3042182, -32'sd381247, -32'sd3102012, -32'sd785830, -32'sd188468, -32'sd1129441, -32'sd668879, 32'sd209082, 32'sd1409067, 32'sd92594, 32'sd429887, -32'sd471230, 32'sd0, 32'sd1273046, -32'sd766611, 32'sd1606023, 32'sd992609, -32'sd1294017, 32'sd346955, 32'sd609077, 32'sd320856, -32'sd404310, -32'sd343981, -32'sd1905728, -32'sd119346, -32'sd442899, -32'sd578682, 32'sd941711, -32'sd875741, -32'sd2119035, -32'sd1944555, -32'sd1496220, -32'sd909553, -32'sd1635478, -32'sd651117, -32'sd2439863, -32'sd1654704, -32'sd1234014, -32'sd1140555, 32'sd163070, 32'sd0, 32'sd565102, 32'sd581800, -32'sd2050380, -32'sd764806, -32'sd828334, 32'sd423624, -32'sd1860695, -32'sd1395362, -32'sd1084625, -32'sd2498452, -32'sd656991, 32'sd275375, -32'sd889208, -32'sd360702, -32'sd1052115, -32'sd2253172, -32'sd2363888, -32'sd979165, -32'sd3452391, -32'sd1557091, -32'sd792082, 32'sd280975, 32'sd1021205, -32'sd2621489, -32'sd3294865, -32'sd972896, -32'sd568282, 32'sd615021, -32'sd126548, -32'sd1808803, 32'sd644664, 32'sd55768, 32'sd83651, -32'sd410647, -32'sd271310, -32'sd3027589, -32'sd3017430, -32'sd1684546, -32'sd1109486, -32'sd1817506, -32'sd486426, -32'sd3526210, -32'sd992882, -32'sd441509, 32'sd886659, 32'sd351300, -32'sd765139, -32'sd895543, 32'sd881990, -32'sd655139, 32'sd248364, -32'sd341428, -32'sd1057732, 32'sd22789, 32'sd1503925, -32'sd774136, -32'sd1136058, 32'sd1438291, -32'sd499329, 32'sd153718, -32'sd1065794, -32'sd611981, 32'sd603592, -32'sd1058490, -32'sd1748648, -32'sd1683823, -32'sd931225, -32'sd863225, -32'sd1202364, -32'sd979439, -32'sd104868, 32'sd1298719, 32'sd2228171, -32'sd245852, -32'sd2024192, -32'sd1429988, -32'sd1234659, 32'sd509113, -32'sd934133, 32'sd1806337, -32'sd332618, 32'sd1313979, -32'sd59727, 32'sd436768, -32'sd157093, 32'sd1034573, -32'sd249021, -32'sd426366, -32'sd1700796, 32'sd273015, 32'sd160059, -32'sd1610541, -32'sd2192472, -32'sd514142, 32'sd900916, -32'sd615067, -32'sd563894, -32'sd2011847, 32'sd17001, 32'sd1363107, 32'sd1439073, 32'sd2693094, 32'sd1606562, -32'sd59857, -32'sd1488343, -32'sd1502302, 32'sd582568, 32'sd1605481, 32'sd544079, 32'sd397167, 32'sd744417, -32'sd332944, 32'sd668300, 32'sd1464538, 32'sd381055, 32'sd1082745, -32'sd330081, -32'sd155918, -32'sd657437, -32'sd1894020, 32'sd958930, 32'sd611316, 32'sd1770640, -32'sd1244414, -32'sd412216, 32'sd509272, 32'sd2864309, 32'sd2447280, 32'sd1444687, 32'sd2622926, 32'sd2709007, -32'sd822421, -32'sd1827944, -32'sd3074101, -32'sd848604, 32'sd309671, 32'sd871870, -32'sd883021, -32'sd1443482, -32'sd800399, 32'sd1509849, 32'sd2190120, 32'sd373057, -32'sd1113988, -32'sd1130017, 32'sd1474208, 32'sd652319, -32'sd419198, -32'sd5271, -32'sd1070248, 32'sd364528, 32'sd1856676, 32'sd45913, -32'sd2008415, -32'sd975640, 32'sd2140927, 32'sd1725251, 32'sd3909202, 32'sd1758408, -32'sd40354, 32'sd689152, -32'sd174660, -32'sd252499, -32'sd767908, -32'sd78246, -32'sd1023470, -32'sd47708, 32'sd1191544, 32'sd287121, 32'sd215995, 32'sd420359, 32'sd265989, -32'sd1784989, 32'sd1187898, -32'sd352732, 32'sd544801, 32'sd1196825, 32'sd1492693, 32'sd1954095, 32'sd2028872, -32'sd1259612, -32'sd1923458, -32'sd361579, -32'sd105021, 32'sd78645, 32'sd1273257, 32'sd2906943, 32'sd501138, -32'sd860552, 32'sd1031922, -32'sd1156712, 32'sd550458, 32'sd681187, -32'sd614617, 32'sd275483, 32'sd585734, 32'sd532640, -32'sd299725, -32'sd273735, 32'sd554666, 32'sd72777, 32'sd930951, 32'sd759259, 32'sd1166393, -32'sd973419, 32'sd314442, 32'sd2204696, 32'sd2292017, -32'sd354814, -32'sd1584014, -32'sd875656, -32'sd1303399, 32'sd2736005, 32'sd2589934, 32'sd3095661, 32'sd232519, 32'sd657202, -32'sd250725, 32'sd1181204, -32'sd1051608, 32'sd725278, 32'sd664163, -32'sd679037, -32'sd746354, -32'sd764281, -32'sd228408, -32'sd964193, -32'sd1579157, -32'sd340656, 32'sd1331207, 32'sd944519, -32'sd747004, 32'sd1900609, -32'sd64780, -32'sd218172, 32'sd1044028, -32'sd1445269, -32'sd1175884, 32'sd1423626, 32'sd658113, 32'sd4246735, 32'sd2117214, 32'sd3669639, 32'sd672934, -32'sd2027223, -32'sd1450128, -32'sd555149, -32'sd1707006, 32'sd1583952, -32'sd1812866, 32'sd1926206, 32'sd70309, -32'sd286195, 32'sd989972, 32'sd444847, 32'sd1628068, 32'sd1304466, -32'sd581467, 32'sd623748, 32'sd1414209, 32'sd1678751, -32'sd92488, 32'sd591397, 32'sd2347491, -32'sd1880379, -32'sd1854294, 32'sd740085, -32'sd212870, 32'sd1906838, 32'sd4720668, 32'sd174186, -32'sd2622907, -32'sd645998, -32'sd258553, -32'sd456284, 32'sd114156, -32'sd483306, 32'sd1280684, -32'sd803590, 32'sd806947, -32'sd504498, 32'sd376195, -32'sd904820, -32'sd1114933, 32'sd1314663, -32'sd1008798, 32'sd1376748, 32'sd1101860, 32'sd2380878, 32'sd1435321, 32'sd1728249, 32'sd1567909, -32'sd2818267, -32'sd3575941, -32'sd1083973, 32'sd1146593, 32'sd4081499, 32'sd2193063, -32'sd1352715, -32'sd2377971, -32'sd1671898, -32'sd1176647, -32'sd613237, -32'sd2125345, -32'sd1655243, 32'sd654395, -32'sd761650, 32'sd0, 32'sd1107231, 32'sd1321437, -32'sd2214370, 32'sd646547, -32'sd148877, 32'sd1359539, 32'sd295156, 32'sd1219249, 32'sd2987808, 32'sd1361717, 32'sd2942323, -32'sd209445, -32'sd1116846, -32'sd703583, 32'sd2802499, 32'sd1778365, 32'sd216602, 32'sd1290304, -32'sd878288, -32'sd2691456, -32'sd1024449, -32'sd305114, 32'sd403177, -32'sd486437, 32'sd51680, 32'sd1041687, -32'sd386761, -32'sd1161235, -32'sd661712, 32'sd709569, -32'sd1156456, -32'sd341607, -32'sd1385760, -32'sd664806, 32'sd934275, 32'sd2781834, 32'sd1901009, -32'sd303197, 32'sd568944, -32'sd798318, -32'sd1877332, 32'sd851678, 32'sd1663533, -32'sd50497, -32'sd752418, -32'sd595002, -32'sd1139317, -32'sd1925194, -32'sd1899253, -32'sd352641, 32'sd761817, -32'sd2463674, 32'sd1284046, -32'sd793714, -32'sd877681, 32'sd56468, 32'sd129715, 32'sd660371, 32'sd1224794, 32'sd505466, -32'sd639071, -32'sd664853, 32'sd2477888, 32'sd1861967, -32'sd1920446, -32'sd783011, -32'sd402205, -32'sd1083364, -32'sd2115915, -32'sd976652, 32'sd519708, -32'sd2605719, 32'sd56634, -32'sd974597, 32'sd810560, -32'sd1432354, -32'sd104196, -32'sd322650, -32'sd1772770, -32'sd636148, 32'sd1172422, -32'sd1387309, 32'sd1544887, 32'sd0, -32'sd331584, 32'sd822897, 32'sd361495, 32'sd230639, -32'sd579525, -32'sd962843, 32'sd981988, -32'sd1840965, -32'sd2926021, -32'sd1218659, -32'sd1676144, -32'sd347434, -32'sd947430, -32'sd2156730, -32'sd3799041, -32'sd1033279, -32'sd331361, 32'sd656992, -32'sd871350, -32'sd978267, 32'sd218880, -32'sd766276, -32'sd423539, 32'sd465131, -32'sd133229, -32'sd989555, 32'sd543068, -32'sd107122, 32'sd634306, -32'sd398426, -32'sd246766, -32'sd628277, 32'sd2202947, 32'sd178776, -32'sd419327, -32'sd1171778, -32'sd1036979, -32'sd2166260, -32'sd2415399, -32'sd1344806, -32'sd2104612, -32'sd2394752, -32'sd3320818, -32'sd655967, -32'sd675780, -32'sd1776032, 32'sd1518651, -32'sd96297, -32'sd706309, 32'sd985316, -32'sd83559, -32'sd60659, 32'sd1022733, 32'sd889529, 32'sd905912, 32'sd661661, 32'sd17778, 32'sd1669631, -32'sd555338, -32'sd90002, -32'sd57105, 32'sd395581, -32'sd1559705, -32'sd3080681, -32'sd941327, -32'sd1101018, 32'sd441059, -32'sd913866, -32'sd2142401, -32'sd254265, -32'sd1568924, -32'sd1094718, -32'sd1952027, -32'sd1735964, 32'sd164767, -32'sd1119018, 32'sd824171, 32'sd1027447, -32'sd1007111, -32'sd354022, 32'sd753433, 32'sd99377, 32'sd2440808, 32'sd0, 32'sd614260, -32'sd573066, -32'sd320143, -32'sd2341333, -32'sd2109659, -32'sd1478296, -32'sd874984, -32'sd652122, -32'sd253145, 32'sd706319, -32'sd979797, -32'sd615685, -32'sd817825, 32'sd114703, -32'sd670409, -32'sd259671, -32'sd1503682, -32'sd1998936, 32'sd125761, 32'sd663252, -32'sd41607, 32'sd737768, 32'sd623104, 32'sd1676481, 32'sd94892, -32'sd1264705, 32'sd0, 32'sd0, 32'sd0, 32'sd33370, -32'sd833101, -32'sd732180, -32'sd945571, -32'sd2614733, -32'sd169626, 32'sd640925, 32'sd36492, -32'sd784422, -32'sd1621326, 32'sd40273, 32'sd414056, -32'sd1059953, -32'sd1269573, 32'sd32036, -32'sd556026, -32'sd984394, 32'sd1462201, -32'sd7503, 32'sd1246775, 32'sd1901019, 32'sd1752604, 32'sd42497, 32'sd62966, 32'sd905684, 32'sd0, 32'sd0, 32'sd0, 32'sd1309159, -32'sd1272254, -32'sd562901, -32'sd202900, -32'sd778004, -32'sd826568, 32'sd244620, 32'sd60553, -32'sd997260, -32'sd178022, 32'sd433532, -32'sd1137001, 32'sd401364, 32'sd751505, -32'sd491854, -32'sd1023159, 32'sd1049493, -32'sd365714, 32'sd1183472, 32'sd365848, 32'sd1321193, -32'sd454184, -32'sd1287363, 32'sd1644268, -32'sd218375, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1495706, -32'sd398260, 32'sd1407830, 32'sd1644173, 32'sd935021, -32'sd332736, 32'sd505640, -32'sd1314504, 32'sd1784923, 32'sd865202, 32'sd854687, -32'sd675263, 32'sd494238, -32'sd103759, -32'sd1304294, -32'sd426242, -32'sd845784, -32'sd1261263, 32'sd428507, -32'sd311436, 32'sd254396, 32'sd1385800, 32'sd744418, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1594414, 32'sd866715, 32'sd114438, 32'sd871610, -32'sd1263173, 32'sd762248, 32'sd1515707, 32'sd255649, -32'sd210194, 32'sd1656678, 32'sd231893, 32'sd357102, 32'sd577456, -32'sd482761, -32'sd51952, 32'sd1017199, 32'sd867409, -32'sd704125, 32'sd2110349, -32'sd88845, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd597803, 32'sd269396, -32'sd872446, 32'sd162620, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1911541, -32'sd434373, -32'sd119520, 32'sd1540983, 32'sd398297, 32'sd634908, 32'sd847487, -32'sd1516710, -32'sd145256, 32'sd1929528, -32'sd105612, 32'sd449168, 32'sd979130, 32'sd274902, 32'sd1836889, -32'sd459841, 32'sd836385, 32'sd2494553, 32'sd2457415, 32'sd793311, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1651903, 32'sd881229, 32'sd898957, 32'sd218402, -32'sd1802319, 32'sd234946, 32'sd198666, 32'sd2212091, -32'sd47448, 32'sd856605, 32'sd498473, 32'sd771440, -32'sd1619557, 32'sd87827, 32'sd1113234, 32'sd2401454, 32'sd1524938, 32'sd1218228, 32'sd891481, -32'sd283261, 32'sd3002349, 32'sd1529822, 32'sd1162288, 32'sd3220770, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2413073, -32'sd456247, 32'sd1159978, -32'sd651813, -32'sd569591, 32'sd915002, 32'sd276516, 32'sd39184, 32'sd2112714, -32'sd8828, 32'sd1414332, -32'sd682888, -32'sd15870, 32'sd850086, 32'sd91746, -32'sd319424, -32'sd1312224, -32'sd163235, -32'sd433188, -32'sd388470, -32'sd944220, 32'sd615266, -32'sd670327, -32'sd419670, 32'sd17224, 32'sd0, 32'sd0, 32'sd484043, 32'sd1795726, -32'sd520561, -32'sd113313, -32'sd3107429, -32'sd1710713, 32'sd2022822, 32'sd515851, 32'sd729904, -32'sd202141, -32'sd1639615, 32'sd250708, 32'sd77481, 32'sd1097811, -32'sd361980, -32'sd383316, -32'sd815686, 32'sd998677, 32'sd967479, 32'sd157357, -32'sd1380580, -32'sd92308, -32'sd852093, -32'sd30943, -32'sd958845, 32'sd1024452, 32'sd1463828, 32'sd0, -32'sd484475, -32'sd314175, -32'sd1811429, 32'sd861909, 32'sd1119899, 32'sd275108, -32'sd903585, -32'sd245719, 32'sd96274, -32'sd2895525, -32'sd1807073, -32'sd1822790, 32'sd542810, 32'sd2456180, 32'sd1328170, 32'sd1257064, 32'sd1141475, -32'sd2308124, -32'sd606778, 32'sd230872, -32'sd1357577, -32'sd1112430, 32'sd620957, 32'sd1975442, -32'sd575806, -32'sd1898363, 32'sd373084, 32'sd0, 32'sd1518391, 32'sd1435949, -32'sd1451053, 32'sd1259523, 32'sd508886, -32'sd632364, 32'sd218599, -32'sd364121, -32'sd1758091, -32'sd1789995, 32'sd1195510, 32'sd235921, 32'sd923585, 32'sd2801756, -32'sd430808, 32'sd216376, -32'sd1197346, -32'sd1087490, 32'sd226239, -32'sd1911380, -32'sd1567858, 32'sd628714, -32'sd548655, 32'sd498906, -32'sd2213261, 32'sd512796, -32'sd323304, 32'sd2170244, 32'sd2032493, -32'sd619372, 32'sd671787, 32'sd1429367, 32'sd1256755, -32'sd1303252, 32'sd1517915, 32'sd287695, 32'sd1372472, -32'sd1335046, -32'sd1348877, -32'sd842220, -32'sd919946, 32'sd1782260, -32'sd1613829, -32'sd4104334, -32'sd2099024, -32'sd1872609, -32'sd2723213, -32'sd2372238, -32'sd2243618, -32'sd750487, -32'sd1189134, -32'sd2743715, -32'sd2422257, 32'sd37125, 32'sd1168137, 32'sd1566854, 32'sd341324, -32'sd624874, -32'sd711472, 32'sd1769394, 32'sd320169, -32'sd428030, -32'sd224417, 32'sd389838, -32'sd46633, -32'sd86679, 32'sd819, -32'sd267184, -32'sd1562623, -32'sd2032146, -32'sd1484491, -32'sd4320884, -32'sd5067666, -32'sd3279951, -32'sd3899208, -32'sd4094874, -32'sd294642, -32'sd919775, -32'sd1411947, -32'sd1162182, -32'sd1203032, 32'sd1617898, -32'sd450175, 32'sd512471, 32'sd1908613, -32'sd1567842, 32'sd999335, 32'sd1133249, 32'sd1264832, 32'sd113936, 32'sd168892, 32'sd886665, -32'sd819373, -32'sd353924, 32'sd403682, 32'sd653809, -32'sd282700, 32'sd1356149, -32'sd2851075, -32'sd6133316, -32'sd2332199, -32'sd749814, -32'sd1090783, -32'sd587980, -32'sd201869, -32'sd87924, 32'sd1307500, 32'sd75401, 32'sd525996, 32'sd1475371, 32'sd1532815, 32'sd959498, 32'sd1150541, -32'sd337851, -32'sd1379292, 32'sd550335, 32'sd500985, 32'sd128702, -32'sd557907, -32'sd781789, -32'sd101444, 32'sd940220, 32'sd3085833, 32'sd1629489, 32'sd1848723, 32'sd2876181, -32'sd423786, -32'sd2734522, -32'sd636678, 32'sd361561, -32'sd282984, 32'sd1783415, 32'sd1211998, 32'sd1703251, 32'sd831867, 32'sd1788320, 32'sd797674, -32'sd875826, -32'sd1436747, 32'sd1537957, 32'sd830564, -32'sd654733, 32'sd932417, -32'sd171700, -32'sd532446, 32'sd1367530, -32'sd841218, -32'sd852749, 32'sd2193987, 32'sd433215, 32'sd2371706, 32'sd1028260, 32'sd4445290, 32'sd4070590, 32'sd16896, -32'sd1900726, 32'sd1001462, 32'sd3358912, 32'sd1083506, 32'sd1197039, 32'sd2713751, 32'sd1994557, 32'sd1523566, -32'sd830845, 32'sd221226, -32'sd485800, 32'sd739907, 32'sd792502, 32'sd742098, 32'sd1586150, 32'sd1566934, -32'sd7968, 32'sd432916, -32'sd1155925, -32'sd2552177, 32'sd461784, 32'sd1369165, -32'sd1481124, 32'sd1583793, 32'sd3190550, 32'sd3908682, 32'sd3446010, -32'sd367461, -32'sd2285755, 32'sd788690, 32'sd370941, 32'sd1649228, 32'sd3130232, 32'sd1589494, 32'sd4097200, 32'sd2249170, -32'sd1726086, -32'sd1439124, 32'sd1435087, 32'sd2335126, 32'sd1484840, 32'sd1436676, 32'sd695379, 32'sd623146, -32'sd1813644, 32'sd2344466, -32'sd1422430, -32'sd826506, -32'sd1025129, -32'sd1883064, -32'sd1654670, -32'sd621291, 32'sd1433554, 32'sd2188764, 32'sd143071, 32'sd1351360, -32'sd175223, 32'sd872081, -32'sd356638, 32'sd894846, 32'sd1561450, 32'sd3818645, 32'sd1392749, 32'sd2587248, -32'sd363458, -32'sd292446, -32'sd5986, -32'sd556043, 32'sd2229575, -32'sd388582, 32'sd492913, 32'sd1327499, -32'sd1740826, -32'sd181347, 32'sd346642, 32'sd20754, -32'sd97130, 32'sd152680, 32'sd1071282, -32'sd717983, 32'sd1566392, -32'sd8339, 32'sd1538496, 32'sd1517217, 32'sd2082733, 32'sd297249, 32'sd1249851, -32'sd187272, 32'sd1519612, 32'sd2761323, 32'sd1111174, -32'sd55308, -32'sd480997, -32'sd526340, -32'sd1540985, -32'sd932908, 32'sd653248, -32'sd114061, 32'sd741319, -32'sd357187, -32'sd981341, -32'sd1123368, -32'sd309772, 32'sd1855319, 32'sd1388198, 32'sd68159, 32'sd352095, -32'sd888872, 32'sd39218, 32'sd2277830, 32'sd2548757, 32'sd1635215, -32'sd624430, -32'sd266101, 32'sd1108036, 32'sd728186, 32'sd865521, 32'sd1244152, 32'sd1058559, -32'sd131497, 32'sd43938, 32'sd696622, -32'sd54489, 32'sd679516, 32'sd600958, -32'sd851663, 32'sd490077, 32'sd1054534, 32'sd239871, 32'sd1199690, 32'sd1526889, 32'sd1103759, 32'sd1100936, -32'sd1085782, -32'sd495872, -32'sd1069389, -32'sd419947, -32'sd399312, 32'sd1811479, -32'sd472344, -32'sd2702298, -32'sd1612160, -32'sd541144, -32'sd1367450, 32'sd14522, 32'sd470196, -32'sd1451939, -32'sd1156915, -32'sd343948, -32'sd893096, 32'sd64932, -32'sd984372, 32'sd0, 32'sd1094988, 32'sd632640, -32'sd877553, 32'sd559348, 32'sd286840, -32'sd2082850, -32'sd1772791, 32'sd904497, -32'sd372872, -32'sd952451, -32'sd782957, -32'sd1574929, 32'sd286091, 32'sd1238359, -32'sd284934, -32'sd1354230, -32'sd961156, 32'sd178310, 32'sd671307, 32'sd488578, 32'sd88054, -32'sd581753, -32'sd2101156, -32'sd1997295, -32'sd1399111, 32'sd1081247, -32'sd461857, -32'sd603976, 32'sd435026, -32'sd281219, -32'sd75266, -32'sd24902, 32'sd295850, -32'sd2183091, -32'sd2657668, -32'sd557170, 32'sd485629, -32'sd2294490, -32'sd1535613, -32'sd1055011, 32'sd1941725, 32'sd923539, -32'sd954787, -32'sd2701041, 32'sd141115, 32'sd733961, 32'sd394484, 32'sd809443, -32'sd1623944, -32'sd2534970, -32'sd3973759, -32'sd2258981, -32'sd33494, 32'sd86967, 32'sd926470, 32'sd969345, -32'sd793181, 32'sd148324, -32'sd893056, 32'sd1091508, -32'sd454566, -32'sd1467309, -32'sd2309900, 32'sd642507, -32'sd809171, -32'sd2339162, -32'sd2193948, -32'sd2078034, 32'sd1157460, 32'sd1029598, 32'sd249955, -32'sd594443, -32'sd1256328, 32'sd952856, -32'sd786059, -32'sd1515395, -32'sd1624338, -32'sd1983140, -32'sd1416233, -32'sd1949929, -32'sd446055, 32'sd1252466, 32'sd931048, 32'sd0, -32'sd256906, -32'sd1098731, 32'sd1315118, 32'sd3388469, 32'sd1193255, -32'sd880999, -32'sd1547312, 32'sd69975, -32'sd924153, -32'sd2342715, -32'sd803712, 32'sd263280, 32'sd164906, 32'sd629646, 32'sd2799337, 32'sd1204542, 32'sd1126213, 32'sd563192, -32'sd1003675, -32'sd1274845, -32'sd1452955, -32'sd3256069, -32'sd1933929, 32'sd222272, 32'sd656790, 32'sd271043, -32'sd244333, 32'sd433019, -32'sd238108, 32'sd935075, -32'sd2584299, -32'sd423310, 32'sd36642, 32'sd1243025, -32'sd1106774, -32'sd1202488, 32'sd1547008, 32'sd240788, 32'sd1098493, 32'sd954966, 32'sd1087307, 32'sd288966, 32'sd1279273, 32'sd3149618, 32'sd2130726, 32'sd246357, 32'sd388274, 32'sd1516202, -32'sd1048172, 32'sd40846, -32'sd936814, -32'sd1142174, -32'sd15236, 32'sd1106265, 32'sd1590531, 32'sd1738743, 32'sd1126685, -32'sd974686, -32'sd1615595, 32'sd319938, -32'sd898999, -32'sd1318427, 32'sd284237, -32'sd1573350, 32'sd440805, -32'sd958220, 32'sd891177, -32'sd211524, 32'sd772661, 32'sd178449, 32'sd133319, 32'sd3326506, -32'sd163416, 32'sd1712763, 32'sd476407, 32'sd500934, -32'sd1153542, -32'sd1615857, -32'sd346460, 32'sd1110822, -32'sd863447, -32'sd123842, 32'sd1382350, 32'sd0, 32'sd1613066, 32'sd1692235, 32'sd367434, 32'sd276717, 32'sd315552, 32'sd868593, -32'sd1588101, -32'sd1851167, -32'sd248692, -32'sd1247180, -32'sd3774273, -32'sd13784, -32'sd430539, 32'sd1898898, -32'sd216498, 32'sd318982, 32'sd407470, 32'sd294538, 32'sd500220, 32'sd1284579, -32'sd229253, -32'sd1763367, -32'sd18717, -32'sd1089541, 32'sd285351, -32'sd54959, 32'sd0, 32'sd0, 32'sd0, -32'sd534733, 32'sd279772, 32'sd1009418, 32'sd1899801, 32'sd856511, -32'sd84604, -32'sd174479, -32'sd755441, 32'sd99682, 32'sd23760, -32'sd1343705, -32'sd358152, -32'sd734777, -32'sd171070, -32'sd1149202, 32'sd997340, 32'sd251820, -32'sd572463, -32'sd268828, -32'sd931849, -32'sd1826826, -32'sd182664, 32'sd416155, 32'sd546685, -32'sd369006, 32'sd0, 32'sd0, 32'sd0, 32'sd1008222, 32'sd2442551, -32'sd702466, -32'sd1262979, 32'sd1722473, 32'sd706353, -32'sd294967, 32'sd101363, 32'sd151284, 32'sd524024, 32'sd963551, -32'sd124352, 32'sd795901, -32'sd1841207, -32'sd308499, 32'sd1906170, 32'sd906916, -32'sd1297311, 32'sd828605, -32'sd969164, 32'sd1262478, 32'sd162159, -32'sd1574935, -32'sd1199424, 32'sd524524, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2354680, -32'sd386846, -32'sd1570430, 32'sd529780, -32'sd931513, -32'sd1369484, 32'sd2764713, 32'sd185630, 32'sd1423349, 32'sd640927, 32'sd1922463, -32'sd205767, -32'sd1113154, 32'sd569303, 32'sd720635, -32'sd10041, 32'sd1398135, -32'sd1124311, 32'sd1588434, 32'sd899581, 32'sd367088, 32'sd434543, 32'sd1800413, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2534512, 32'sd1399827, 32'sd1322783, 32'sd1031824, 32'sd1737123, -32'sd85207, 32'sd69678, 32'sd1417754, 32'sd96594, -32'sd685744, 32'sd566803, 32'sd526723, 32'sd1239773, 32'sd1722862, 32'sd350803, 32'sd1355804, -32'sd435547, 32'sd1802779, 32'sd1611475, 32'sd1442077, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd836875, 32'sd1940371, -32'sd405677, 32'sd1937758, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd346684, -32'sd1474340, 32'sd1055271, 32'sd2098073, -32'sd172863, 32'sd425710, 32'sd1738269, 32'sd142482, 32'sd1107910, -32'sd582973, -32'sd1618006, 32'sd287275, 32'sd704455, 32'sd1091386, 32'sd1079444, 32'sd157739, 32'sd1076964, 32'sd961416, 32'sd1333799, -32'sd72555, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd545326, -32'sd762169, 32'sd381789, 32'sd506484, 32'sd1353955, 32'sd568700, 32'sd2136986, 32'sd601336, -32'sd245662, 32'sd2405492, 32'sd2204703, -32'sd143703, -32'sd465431, 32'sd1371663, -32'sd58435, 32'sd1507666, -32'sd188779, 32'sd81740, -32'sd201104, 32'sd645998, 32'sd276620, -32'sd550458, 32'sd996124, 32'sd1822041, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd697754, 32'sd1330054, 32'sd1711413, 32'sd1977547, 32'sd1924609, 32'sd2092561, 32'sd566537, -32'sd594245, 32'sd986655, 32'sd2064100, 32'sd1032912, 32'sd2067190, -32'sd146948, -32'sd1040453, 32'sd642392, 32'sd342758, -32'sd1641539, -32'sd991960, -32'sd757768, 32'sd1065577, 32'sd684094, 32'sd1565518, 32'sd1646677, 32'sd183529, 32'sd1589158, 32'sd0, 32'sd0, 32'sd738759, -32'sd77015, 32'sd34320, -32'sd211725, 32'sd1302965, 32'sd1789650, 32'sd795732, 32'sd582170, -32'sd407505, 32'sd1874509, 32'sd972038, 32'sd778422, -32'sd733990, 32'sd788881, 32'sd138303, 32'sd1281341, 32'sd826264, 32'sd666373, 32'sd590225, 32'sd650619, -32'sd905410, -32'sd738248, 32'sd128252, 32'sd372302, -32'sd222885, -32'sd412535, 32'sd1095333, 32'sd0, 32'sd872508, 32'sd171107, 32'sd1028578, 32'sd700913, 32'sd529363, 32'sd856155, -32'sd1741461, -32'sd186166, -32'sd1239757, -32'sd39255, -32'sd27961, -32'sd1740315, -32'sd1842653, -32'sd1299877, 32'sd62453, 32'sd218181, 32'sd278494, 32'sd397297, 32'sd2242015, -32'sd105805, -32'sd1816039, -32'sd1471157, -32'sd538140, -32'sd1524337, -32'sd1224604, 32'sd701018, 32'sd1299816, 32'sd0, 32'sd109906, 32'sd254730, 32'sd25149, 32'sd1356221, 32'sd719831, 32'sd564044, -32'sd938791, -32'sd590742, 32'sd1215219, -32'sd1277793, 32'sd367275, -32'sd3619910, -32'sd2825241, -32'sd1445792, -32'sd978553, 32'sd989015, 32'sd1619251, 32'sd1728301, 32'sd1995132, -32'sd343701, -32'sd875265, -32'sd1054278, -32'sd2444818, -32'sd4079209, -32'sd1578440, 32'sd1478147, -32'sd279634, 32'sd1393180, -32'sd246274, 32'sd877328, 32'sd1211398, -32'sd1460443, -32'sd519229, -32'sd793505, 32'sd594699, 32'sd1194208, -32'sd159031, -32'sd698261, -32'sd2476912, -32'sd2633178, -32'sd2097013, 32'sd1279759, -32'sd46510, -32'sd2275577, 32'sd344482, 32'sd1453599, 32'sd1324226, -32'sd389292, 32'sd565130, -32'sd105088, -32'sd604278, 32'sd300045, -32'sd756542, 32'sd193327, -32'sd94848, 32'sd913033, 32'sd1163248, 32'sd1256438, -32'sd12121, -32'sd1085832, -32'sd1069353, 32'sd422772, -32'sd1144093, -32'sd1046265, -32'sd2023526, -32'sd698883, -32'sd476026, 32'sd698021, 32'sd381387, 32'sd1307946, 32'sd1455256, 32'sd888630, -32'sd608459, -32'sd246545, 32'sd619535, -32'sd478793, -32'sd961047, 32'sd50243, 32'sd697040, -32'sd636912, -32'sd809920, 32'sd1646366, -32'sd298489, 32'sd739884, -32'sd1523131, -32'sd84960, -32'sd964089, 32'sd781746, 32'sd1190019, -32'sd146928, -32'sd465682, -32'sd1113964, -32'sd1713688, -32'sd2154796, -32'sd1277741, 32'sd425784, 32'sd2649335, -32'sd128943, -32'sd946807, -32'sd1606511, -32'sd225218, -32'sd861792, -32'sd590075, -32'sd22505, -32'sd1079449, 32'sd1487739, 32'sd1370888, 32'sd756243, -32'sd1616621, 32'sd1568120, -32'sd620551, -32'sd208607, -32'sd217925, 32'sd348409, -32'sd1047571, 32'sd312284, 32'sd2244763, -32'sd326515, -32'sd2337421, -32'sd1273976, -32'sd786150, -32'sd1741396, -32'sd1621016, 32'sd2398947, -32'sd282321, -32'sd879155, -32'sd1945532, -32'sd2452763, -32'sd1729496, -32'sd1191174, -32'sd1310717, -32'sd120074, 32'sd348474, 32'sd356537, 32'sd1665181, -32'sd132326, -32'sd749635, 32'sd1071973, 32'sd303359, -32'sd935662, 32'sd1070754, 32'sd310549, -32'sd1331981, -32'sd1471755, 32'sd394366, 32'sd18742, -32'sd735169, 32'sd464299, 32'sd1793711, -32'sd2095587, 32'sd1291457, -32'sd364484, -32'sd870497, -32'sd2856925, -32'sd4036760, -32'sd3609974, -32'sd1050810, -32'sd1835782, -32'sd1827392, 32'sd1944465, 32'sd1058752, 32'sd1381995, -32'sd77522, 32'sd514880, 32'sd312877, 32'sd448773, 32'sd1385093, 32'sd988526, 32'sd802835, -32'sd1282799, -32'sd757563, 32'sd1295023, 32'sd616838, 32'sd145386, -32'sd486245, -32'sd677422, 32'sd825281, 32'sd373665, 32'sd142215, 32'sd229230, -32'sd784217, -32'sd751523, -32'sd174596, 32'sd163733, 32'sd995877, 32'sd1773485, -32'sd137520, 32'sd932631, 32'sd1929662, 32'sd725854, 32'sd2081306, 32'sd501442, -32'sd84102, -32'sd323195, 32'sd251457, 32'sd910662, -32'sd888840, -32'sd1271901, -32'sd879480, 32'sd755297, 32'sd1186707, -32'sd1052989, 32'sd560948, -32'sd543341, 32'sd1820935, -32'sd638681, 32'sd922624, -32'sd1586226, -32'sd175827, 32'sd2053194, 32'sd1866654, 32'sd3294458, 32'sd561836, 32'sd1678963, -32'sd129179, 32'sd1218092, 32'sd753025, 32'sd2822304, 32'sd1293284, -32'sd503613, 32'sd214286, 32'sd363610, 32'sd970665, 32'sd493714, 32'sd334067, -32'sd348774, -32'sd1588716, -32'sd14036, 32'sd1849018, -32'sd111062, 32'sd1582213, 32'sd942330, 32'sd1513924, 32'sd1377701, -32'sd219892, -32'sd1422505, -32'sd881224, -32'sd439381, 32'sd3581875, 32'sd2626076, 32'sd1461737, -32'sd544156, -32'sd1117847, -32'sd303696, 32'sd299327, -32'sd127535, 32'sd1140604, -32'sd1099702, 32'sd4792, 32'sd19138, 32'sd1273199, -32'sd400538, 32'sd404313, 32'sd1011686, -32'sd1672353, -32'sd2061439, 32'sd697988, 32'sd1521425, 32'sd581602, 32'sd948395, 32'sd2593755, -32'sd138128, -32'sd921576, -32'sd1117068, -32'sd958871, 32'sd2024718, 32'sd2760059, 32'sd1756982, -32'sd907293, 32'sd10286, 32'sd175917, -32'sd228537, 32'sd915069, -32'sd134616, 32'sd1003340, 32'sd776311, -32'sd1165281, 32'sd872554, 32'sd488598, 32'sd641246, 32'sd1841496, 32'sd936829, -32'sd1624942, -32'sd854387, 32'sd1092055, -32'sd481099, -32'sd388423, 32'sd294504, 32'sd1797490, 32'sd1147261, 32'sd2710758, 32'sd3095535, 32'sd1627051, 32'sd1545873, 32'sd713861, -32'sd556530, -32'sd2232900, -32'sd966897, -32'sd1803252, -32'sd1166819, -32'sd2160877, -32'sd2030805, -32'sd62984, -32'sd1092221, 32'sd688595, -32'sd421003, -32'sd165049, 32'sd0, -32'sd51755, 32'sd737732, 32'sd758997, -32'sd67585, 32'sd2028540, 32'sd1249749, -32'sd1209455, -32'sd635445, -32'sd1136344, 32'sd1765041, 32'sd908588, 32'sd1044420, -32'sd663175, -32'sd733728, 32'sd1117271, 32'sd20550, -32'sd1786827, 32'sd863192, -32'sd856560, -32'sd1183989, -32'sd75706, -32'sd415715, 32'sd502041, -32'sd897705, 32'sd1529967, -32'sd1133291, 32'sd886015, 32'sd755459, 32'sd1585962, -32'sd608324, 32'sd8086, 32'sd539211, -32'sd26280, 32'sd697449, -32'sd65141, 32'sd295796, 32'sd744897, 32'sd2105135, 32'sd2054617, 32'sd655087, 32'sd1070403, -32'sd746301, 32'sd162456, -32'sd909582, 32'sd156016, 32'sd1254575, 32'sd122035, -32'sd212135, -32'sd847706, 32'sd635953, -32'sd248657, -32'sd2430866, 32'sd362838, -32'sd1353702, -32'sd383118, 32'sd821858, -32'sd809015, 32'sd662425, 32'sd574231, -32'sd967759, 32'sd1870242, -32'sd764394, 32'sd483768, -32'sd847719, 32'sd935419, 32'sd1862889, 32'sd2042176, 32'sd1338985, 32'sd21721, -32'sd115116, 32'sd258136, 32'sd247239, 32'sd1164871, 32'sd1671837, 32'sd965616, 32'sd414127, 32'sd272340, -32'sd1435089, -32'sd1048070, 32'sd621370, -32'sd726550, 32'sd1641077, -32'sd663014, 32'sd0, 32'sd336960, -32'sd428958, 32'sd1186626, -32'sd113656, 32'sd1192275, -32'sd210805, 32'sd459646, -32'sd104464, 32'sd1903437, -32'sd149851, 32'sd29584, -32'sd354025, 32'sd1200260, 32'sd2008219, 32'sd2656828, 32'sd1430843, 32'sd1126442, 32'sd2929452, 32'sd1772770, 32'sd228926, -32'sd1389598, -32'sd2420568, -32'sd3226142, -32'sd838390, -32'sd878159, 32'sd664232, 32'sd925968, 32'sd1739317, 32'sd1610084, -32'sd262558, 32'sd586283, 32'sd1361745, -32'sd385303, -32'sd1242585, -32'sd396936, 32'sd1218993, -32'sd416636, 32'sd195184, -32'sd152775, 32'sd1937312, 32'sd2215903, 32'sd2450097, 32'sd868510, 32'sd807003, 32'sd544316, 32'sd1700164, 32'sd101526, -32'sd1502085, -32'sd2008253, -32'sd1550334, -32'sd1649032, -32'sd1407422, 32'sd1130185, 32'sd193235, 32'sd575812, 32'sd1789255, 32'sd1466426, 32'sd676879, -32'sd347128, 32'sd2106456, -32'sd665975, -32'sd610350, -32'sd1111590, -32'sd891716, -32'sd123997, 32'sd879940, -32'sd216720, -32'sd1230217, -32'sd1450710, -32'sd667736, 32'sd3171446, -32'sd251886, 32'sd277481, -32'sd1832508, -32'sd1826259, -32'sd1640090, -32'sd2316519, -32'sd2953410, -32'sd1941821, -32'sd924541, 32'sd485916, 32'sd118238, -32'sd809372, 32'sd0, 32'sd814832, 32'sd957641, -32'sd1213728, -32'sd594787, -32'sd408501, -32'sd565394, 32'sd256174, -32'sd1539962, 32'sd997914, -32'sd577859, -32'sd1926261, 32'sd337224, -32'sd60442, 32'sd136969, 32'sd1431282, 32'sd1030918, 32'sd118768, -32'sd550311, 32'sd182144, -32'sd144200, -32'sd1169245, -32'sd290198, -32'sd1168297, -32'sd769370, -32'sd500407, -32'sd422960, 32'sd0, 32'sd0, 32'sd0, 32'sd288747, -32'sd1076947, 32'sd1333900, -32'sd1182306, -32'sd912038, -32'sd1487631, 32'sd1320456, 32'sd367934, -32'sd516509, -32'sd1726375, 32'sd989903, -32'sd768396, 32'sd1260183, 32'sd439865, -32'sd17429, -32'sd384387, -32'sd17980, -32'sd381788, -32'sd1752777, -32'sd1995318, -32'sd1188992, -32'sd23252, 32'sd760849, 32'sd656106, 32'sd953690, 32'sd0, 32'sd0, 32'sd0, -32'sd400763, -32'sd33164, 32'sd514685, -32'sd1197543, -32'sd431111, 32'sd749470, -32'sd113315, 32'sd708352, -32'sd858812, -32'sd115307, -32'sd133857, 32'sd2263559, 32'sd486930, 32'sd432242, 32'sd1798230, 32'sd1047587, -32'sd1644859, -32'sd1388612, 32'sd1432971, 32'sd534289, -32'sd751920, -32'sd1531419, -32'sd789352, 32'sd931117, 32'sd304922, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd892981, -32'sd252335, -32'sd190283, -32'sd532966, 32'sd416826, 32'sd986575, -32'sd510930, -32'sd70269, 32'sd275558, 32'sd83276, 32'sd278386, -32'sd563372, 32'sd582606, 32'sd1704084, -32'sd73165, -32'sd48477, 32'sd1250717, 32'sd2176699, -32'sd81467, -32'sd1101402, 32'sd537830, 32'sd944779, -32'sd221393, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2001787, 32'sd48885, 32'sd835286, 32'sd1456525, -32'sd212980, 32'sd1547028, 32'sd1035502, 32'sd405818, 32'sd2046243, 32'sd216186, 32'sd1350939, -32'sd1337715, 32'sd342422, 32'sd401169, 32'sd732156, 32'sd869945, 32'sd791854, 32'sd1432243, -32'sd1243228, 32'sd1124714, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd179957, -32'sd673982, -32'sd432104, -32'sd848767, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd99699, -32'sd1031803, -32'sd725531, -32'sd242688, -32'sd1030100, -32'sd493113, -32'sd279596, 32'sd807244, 32'sd133860, -32'sd167539, -32'sd877333, -32'sd621671, -32'sd1765229, -32'sd1632598, -32'sd1304547, -32'sd262360, -32'sd1350346, -32'sd1256776, -32'sd895347, -32'sd231230, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd689624, -32'sd1009323, 32'sd1223185, 32'sd320622, -32'sd1412232, -32'sd86274, 32'sd101269, -32'sd552329, -32'sd87139, -32'sd1100745, -32'sd1860899, -32'sd1330339, -32'sd1516685, -32'sd363394, -32'sd320534, -32'sd444115, 32'sd1258142, 32'sd217414, 32'sd232106, -32'sd839199, -32'sd128048, 32'sd1089707, 32'sd265032, -32'sd767264, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd310280, -32'sd1055470, 32'sd446456, 32'sd644748, -32'sd1856928, -32'sd1420455, -32'sd929549, -32'sd294309, -32'sd861297, -32'sd1616988, -32'sd2611989, -32'sd2989057, -32'sd2041599, 32'sd515219, -32'sd667893, -32'sd571743, 32'sd1465050, 32'sd1065918, -32'sd413899, 32'sd1174894, 32'sd1203379, -32'sd1052432, 32'sd697801, 32'sd999161, -32'sd177995, 32'sd0, 32'sd0, -32'sd667059, 32'sd336175, -32'sd2397247, -32'sd437826, -32'sd1345011, -32'sd95004, -32'sd1934031, -32'sd1068453, -32'sd1040768, -32'sd911588, -32'sd457907, 32'sd576465, -32'sd1648149, -32'sd165796, -32'sd372488, 32'sd1539771, 32'sd985002, 32'sd528277, -32'sd2181086, -32'sd1364975, 32'sd37738, 32'sd102649, -32'sd516839, 32'sd1256815, 32'sd502000, 32'sd1105439, -32'sd1465341, 32'sd0, 32'sd98870, -32'sd761077, -32'sd801836, -32'sd313488, -32'sd551067, -32'sd770295, -32'sd1590939, -32'sd349716, -32'sd1169102, -32'sd244610, 32'sd495889, 32'sd1470132, 32'sd1097024, 32'sd1616031, 32'sd134644, 32'sd903852, 32'sd107837, -32'sd640653, -32'sd1804157, -32'sd1372556, 32'sd572566, 32'sd758929, -32'sd1488771, -32'sd1704964, -32'sd106726, 32'sd269169, 32'sd783225, 32'sd0, 32'sd642113, -32'sd1465337, 32'sd868730, -32'sd2026492, 32'sd1733703, 32'sd278678, -32'sd1223180, -32'sd1215097, 32'sd317847, 32'sd2094894, 32'sd612468, -32'sd635066, -32'sd2297633, 32'sd18188, -32'sd3248566, -32'sd2543680, -32'sd3094925, -32'sd105980, -32'sd553824, -32'sd201786, -32'sd1506051, -32'sd757448, 32'sd1294073, -32'sd366469, -32'sd410753, -32'sd788806, 32'sd607125, -32'sd884901, 32'sd1011785, -32'sd200031, -32'sd1193928, -32'sd2112961, -32'sd578832, -32'sd1055176, -32'sd1666319, 32'sd194580, 32'sd464647, 32'sd1553651, -32'sd1817639, -32'sd2224084, -32'sd493642, -32'sd2654173, -32'sd337560, 32'sd24891, -32'sd802400, 32'sd740469, 32'sd2200069, 32'sd1555286, 32'sd554556, 32'sd2643353, 32'sd39708, -32'sd207112, 32'sd405121, 32'sd1073087, -32'sd686173, -32'sd373915, 32'sd262438, 32'sd657478, -32'sd1352409, -32'sd1234158, -32'sd1445368, -32'sd265946, 32'sd516211, 32'sd2378619, 32'sd162304, -32'sd482006, -32'sd1313536, -32'sd1036963, -32'sd998605, 32'sd2148574, 32'sd961278, 32'sd1523018, 32'sd1182934, 32'sd1134117, 32'sd658745, 32'sd2655402, 32'sd2114940, 32'sd975832, 32'sd385352, 32'sd979840, -32'sd1643536, 32'sd384198, -32'sd1460679, -32'sd1022156, -32'sd64489, -32'sd896802, -32'sd1564784, -32'sd255272, 32'sd945607, -32'sd530624, 32'sd727562, 32'sd1306903, 32'sd863198, -32'sd430503, -32'sd851572, 32'sd763045, 32'sd1250892, 32'sd656834, 32'sd2251447, 32'sd2458448, 32'sd297315, 32'sd223108, 32'sd937888, -32'sd665047, 32'sd396094, 32'sd1651756, 32'sd1510287, -32'sd1075728, -32'sd292073, -32'sd426090, -32'sd1310951, -32'sd969540, -32'sd1349203, -32'sd1467848, -32'sd2274998, -32'sd117304, 32'sd309248, -32'sd195098, 32'sd1209136, 32'sd1781601, -32'sd284803, 32'sd517369, -32'sd2684020, 32'sd283012, -32'sd1840013, -32'sd899145, -32'sd295648, -32'sd455850, 32'sd753489, -32'sd390399, 32'sd339923, -32'sd461531, -32'sd946789, 32'sd1795837, 32'sd326327, 32'sd1058545, 32'sd1996637, 32'sd75787, 32'sd1043460, -32'sd166026, -32'sd131755, -32'sd1390848, -32'sd2160286, -32'sd151530, 32'sd1200365, 32'sd1032214, 32'sd744910, -32'sd533557, 32'sd3803048, 32'sd3069189, -32'sd148238, -32'sd1195904, -32'sd3261153, -32'sd2895185, -32'sd2368607, -32'sd20136, 32'sd201171, -32'sd1288483, 32'sd59297, -32'sd1474165, 32'sd740687, 32'sd2195987, 32'sd750541, 32'sd859220, 32'sd583109, 32'sd2933111, -32'sd569075, 32'sd463747, 32'sd767530, -32'sd716226, -32'sd15705, 32'sd393693, 32'sd1283108, -32'sd354401, 32'sd1685274, 32'sd3667294, 32'sd5159523, 32'sd3439789, 32'sd2409798, -32'sd133017, -32'sd1056151, -32'sd3131642, -32'sd2298406, -32'sd886859, 32'sd1951563, -32'sd722083, 32'sd125714, -32'sd525122, -32'sd293578, 32'sd868583, 32'sd2909603, 32'sd1058747, 32'sd737949, 32'sd1740159, 32'sd858580, -32'sd599967, 32'sd2001451, 32'sd1061283, -32'sd1863327, -32'sd1050469, -32'sd2019958, -32'sd2807824, -32'sd832079, 32'sd931134, 32'sd4729048, 32'sd3278970, 32'sd3100749, 32'sd2028710, 32'sd3521837, 32'sd1349461, 32'sd412859, 32'sd1271080, -32'sd251152, 32'sd128727, -32'sd130832, 32'sd168045, 32'sd286398, 32'sd1404199, 32'sd793928, -32'sd1241033, 32'sd1115820, 32'sd648590, 32'sd505112, -32'sd364392, 32'sd953575, -32'sd885538, -32'sd12692, -32'sd803731, -32'sd439169, -32'sd2619216, -32'sd2220626, -32'sd221569, 32'sd240151, 32'sd2998701, 32'sd2593971, 32'sd3626505, 32'sd3377154, 32'sd1749368, -32'sd2218923, -32'sd2065298, 32'sd1060767, -32'sd1628987, -32'sd88102, -32'sd94937, 32'sd557128, -32'sd176807, -32'sd778866, -32'sd1291491, 32'sd1149255, 32'sd528944, -32'sd934407, 32'sd1419985, -32'sd282326, -32'sd1471808, 32'sd1032106, -32'sd1182023, -32'sd1431109, -32'sd3786135, -32'sd4644697, -32'sd3545262, -32'sd1040358, 32'sd2201183, 32'sd1810707, 32'sd983848, 32'sd1555692, 32'sd1994679, 32'sd343444, -32'sd210657, -32'sd457381, -32'sd398482, -32'sd449018, -32'sd1178177, -32'sd838630, -32'sd3350984, -32'sd123375, -32'sd3780639, -32'sd2026431, -32'sd2765611, -32'sd394501, 32'sd83330, -32'sd1424670, -32'sd2504564, 32'sd2744486, 32'sd204317, -32'sd2520193, -32'sd5507198, -32'sd4504669, -32'sd4599798, -32'sd2312205, -32'sd2642672, -32'sd3348232, -32'sd1126908, 32'sd899551, 32'sd224185, 32'sd907916, -32'sd985186, -32'sd394554, -32'sd1877630, -32'sd2529176, -32'sd3172013, -32'sd3236217, -32'sd1519986, -32'sd1250324, -32'sd3520702, -32'sd2577786, 32'sd394662, -32'sd564582, 32'sd0, 32'sd643333, -32'sd1168391, -32'sd148830, 32'sd1228500, -32'sd280331, -32'sd1619203, -32'sd3028176, -32'sd5822823, -32'sd2632991, -32'sd5044955, -32'sd3575155, -32'sd2103127, 32'sd1500277, -32'sd332703, -32'sd1032697, -32'sd1623409, -32'sd816646, 32'sd158737, -32'sd2111263, -32'sd990662, -32'sd2833968, -32'sd2302619, -32'sd1330602, -32'sd2771270, 32'sd502444, 32'sd910157, 32'sd15666, 32'sd12405, 32'sd843552, 32'sd118697, -32'sd7353, 32'sd1898503, 32'sd2034280, -32'sd545868, -32'sd1371649, -32'sd859376, -32'sd2979481, -32'sd1544643, -32'sd1343443, -32'sd1312262, 32'sd886181, 32'sd292948, 32'sd801442, -32'sd1201521, -32'sd87942, -32'sd1399725, -32'sd608213, 32'sd264246, -32'sd808009, -32'sd1156900, -32'sd1173269, -32'sd2039113, 32'sd876846, 32'sd925578, -32'sd387818, -32'sd658115, -32'sd389348, 32'sd90574, -32'sd1203452, -32'sd852271, 32'sd356179, -32'sd843130, 32'sd1238110, 32'sd2880431, -32'sd245696, 32'sd814281, -32'sd2751913, -32'sd348373, 32'sd1540090, 32'sd2044169, 32'sd665084, -32'sd190648, -32'sd1858318, 32'sd674771, 32'sd130077, 32'sd1157116, -32'sd2073267, -32'sd198129, -32'sd2664568, -32'sd868035, 32'sd479648, -32'sd1160980, 32'sd130292, 32'sd0, -32'sd100044, 32'sd57417, 32'sd755403, -32'sd1965684, -32'sd1112510, -32'sd752729, 32'sd1750096, 32'sd1244227, 32'sd1921036, 32'sd331597, -32'sd272632, -32'sd832569, 32'sd976189, -32'sd1520672, -32'sd247298, -32'sd1327736, -32'sd529130, 32'sd105004, -32'sd315012, 32'sd372871, -32'sd1949866, -32'sd572157, -32'sd1684217, -32'sd1108110, -32'sd463494, 32'sd124466, -32'sd215394, -32'sd907127, -32'sd1444380, -32'sd1134688, -32'sd1873893, -32'sd354655, -32'sd66700, -32'sd250224, 32'sd603597, 32'sd1183589, 32'sd2679785, 32'sd1227674, 32'sd1673405, -32'sd167111, 32'sd575343, -32'sd1182768, 32'sd381910, -32'sd486112, 32'sd1012626, 32'sd1683753, -32'sd2103545, -32'sd413209, -32'sd1414311, 32'sd896700, -32'sd1435723, -32'sd2008448, -32'sd1069472, -32'sd930859, 32'sd179762, -32'sd503458, 32'sd301089, -32'sd343609, -32'sd880628, -32'sd190920, -32'sd1699856, -32'sd379498, 32'sd2024024, 32'sd1440155, 32'sd758377, 32'sd465325, 32'sd267823, 32'sd161708, 32'sd908273, 32'sd2902008, 32'sd1957238, -32'sd73821, 32'sd2183172, -32'sd583650, -32'sd881765, -32'sd2300144, -32'sd1273963, -32'sd1088145, 32'sd682243, -32'sd688987, -32'sd569473, -32'sd275166, -32'sd750664, 32'sd0, -32'sd785833, -32'sd445646, -32'sd1011182, -32'sd596933, 32'sd1193001, -32'sd827303, 32'sd779871, 32'sd497640, 32'sd74323, -32'sd848198, 32'sd1497547, 32'sd1164450, 32'sd791586, -32'sd133187, 32'sd1251692, 32'sd99824, 32'sd1705486, -32'sd955035, -32'sd1100495, 32'sd1112626, -32'sd1533365, -32'sd1629552, 32'sd1271094, 32'sd481428, -32'sd2504306, -32'sd1294966, 32'sd0, 32'sd0, 32'sd0, -32'sd17962, 32'sd197086, -32'sd960951, -32'sd122951, -32'sd954595, 32'sd194089, -32'sd1249809, -32'sd3128416, -32'sd449037, 32'sd672966, -32'sd967975, 32'sd1256814, 32'sd94790, 32'sd600934, -32'sd298098, -32'sd1322956, 32'sd2025801, 32'sd2262581, 32'sd88364, -32'sd797543, -32'sd1703084, 32'sd1301726, -32'sd596041, -32'sd1127042, -32'sd975876, 32'sd0, 32'sd0, 32'sd0, -32'sd527735, -32'sd279294, -32'sd520677, 32'sd826061, 32'sd113070, -32'sd807659, -32'sd34282, -32'sd1399997, -32'sd466927, -32'sd373570, -32'sd461398, 32'sd929701, 32'sd900990, 32'sd180404, 32'sd429642, 32'sd1172141, 32'sd508837, 32'sd1600252, 32'sd591875, -32'sd417229, 32'sd352660, -32'sd73239, -32'sd816729, 32'sd172730, -32'sd135703, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd909443, 32'sd746041, 32'sd79617, 32'sd2045486, -32'sd670715, 32'sd2480023, -32'sd135840, -32'sd116742, -32'sd58362, 32'sd1462319, -32'sd1054996, 32'sd2193976, 32'sd1926547, 32'sd1323362, 32'sd793999, 32'sd1196391, -32'sd394261, -32'sd1267544, 32'sd472385, -32'sd102399, 32'sd620413, 32'sd795873, -32'sd709681, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd781363, -32'sd241571, -32'sd1680959, 32'sd1029144, -32'sd403166, 32'sd315069, 32'sd625934, -32'sd227843, 32'sd1001712, 32'sd997838, -32'sd802660, 32'sd566123, 32'sd90318, 32'sd325418, 32'sd525055, 32'sd502724, 32'sd551053, -32'sd200908, -32'sd607777, -32'sd265539, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd957511, -32'sd134910, -32'sd587774, -32'sd1202374, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1369841, -32'sd925727, -32'sd987468, -32'sd1400240, -32'sd1593552, -32'sd2182827, -32'sd1129807, 32'sd293231, -32'sd1149332, -32'sd615413, -32'sd1328683, -32'sd1829154, -32'sd867963, -32'sd1938161, -32'sd2044416, -32'sd1981456, -32'sd1410061, -32'sd715916, 32'sd213752, 32'sd649116, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1219426, -32'sd971796, -32'sd1533099, 32'sd915844, 32'sd1654566, -32'sd257129, 32'sd830853, -32'sd1780021, -32'sd262936, -32'sd872294, -32'sd613567, -32'sd1383053, -32'sd565818, -32'sd732767, -32'sd852936, -32'sd1601580, -32'sd1086668, -32'sd1820719, -32'sd2198759, -32'sd2094023, -32'sd715274, 32'sd541052, -32'sd391992, -32'sd1782884, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1531351, -32'sd393740, -32'sd1386658, -32'sd987812, -32'sd545143, 32'sd1777136, 32'sd135034, -32'sd1234306, -32'sd77045, -32'sd955561, -32'sd623643, 32'sd1359377, 32'sd3379136, -32'sd265608, 32'sd105417, -32'sd478994, -32'sd821445, -32'sd4148862, -32'sd2234251, -32'sd49780, 32'sd634601, 32'sd878924, -32'sd719989, -32'sd975708, -32'sd1466268, 32'sd0, 32'sd0, 32'sd339164, -32'sd225722, -32'sd441270, 32'sd1877302, 32'sd1432102, 32'sd1669640, 32'sd163019, 32'sd416566, -32'sd1229459, -32'sd68814, -32'sd614334, 32'sd2208909, 32'sd3067577, 32'sd111363, 32'sd494833, -32'sd756344, 32'sd1262956, -32'sd1316346, -32'sd1744639, -32'sd2983318, -32'sd2365342, 32'sd900493, -32'sd1252962, 32'sd251309, -32'sd274737, -32'sd740786, -32'sd727955, 32'sd0, -32'sd1103396, 32'sd457839, -32'sd1874685, -32'sd469870, 32'sd390543, -32'sd857755, -32'sd2220307, -32'sd2238252, -32'sd1922070, -32'sd1100225, 32'sd194485, 32'sd1372633, 32'sd214635, 32'sd1014995, 32'sd3597856, 32'sd3733243, 32'sd243549, 32'sd1345571, 32'sd2500130, -32'sd2046185, -32'sd1616502, -32'sd812721, 32'sd898146, 32'sd377131, 32'sd689127, 32'sd896395, -32'sd1635305, 32'sd0, 32'sd878793, 32'sd177071, -32'sd1103188, -32'sd733543, -32'sd572092, -32'sd940089, -32'sd2174865, -32'sd615845, 32'sd1116508, 32'sd912463, 32'sd869774, 32'sd1863995, 32'sd2085752, 32'sd3099593, 32'sd2818840, 32'sd1435241, 32'sd2308056, 32'sd1196547, -32'sd1009591, -32'sd930321, -32'sd966698, 32'sd1613445, 32'sd354111, 32'sd1044914, -32'sd977152, 32'sd1116704, 32'sd608141, -32'sd431185, -32'sd865212, -32'sd1135071, -32'sd8319, -32'sd1982267, 32'sd938659, -32'sd254746, 32'sd256034, -32'sd1342829, 32'sd1036552, 32'sd1973344, 32'sd1114743, 32'sd2117000, -32'sd60673, -32'sd811499, -32'sd1233516, -32'sd517606, 32'sd397942, -32'sd1002847, -32'sd818103, -32'sd1794695, -32'sd2778219, 32'sd51264, 32'sd161316, 32'sd711697, -32'sd1841854, -32'sd898106, -32'sd703411, -32'sd1558506, -32'sd1200110, 32'sd698697, 32'sd1025811, 32'sd482675, 32'sd224182, 32'sd832740, 32'sd493559, 32'sd2419724, 32'sd2969237, 32'sd230942, 32'sd452039, -32'sd336697, -32'sd3488291, -32'sd2217311, -32'sd1034999, 32'sd391388, 32'sd1581876, 32'sd3519390, 32'sd1455019, -32'sd585302, -32'sd753965, -32'sd136246, 32'sd242425, -32'sd669456, 32'sd432500, -32'sd305348, 32'sd149454, -32'sd469629, -32'sd2216831, -32'sd326757, -32'sd490839, 32'sd452959, -32'sd38484, 32'sd1284094, 32'sd1837746, 32'sd2791169, 32'sd1248890, 32'sd951130, -32'sd611629, -32'sd3409160, -32'sd2545721, -32'sd3859004, 32'sd909639, 32'sd2740838, 32'sd5733443, 32'sd3127209, 32'sd3263244, 32'sd1032008, 32'sd621123, -32'sd203579, -32'sd1036907, -32'sd3336082, -32'sd904601, 32'sd434104, 32'sd1055952, -32'sd1021114, -32'sd442799, -32'sd940015, 32'sd1130608, -32'sd489991, 32'sd1389103, -32'sd512428, 32'sd666016, -32'sd34345, 32'sd840106, -32'sd2339531, -32'sd1916228, -32'sd4997096, -32'sd3984653, -32'sd1877767, 32'sd164823, 32'sd2927967, 32'sd3419803, 32'sd1715793, 32'sd3409324, 32'sd1999708, 32'sd888163, 32'sd1127019, -32'sd1650326, -32'sd2934578, 32'sd726109, -32'sd234127, 32'sd1067264, -32'sd1032015, -32'sd2099897, -32'sd22498, -32'sd1109685, -32'sd202940, 32'sd1173945, -32'sd731987, -32'sd222301, 32'sd901782, -32'sd176906, -32'sd560475, -32'sd4086388, -32'sd3344133, -32'sd1740594, 32'sd1200528, 32'sd1914177, 32'sd2146398, 32'sd2535610, 32'sd2620319, 32'sd3705375, 32'sd2484917, -32'sd165786, 32'sd902744, 32'sd528320, -32'sd2884251, -32'sd1682339, -32'sd1169424, -32'sd1721773, -32'sd1115431, -32'sd573171, 32'sd814042, -32'sd977932, 32'sd735359, 32'sd667869, -32'sd1849343, 32'sd286904, -32'sd283954, -32'sd484021, -32'sd910558, -32'sd1273239, -32'sd387492, 32'sd268331, 32'sd621023, 32'sd783227, -32'sd87120, -32'sd1059793, 32'sd2002122, 32'sd804339, 32'sd523236, 32'sd1271195, 32'sd414918, 32'sd1958473, -32'sd1381834, -32'sd1925714, 32'sd2163699, -32'sd322326, -32'sd933744, -32'sd1844666, -32'sd1058183, 32'sd1446475, 32'sd187409, 32'sd291206, -32'sd1565350, -32'sd642637, -32'sd570486, -32'sd2336253, -32'sd798855, 32'sd286914, 32'sd1726008, 32'sd2263652, 32'sd120508, 32'sd543233, 32'sd403958, -32'sd1085821, 32'sd1982462, 32'sd1624867, 32'sd1888122, 32'sd2191385, 32'sd1089130, 32'sd988997, -32'sd432859, 32'sd1029462, 32'sd1090416, -32'sd1673834, -32'sd564380, -32'sd1393028, 32'sd207163, -32'sd524676, -32'sd928628, -32'sd1400321, -32'sd2681923, -32'sd703676, 32'sd1029408, 32'sd457077, 32'sd1461926, -32'sd653439, 32'sd1505259, -32'sd538816, 32'sd578702, -32'sd1514891, -32'sd218212, 32'sd2010076, -32'sd119662, 32'sd1346421, 32'sd3183515, 32'sd5705601, 32'sd2230424, 32'sd33446, -32'sd1139605, 32'sd856284, -32'sd4075, -32'sd1008757, -32'sd439854, 32'sd990604, -32'sd149474, -32'sd163413, -32'sd689326, 32'sd852686, -32'sd757089, 32'sd25362, 32'sd452339, -32'sd86068, -32'sd306736, 32'sd1014820, 32'sd881427, -32'sd873245, -32'sd1302548, -32'sd2619843, -32'sd1699848, 32'sd1063075, -32'sd1350147, 32'sd2362989, 32'sd2089412, 32'sd3287761, 32'sd535656, -32'sd1080647, -32'sd2450470, 32'sd682441, 32'sd206366, -32'sd1307778, 32'sd266179, 32'sd1024941, 32'sd121794, -32'sd1026385, 32'sd54065, 32'sd1559763, -32'sd2244035, -32'sd605094, -32'sd3711977, -32'sd1204047, 32'sd1387949, 32'sd1278016, 32'sd1656512, 32'sd49303, -32'sd211137, -32'sd3591101, 32'sd4831, 32'sd1863986, -32'sd665680, 32'sd2251481, 32'sd2300194, 32'sd531036, 32'sd108822, -32'sd1363000, -32'sd40330, -32'sd349305, 32'sd1545983, -32'sd1384422, 32'sd0, -32'sd1154536, -32'sd313979, -32'sd255438, 32'sd667562, 32'sd792635, -32'sd2997531, -32'sd2965945, -32'sd2587673, 32'sd582086, 32'sd1934393, -32'sd1954250, -32'sd1384445, 32'sd690286, -32'sd62878, -32'sd545172, 32'sd1733756, 32'sd1637358, 32'sd901316, 32'sd431381, -32'sd1192424, -32'sd487749, -32'sd1824325, -32'sd2571938, -32'sd239377, -32'sd303751, -32'sd1127116, -32'sd1628398, -32'sd1275000, 32'sd719845, 32'sd1939384, 32'sd700849, -32'sd2298122, 32'sd1983233, -32'sd110252, -32'sd2915020, -32'sd144580, -32'sd1120764, -32'sd229660, 32'sd147347, -32'sd789099, -32'sd1979181, -32'sd968186, 32'sd1328100, 32'sd2129790, 32'sd1972748, 32'sd267605, 32'sd1415352, -32'sd1278074, 32'sd383333, 32'sd25098, -32'sd446688, -32'sd1385970, 32'sd239107, -32'sd1467169, -32'sd1716910, 32'sd714185, -32'sd839601, -32'sd144104, 32'sd1579482, -32'sd1201649, 32'sd2167818, 32'sd292417, 32'sd1116249, 32'sd427779, 32'sd1201520, -32'sd502894, -32'sd1224930, -32'sd903099, -32'sd2327964, 32'sd262937, 32'sd2546939, 32'sd1967380, -32'sd1825009, 32'sd1401134, -32'sd720131, -32'sd1499364, -32'sd821864, -32'sd1640510, -32'sd835092, -32'sd1167161, 32'sd1229788, 32'sd155631, -32'sd651933, 32'sd0, 32'sd312771, 32'sd1099819, 32'sd596406, -32'sd419169, 32'sd1436414, -32'sd459866, 32'sd494100, 32'sd513156, 32'sd13289, -32'sd475660, -32'sd1266281, 32'sd1138920, -32'sd1787727, -32'sd540237, 32'sd438788, 32'sd342560, 32'sd1506362, -32'sd431099, -32'sd400862, 32'sd571788, -32'sd457116, -32'sd1443346, -32'sd129018, -32'sd1118559, -32'sd202751, -32'sd205073, -32'sd1612565, -32'sd1167520, -32'sd611474, 32'sd399971, 32'sd611440, -32'sd1323928, -32'sd352736, 32'sd1107517, -32'sd175293, -32'sd2022468, -32'sd891811, -32'sd466978, -32'sd1237806, 32'sd745340, 32'sd1898296, 32'sd746752, 32'sd1041261, -32'sd992175, -32'sd1235371, -32'sd1699891, 32'sd1202687, 32'sd623374, -32'sd294040, -32'sd2624821, -32'sd1112869, -32'sd1167081, 32'sd388379, 32'sd2254359, -32'sd1312909, -32'sd970154, 32'sd1006059, 32'sd1341777, 32'sd729879, -32'sd1502267, 32'sd533917, -32'sd691882, -32'sd787422, 32'sd370138, -32'sd298943, 32'sd1583445, -32'sd656777, 32'sd799829, 32'sd2245118, 32'sd1090293, 32'sd820453, -32'sd1641281, -32'sd1814121, -32'sd1226397, -32'sd823807, 32'sd560511, -32'sd317514, -32'sd471150, -32'sd2498011, -32'sd1609143, 32'sd1371026, 32'sd1890741, -32'sd412055, 32'sd0, -32'sd1012582, 32'sd313464, -32'sd604093, -32'sd255091, -32'sd775463, -32'sd363381, 32'sd861102, -32'sd165695, -32'sd446184, 32'sd578485, 32'sd2143102, 32'sd1618557, 32'sd1222297, -32'sd959976, -32'sd1796175, -32'sd1641020, -32'sd489594, 32'sd402652, 32'sd771918, 32'sd1174011, -32'sd572055, -32'sd127014, 32'sd71589, -32'sd1578183, 32'sd1186628, -32'sd122564, 32'sd0, 32'sd0, 32'sd0, 32'sd1218120, -32'sd286419, -32'sd343924, -32'sd224995, -32'sd1405771, 32'sd274368, 32'sd601124, -32'sd1432246, 32'sd131369, -32'sd313145, 32'sd76679, 32'sd288523, -32'sd863726, -32'sd495007, 32'sd475311, -32'sd332655, -32'sd2430282, 32'sd308128, 32'sd1900063, 32'sd2617582, -32'sd476494, -32'sd915864, -32'sd93108, 32'sd1019155, -32'sd1054044, 32'sd0, 32'sd0, 32'sd0, -32'sd1274731, -32'sd953685, -32'sd979349, -32'sd1323366, -32'sd2058102, -32'sd1622599, 32'sd98108, 32'sd468920, 32'sd1157559, 32'sd248302, 32'sd10339, 32'sd1752421, 32'sd459119, -32'sd185343, -32'sd981135, -32'sd561569, -32'sd3871092, 32'sd311900, 32'sd904096, 32'sd2172761, 32'sd141894, -32'sd311498, 32'sd1551369, -32'sd1580211, -32'sd106552, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd109324, 32'sd22455, -32'sd2758814, -32'sd1648689, -32'sd1935261, 32'sd2116618, -32'sd277698, 32'sd1190680, -32'sd547379, -32'sd2195569, -32'sd2098895, 32'sd66671, -32'sd1970379, -32'sd590697, -32'sd454454, -32'sd253587, -32'sd1980695, -32'sd1257798, -32'sd195008, 32'sd1085111, 32'sd1675460, 32'sd414550, -32'sd511982, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1605212, 32'sd592795, -32'sd165626, -32'sd1278870, -32'sd163465, -32'sd94583, -32'sd2495086, -32'sd947822, -32'sd1401823, -32'sd1559021, -32'sd2269269, -32'sd2203289, -32'sd1292525, -32'sd1421510, -32'sd1055937, -32'sd545825, 32'sd33642, 32'sd1617190, -32'sd491590, 32'sd1436345, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd890743, 32'sd704255, 32'sd1082117, 32'sd888528, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd220040, 32'sd1547862, 32'sd93639, -32'sd1809685, -32'sd28183, -32'sd1703940, -32'sd1703915, 32'sd181320, 32'sd882837, -32'sd829952, 32'sd765054, -32'sd107588, 32'sd2374465, 32'sd1398656, 32'sd1407781, 32'sd39614, 32'sd472876, 32'sd1757251, 32'sd1736605, 32'sd210152, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd355554, 32'sd937681, 32'sd412012, 32'sd509728, 32'sd162209, 32'sd1833440, 32'sd350054, -32'sd2370488, -32'sd2522309, -32'sd2352897, -32'sd150812, -32'sd1484759, 32'sd973215, 32'sd466820, 32'sd1095755, 32'sd2575381, 32'sd516501, 32'sd2109096, 32'sd2000312, -32'sd570182, 32'sd623719, 32'sd110583, -32'sd288887, -32'sd217332, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd60371, 32'sd1332599, 32'sd879571, -32'sd1162966, 32'sd145257, -32'sd176195, -32'sd263207, 32'sd98972, -32'sd1297792, 32'sd322397, 32'sd1937567, 32'sd1958022, 32'sd154371, 32'sd1100019, 32'sd839262, -32'sd742093, -32'sd653268, -32'sd2656776, -32'sd442106, 32'sd203170, -32'sd1164605, 32'sd270250, -32'sd937459, -32'sd998876, 32'sd132695, 32'sd0, 32'sd0, 32'sd282198, 32'sd1003113, 32'sd391341, 32'sd698023, 32'sd267085, -32'sd588235, -32'sd1940188, 32'sd366605, 32'sd1171430, 32'sd1770676, -32'sd1136132, -32'sd1325041, 32'sd779345, 32'sd1864909, -32'sd862205, 32'sd1051237, 32'sd101964, -32'sd1515192, -32'sd843909, -32'sd2544975, -32'sd1915587, -32'sd40298, -32'sd1928342, -32'sd1458253, -32'sd710710, 32'sd609511, 32'sd425203, 32'sd0, 32'sd127922, 32'sd1104400, 32'sd774086, 32'sd692789, 32'sd1281537, 32'sd755789, 32'sd50907, -32'sd799711, 32'sd147612, -32'sd1216423, -32'sd88595, 32'sd370404, -32'sd1380762, 32'sd1123805, 32'sd337494, 32'sd189508, -32'sd749677, -32'sd2766248, 32'sd130027, 32'sd375142, -32'sd730076, -32'sd1201215, -32'sd1671547, -32'sd15677, 32'sd83763, -32'sd1880511, 32'sd916292, 32'sd0, -32'sd210902, 32'sd12935, 32'sd1392384, -32'sd1581542, 32'sd858950, 32'sd1803166, 32'sd964723, 32'sd682058, -32'sd1587253, -32'sd2940625, -32'sd605624, 32'sd360851, -32'sd1071698, 32'sd59981, -32'sd1809631, -32'sd575047, -32'sd2704139, -32'sd1420730, -32'sd485115, -32'sd1130876, -32'sd1237345, -32'sd1707259, 32'sd326783, 32'sd883711, 32'sd1369270, -32'sd1132211, -32'sd980103, -32'sd125079, 32'sd540707, 32'sd10970, 32'sd241251, -32'sd508251, -32'sd5033, -32'sd733264, -32'sd505184, 32'sd557025, -32'sd335919, -32'sd886750, 32'sd1489770, -32'sd268386, -32'sd1899170, -32'sd2563103, -32'sd2268398, -32'sd2907179, -32'sd1158653, -32'sd2868220, -32'sd1266139, -32'sd1083324, 32'sd415198, -32'sd270758, -32'sd2402677, -32'sd383316, 32'sd332050, -32'sd1767464, 32'sd912356, 32'sd631383, 32'sd1196119, -32'sd225017, -32'sd61436, -32'sd704185, 32'sd882709, 32'sd20171, -32'sd26679, 32'sd597390, -32'sd407283, 32'sd1735435, 32'sd784499, -32'sd330620, -32'sd2114586, -32'sd3761056, -32'sd3777859, -32'sd3384873, -32'sd2437201, -32'sd3423883, -32'sd2053992, 32'sd489325, 32'sd210724, -32'sd2233392, -32'sd140639, -32'sd1110748, 32'sd447388, 32'sd372922, -32'sd1091077, -32'sd655805, -32'sd1311162, 32'sd1137788, -32'sd2015194, -32'sd1177335, -32'sd1408026, -32'sd732095, 32'sd1470822, -32'sd809704, 32'sd524246, -32'sd206076, 32'sd1017440, 32'sd268473, -32'sd1661472, -32'sd2023947, -32'sd2092023, 32'sd210548, -32'sd1075060, -32'sd2048101, 32'sd79993, 32'sd983508, 32'sd912009, -32'sd451058, -32'sd1380793, 32'sd614393, -32'sd1757044, 32'sd132841, 32'sd79717, 32'sd180531, 32'sd795305, 32'sd788701, -32'sd2287221, -32'sd1936767, -32'sd99679, 32'sd1118051, -32'sd34469, 32'sd1175005, 32'sd240620, 32'sd339729, 32'sd1315351, 32'sd2204468, -32'sd1406874, -32'sd1191244, 32'sd320707, 32'sd2238653, 32'sd1340871, -32'sd769596, 32'sd1237797, 32'sd158360, 32'sd12924, -32'sd685220, -32'sd309320, 32'sd2165184, -32'sd274053, 32'sd80639, 32'sd420677, -32'sd903757, 32'sd2191752, -32'sd1782145, -32'sd2725813, -32'sd1837155, -32'sd268510, 32'sd877204, -32'sd800370, 32'sd1125490, 32'sd1703441, -32'sd1088804, -32'sd1091418, -32'sd1310200, -32'sd1318826, -32'sd1610323, 32'sd1073817, 32'sd1471319, 32'sd73020, 32'sd1515366, 32'sd449379, 32'sd1455012, 32'sd1601599, -32'sd591749, 32'sd484040, 32'sd658709, 32'sd1098965, -32'sd496256, -32'sd1871391, 32'sd432981, 32'sd696620, -32'sd2543918, -32'sd1186150, 32'sd987571, 32'sd1202157, 32'sd479224, -32'sd669240, 32'sd750617, 32'sd415182, -32'sd289238, 32'sd716416, -32'sd2209968, 32'sd209130, 32'sd623850, -32'sd421738, 32'sd1492912, -32'sd1303383, -32'sd390740, -32'sd1240730, 32'sd2008846, 32'sd859226, 32'sd574842, 32'sd88427, -32'sd250138, 32'sd600291, -32'sd167275, -32'sd1307794, 32'sd5595, -32'sd446598, -32'sd1851516, -32'sd2398408, -32'sd1235692, -32'sd50903, -32'sd1527653, -32'sd2113485, -32'sd1930968, -32'sd1058169, -32'sd1697765, -32'sd2086541, -32'sd649755, 32'sd113288, 32'sd348036, -32'sd529038, 32'sd21090, -32'sd1619482, 32'sd788828, -32'sd140677, 32'sd913839, 32'sd2826786, 32'sd1704125, 32'sd1303403, -32'sd1467790, -32'sd1359423, 32'sd746044, -32'sd370221, -32'sd521489, -32'sd700328, -32'sd949060, 32'sd317117, -32'sd2472445, 32'sd149802, -32'sd198511, -32'sd2234688, -32'sd499816, -32'sd1417495, -32'sd318204, -32'sd301845, 32'sd435645, 32'sd2534596, 32'sd3305666, 32'sd1636225, 32'sd136806, -32'sd1787899, -32'sd1973287, 32'sd863640, 32'sd881865, 32'sd533782, 32'sd789300, -32'sd662377, -32'sd230668, 32'sd1180012, -32'sd268516, -32'sd35513, 32'sd975853, 32'sd964113, -32'sd973056, 32'sd731858, 32'sd314532, 32'sd801444, 32'sd489150, -32'sd184402, -32'sd711713, -32'sd833714, -32'sd2048034, -32'sd2339700, 32'sd367904, 32'sd4481597, 32'sd3238063, 32'sd2249202, 32'sd264418, -32'sd2561871, -32'sd1196266, 32'sd17434, 32'sd479264, 32'sd518294, 32'sd533714, -32'sd33571, 32'sd240331, 32'sd708722, 32'sd699934, 32'sd957119, -32'sd53362, -32'sd564489, -32'sd857114, 32'sd151707, 32'sd352066, 32'sd377937, -32'sd1181613, -32'sd1650448, -32'sd909266, -32'sd1154257, -32'sd1143467, 32'sd1019609, 32'sd1128479, 32'sd582678, 32'sd2860921, 32'sd4151221, 32'sd231823, 32'sd1119033, 32'sd753087, 32'sd909304, 32'sd630888, 32'sd320551, -32'sd215140, 32'sd192611, -32'sd2015324, 32'sd463545, 32'sd490119, -32'sd328668, 32'sd0, 32'sd303120, -32'sd908903, 32'sd932821, 32'sd406796, -32'sd1846926, -32'sd1205869, -32'sd4209843, -32'sd1782619, -32'sd917186, -32'sd434129, 32'sd46977, 32'sd1708185, -32'sd1142743, 32'sd801755, 32'sd3317278, 32'sd1692332, 32'sd1629810, 32'sd2441605, 32'sd947384, 32'sd1043006, -32'sd983131, 32'sd1102233, 32'sd268943, 32'sd1772411, 32'sd956869, -32'sd642310, 32'sd375875, 32'sd1255618, -32'sd52041, 32'sd1393381, 32'sd275699, -32'sd978992, -32'sd2005308, -32'sd2648512, -32'sd338663, 32'sd1573923, 32'sd1266949, 32'sd331339, -32'sd1406576, 32'sd1056351, -32'sd1572380, 32'sd2761910, 32'sd2008719, -32'sd80581, -32'sd409942, 32'sd840975, -32'sd910266, -32'sd1426325, 32'sd1111382, -32'sd154258, 32'sd1283316, 32'sd1716046, 32'sd1918397, -32'sd1579567, 32'sd8464, 32'sd447597, -32'sd486292, 32'sd359321, 32'sd1491791, -32'sd1292794, -32'sd2190807, -32'sd3077114, 32'sd652918, 32'sd1882137, 32'sd1620528, 32'sd2878211, 32'sd1392068, -32'sd1336490, -32'sd545861, -32'sd247674, 32'sd1895059, 32'sd1319383, 32'sd1403194, 32'sd1373106, -32'sd786285, 32'sd913702, 32'sd1289553, -32'sd517030, 32'sd1858592, 32'sd1085875, -32'sd2651, 32'sd339442, 32'sd2045031, 32'sd0, -32'sd1593089, 32'sd1001540, 32'sd462270, -32'sd2049790, -32'sd3620478, -32'sd1407669, -32'sd162108, -32'sd798348, 32'sd790603, 32'sd3182776, 32'sd3100896, 32'sd108584, 32'sd113826, -32'sd674442, 32'sd758317, 32'sd536300, 32'sd36307, 32'sd2892748, 32'sd2073538, 32'sd2569309, -32'sd30143, -32'sd145692, -32'sd411574, 32'sd1844769, -32'sd261956, -32'sd986926, 32'sd471947, -32'sd7876, 32'sd404944, 32'sd274730, 32'sd829383, 32'sd229532, -32'sd1730685, -32'sd1199918, -32'sd987939, 32'sd1828332, 32'sd2296812, 32'sd2012511, -32'sd985000, -32'sd1451173, 32'sd1756154, 32'sd1390103, -32'sd473227, 32'sd782040, 32'sd2620352, 32'sd898926, 32'sd306967, 32'sd742126, -32'sd382148, -32'sd2119333, -32'sd2320724, 32'sd193690, 32'sd780651, -32'sd1887294, 32'sd601708, -32'sd12870, 32'sd183032, -32'sd718562, -32'sd906843, 32'sd593625, 32'sd506522, -32'sd1228337, -32'sd2539229, 32'sd115623, -32'sd1332900, -32'sd291992, -32'sd1356861, -32'sd638772, 32'sd592709, 32'sd325276, -32'sd2292610, -32'sd797243, -32'sd311170, -32'sd1188712, -32'sd1317084, -32'sd1722946, -32'sd723862, -32'sd79652, -32'sd1137605, -32'sd1838689, 32'sd1492441, -32'sd1327277, 32'sd977049, 32'sd0, 32'sd479805, -32'sd1588535, -32'sd795129, -32'sd485063, -32'sd665342, -32'sd1396055, -32'sd2063409, -32'sd962931, -32'sd1046977, -32'sd1226608, -32'sd1855367, 32'sd574793, 32'sd1760301, -32'sd1043253, -32'sd863067, -32'sd2009635, -32'sd1181527, -32'sd3371463, -32'sd3126860, 32'sd701176, 32'sd344515, -32'sd614951, -32'sd1601425, -32'sd736439, 32'sd632180, 32'sd378551, 32'sd0, 32'sd0, 32'sd0, 32'sd152835, -32'sd374415, 32'sd1796097, -32'sd1150517, -32'sd245113, -32'sd2056018, -32'sd954855, 32'sd814802, -32'sd288596, -32'sd1721047, -32'sd2698595, -32'sd2253338, -32'sd425584, -32'sd1450694, -32'sd1172622, -32'sd1530816, -32'sd2141155, -32'sd2482575, -32'sd2022943, 32'sd120139, -32'sd1891460, -32'sd2065810, -32'sd79777, -32'sd311806, -32'sd203577, 32'sd0, 32'sd0, 32'sd0, 32'sd428661, 32'sd741574, -32'sd1078887, -32'sd1354902, -32'sd31297, 32'sd628998, -32'sd73034, -32'sd476486, -32'sd664455, -32'sd691677, -32'sd1445254, -32'sd3707752, -32'sd583836, -32'sd1619468, -32'sd2072487, -32'sd3252788, -32'sd1907408, 32'sd162082, -32'sd405548, -32'sd909262, -32'sd1355735, 32'sd442808, -32'sd955920, 32'sd247027, 32'sd550631, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd116246, -32'sd1171772, 32'sd607896, -32'sd610330, 32'sd1269080, -32'sd1457007, 32'sd656828, -32'sd1518959, 32'sd73259, -32'sd405432, -32'sd1356332, -32'sd3031116, -32'sd1333159, 32'sd1980341, 32'sd1389572, -32'sd1272753, -32'sd795240, -32'sd1290586, -32'sd1292497, -32'sd1024106, -32'sd35373, 32'sd241884, 32'sd36082, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd754115, -32'sd220276, 32'sd686689, 32'sd367422, 32'sd352507, -32'sd757188, 32'sd452315, -32'sd14278, -32'sd396159, 32'sd896419, 32'sd765228, 32'sd1658539, 32'sd922073, 32'sd1032235, 32'sd451053, 32'sd395147, 32'sd77082, -32'sd617788, -32'sd26043, -32'sd435749, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd173212, -32'sd813048, 32'sd551157, -32'sd508475, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1055184, -32'sd101630, -32'sd51790, 32'sd266118, 32'sd141038, 32'sd611772, 32'sd471763, 32'sd260023, 32'sd1169166, -32'sd1407264, -32'sd171634, 32'sd391646, 32'sd1583856, -32'sd418974, 32'sd951835, 32'sd195705, 32'sd372531, -32'sd178017, -32'sd331605, 32'sd578428, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd687709, -32'sd278283, 32'sd979662, 32'sd741347, -32'sd1508572, -32'sd1115869, -32'sd1101758, -32'sd335710, -32'sd1333581, 32'sd811888, 32'sd804774, 32'sd113457, 32'sd1270620, -32'sd1170319, -32'sd736213, 32'sd641578, -32'sd938943, 32'sd661694, 32'sd1425955, 32'sd589941, 32'sd145926, 32'sd1017617, -32'sd272549, 32'sd1023464, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1089302, 32'sd420562, 32'sd7145, -32'sd537979, -32'sd243219, -32'sd529141, -32'sd111259, 32'sd142252, 32'sd1635950, 32'sd969349, 32'sd22677, 32'sd529470, 32'sd98211, 32'sd640743, -32'sd1041180, 32'sd1147177, 32'sd729249, 32'sd773141, -32'sd800185, -32'sd2120517, -32'sd1287881, -32'sd1100195, -32'sd906671, -32'sd343496, 32'sd301169, 32'sd0, 32'sd0, 32'sd790776, -32'sd80749, 32'sd1115127, -32'sd782597, 32'sd639034, -32'sd970743, -32'sd780233, -32'sd1631968, 32'sd590986, 32'sd882353, -32'sd243104, 32'sd958530, -32'sd223167, 32'sd1317023, 32'sd913859, 32'sd527774, -32'sd833574, 32'sd409019, 32'sd427827, -32'sd1644230, 32'sd148774, 32'sd1392380, 32'sd22089, -32'sd1024717, -32'sd2308112, -32'sd1188132, 32'sd210957, 32'sd0, -32'sd180924, -32'sd1180187, -32'sd934331, 32'sd315128, 32'sd980875, -32'sd2082091, -32'sd3190369, -32'sd1210887, -32'sd762933, -32'sd1100620, 32'sd1180147, -32'sd679389, -32'sd2060168, -32'sd2080334, -32'sd996214, -32'sd1772845, -32'sd453219, -32'sd1630322, 32'sd515866, -32'sd1435084, -32'sd733632, 32'sd1045558, -32'sd980830, -32'sd1301421, -32'sd1141199, -32'sd1613998, 32'sd44595, 32'sd0, 32'sd250357, -32'sd1251947, -32'sd1279851, -32'sd535155, 32'sd2312005, 32'sd919241, -32'sd1600303, -32'sd987689, -32'sd2443468, -32'sd577106, 32'sd1958705, 32'sd2324517, -32'sd796334, -32'sd1698320, -32'sd4634285, -32'sd379613, -32'sd1406471, -32'sd1396130, -32'sd510107, 32'sd1345565, 32'sd665607, 32'sd1209549, -32'sd250706, -32'sd1463335, -32'sd296873, -32'sd246743, 32'sd552911, -32'sd137011, 32'sd558831, -32'sd300338, -32'sd1086176, -32'sd168955, 32'sd1044038, 32'sd1754043, -32'sd1445524, -32'sd2859175, 32'sd1637256, 32'sd610794, 32'sd3636915, 32'sd2200916, -32'sd1126431, -32'sd155326, -32'sd3274042, -32'sd3266038, -32'sd875286, -32'sd652049, 32'sd2594661, 32'sd817271, 32'sd112356, 32'sd749621, 32'sd1058698, 32'sd725462, -32'sd1709381, -32'sd157056, -32'sd1050508, -32'sd297007, -32'sd1521630, -32'sd1529824, 32'sd273056, -32'sd1498438, -32'sd364302, 32'sd1370171, 32'sd1896943, -32'sd2508345, 32'sd374669, 32'sd1221356, 32'sd1494001, 32'sd125978, -32'sd1620552, -32'sd2657182, -32'sd2271364, -32'sd2247512, 32'sd1083163, 32'sd794511, 32'sd2778694, 32'sd2750367, 32'sd1099135, -32'sd249562, -32'sd670067, 32'sd976953, 32'sd219867, -32'sd969099, -32'sd138835, 32'sd717541, -32'sd482636, -32'sd1577959, -32'sd451313, -32'sd2231842, -32'sd2051463, -32'sd501542, -32'sd600198, -32'sd1131017, -32'sd661069, 32'sd1617992, 32'sd2077646, 32'sd2190865, -32'sd1256792, -32'sd2667198, -32'sd1509193, 32'sd1097421, 32'sd1572606, 32'sd682929, 32'sd556540, 32'sd924762, 32'sd1825086, -32'sd1091674, -32'sd1789879, -32'sd187128, -32'sd1902304, -32'sd1432822, -32'sd654697, 32'sd683303, 32'sd1059331, 32'sd596707, -32'sd634088, 32'sd375473, -32'sd1026683, -32'sd1651549, -32'sd444171, -32'sd1848928, 32'sd1094806, 32'sd2234477, 32'sd3419129, 32'sd3552826, -32'sd85996, -32'sd1267986, -32'sd1190704, -32'sd2976050, 32'sd493995, 32'sd118611, 32'sd971574, -32'sd1425174, -32'sd95264, -32'sd1285098, -32'sd1759333, -32'sd123414, 32'sd3035113, -32'sd1801222, 32'sd1445864, 32'sd1383183, -32'sd46191, 32'sd325152, -32'sd1464633, -32'sd285266, -32'sd851534, 32'sd665336, -32'sd2904011, -32'sd2496524, -32'sd772549, 32'sd980208, -32'sd61681, 32'sd63990, -32'sd698296, -32'sd1168987, -32'sd279516, -32'sd49196, 32'sd457021, -32'sd262701, -32'sd2187889, -32'sd759450, -32'sd1549050, -32'sd2339159, -32'sd1912079, -32'sd1208969, -32'sd323290, 32'sd599613, 32'sd414203, 32'sd430724, -32'sd121991, -32'sd271450, -32'sd55612, -32'sd3249819, -32'sd1727129, -32'sd1021648, -32'sd926971, -32'sd1132429, -32'sd73052, -32'sd231058, 32'sd1662896, 32'sd374779, 32'sd622709, 32'sd2052983, 32'sd873485, 32'sd308381, 32'sd300689, -32'sd2018733, -32'sd2967251, -32'sd46442, -32'sd738623, -32'sd1845202, -32'sd292406, 32'sd840598, 32'sd649021, 32'sd785679, 32'sd138731, 32'sd230464, -32'sd487831, -32'sd1637090, -32'sd1868600, -32'sd2584911, 32'sd603633, -32'sd1157222, 32'sd585934, 32'sd186737, 32'sd77830, 32'sd109396, 32'sd2274883, 32'sd1403269, 32'sd1005216, 32'sd1748930, 32'sd2306186, 32'sd1131796, 32'sd1527882, -32'sd1241377, -32'sd1718413, 32'sd30671, 32'sd136109, 32'sd1636756, 32'sd930355, 32'sd1279361, -32'sd1855146, -32'sd1596043, 32'sd633670, 32'sd444594, 32'sd78390, -32'sd131675, -32'sd146013, -32'sd603464, 32'sd873424, -32'sd982689, -32'sd1041727, 32'sd254508, -32'sd648151, -32'sd1226425, -32'sd428037, 32'sd1189831, 32'sd240203, 32'sd3207258, 32'sd1939847, -32'sd388283, -32'sd1544430, -32'sd553442, 32'sd80449, -32'sd144309, -32'sd1453495, -32'sd395979, 32'sd660556, -32'sd854777, -32'sd520797, -32'sd709890, -32'sd1363680, 32'sd1400116, -32'sd297946, -32'sd1680368, 32'sd1222598, -32'sd165982, -32'sd785942, -32'sd215424, -32'sd511011, -32'sd1275674, -32'sd1389258, 32'sd1431415, -32'sd248726, 32'sd651291, -32'sd1017248, 32'sd875689, 32'sd1053030, 32'sd746055, 32'sd522897, -32'sd560933, 32'sd808919, 32'sd98467, -32'sd1203974, 32'sd268744, 32'sd598971, -32'sd245563, -32'sd1021746, -32'sd1662343, 32'sd378863, -32'sd457, 32'sd531844, -32'sd2295883, 32'sd147745, 32'sd849810, 32'sd773462, 32'sd741936, 32'sd774022, -32'sd76943, -32'sd715077, -32'sd1437845, -32'sd2002570, 32'sd513246, -32'sd17015, 32'sd945355, 32'sd2955092, 32'sd1731338, -32'sd60514, -32'sd126990, 32'sd527666, -32'sd1161402, 32'sd1738503, -32'sd610565, -32'sd225765, -32'sd3124458, -32'sd1642992, -32'sd1469080, -32'sd137301, 32'sd0, 32'sd581914, -32'sd1108304, -32'sd691758, 32'sd1471510, 32'sd350991, 32'sd1954739, 32'sd349721, 32'sd647772, -32'sd42563, -32'sd1908899, -32'sd2600966, -32'sd2431980, 32'sd1474116, 32'sd1664218, 32'sd2344899, 32'sd1514217, -32'sd931971, -32'sd921888, -32'sd2547991, -32'sd849573, -32'sd153579, -32'sd1402528, -32'sd846664, -32'sd548441, 32'sd73041, 32'sd361796, -32'sd1242312, 32'sd803010, 32'sd1231188, -32'sd284393, 32'sd603039, 32'sd584508, 32'sd686383, -32'sd1636948, -32'sd1100131, -32'sd839858, -32'sd2328988, -32'sd712439, -32'sd2778369, -32'sd2444825, 32'sd1739824, 32'sd1467771, 32'sd436296, 32'sd1789298, -32'sd1979208, -32'sd1000529, 32'sd1516461, 32'sd1873839, -32'sd50821, -32'sd1929576, -32'sd762390, -32'sd1236474, -32'sd1443253, -32'sd428262, 32'sd760581, 32'sd647243, -32'sd1285379, 32'sd750055, 32'sd199688, -32'sd1594636, -32'sd1239446, -32'sd3078420, -32'sd471291, -32'sd864396, -32'sd410148, -32'sd3150336, -32'sd3299927, -32'sd3398903, -32'sd384259, 32'sd1668240, 32'sd1088161, 32'sd1207738, -32'sd129334, -32'sd1145995, -32'sd101217, 32'sd899075, -32'sd2143575, -32'sd1521423, -32'sd2977981, -32'sd77381, 32'sd1407165, -32'sd1149773, 32'sd758567, 32'sd0, -32'sd17632, 32'sd455782, 32'sd251582, -32'sd953470, -32'sd1015331, -32'sd1916532, -32'sd2583433, -32'sd616452, -32'sd1515436, -32'sd1728759, -32'sd1624192, -32'sd241398, -32'sd2133399, 32'sd622345, 32'sd1441543, 32'sd844341, -32'sd575387, 32'sd747832, 32'sd758898, -32'sd1048975, -32'sd3518112, -32'sd433590, -32'sd1404006, -32'sd1161483, 32'sd952189, -32'sd758031, 32'sd739403, 32'sd656031, 32'sd818018, 32'sd1584890, -32'sd589924, 32'sd33858, 32'sd1050252, -32'sd1578965, 32'sd353549, 32'sd187487, -32'sd2671, 32'sd161076, -32'sd1023200, 32'sd114306, -32'sd1524165, 32'sd947152, 32'sd2442902, -32'sd72793, 32'sd262282, 32'sd1200389, 32'sd1194070, -32'sd982451, -32'sd1297501, -32'sd762432, -32'sd278175, 32'sd1312748, 32'sd122413, -32'sd143924, -32'sd263065, 32'sd536912, 32'sd1828582, -32'sd204791, -32'sd297363, 32'sd1667693, 32'sd1891286, 32'sd797342, -32'sd418369, 32'sd168533, -32'sd758477, -32'sd301204, 32'sd1547874, 32'sd306040, -32'sd557184, -32'sd1548246, 32'sd797920, 32'sd1163290, -32'sd648576, 32'sd2019375, -32'sd1136633, -32'sd501350, -32'sd573648, -32'sd2015850, 32'sd511085, 32'sd1790351, -32'sd1136995, 32'sd233249, 32'sd336602, 32'sd0, 32'sd655694, 32'sd889289, -32'sd419573, 32'sd987456, 32'sd1901656, 32'sd1193224, 32'sd1220548, 32'sd252327, 32'sd1590427, 32'sd706497, -32'sd154451, -32'sd26821, 32'sd712737, -32'sd1686977, 32'sd412653, 32'sd1779331, 32'sd145454, 32'sd131945, 32'sd369157, -32'sd833945, 32'sd1575318, 32'sd404261, 32'sd73348, -32'sd257310, -32'sd564364, -32'sd653449, 32'sd0, 32'sd0, 32'sd0, 32'sd354109, -32'sd1518157, -32'sd1036632, 32'sd418627, -32'sd1391977, -32'sd269646, -32'sd8156, 32'sd2014782, -32'sd606104, -32'sd749858, 32'sd419129, -32'sd1185399, -32'sd3255089, -32'sd2255816, -32'sd492886, -32'sd1172971, 32'sd1236796, -32'sd208926, 32'sd1222369, -32'sd235876, 32'sd405307, -32'sd276062, -32'sd59643, 32'sd369418, 32'sd49734, 32'sd0, 32'sd0, 32'sd0, -32'sd357972, -32'sd397358, -32'sd631398, -32'sd198713, 32'sd98201, 32'sd1150941, 32'sd760625, 32'sd998243, -32'sd1133358, -32'sd1496458, 32'sd396686, 32'sd120646, 32'sd1329844, 32'sd687584, -32'sd222883, -32'sd3108152, -32'sd379320, -32'sd1039375, -32'sd332833, -32'sd356493, -32'sd168513, -32'sd350441, 32'sd652415, -32'sd101066, 32'sd385165, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd268797, -32'sd402766, -32'sd1250509, -32'sd1294435, -32'sd13837, 32'sd1447074, -32'sd742990, 32'sd576798, -32'sd406504, -32'sd2107511, -32'sd3535216, -32'sd2100063, -32'sd3029310, 32'sd1171171, 32'sd1387522, -32'sd2231218, -32'sd1130276, 32'sd170750, 32'sd1051016, -32'sd2216930, -32'sd88960, 32'sd527818, -32'sd643968, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd637501, -32'sd49357, 32'sd701384, 32'sd1132938, -32'sd1606401, -32'sd118479, -32'sd681613, -32'sd780384, -32'sd665348, -32'sd681954, -32'sd647004, -32'sd451816, -32'sd481317, -32'sd115485, 32'sd973642, -32'sd66703, 32'sd2016797, -32'sd552947, -32'sd748804, 32'sd457212, 32'sd0, 32'sd0, 32'sd0, 32'sd0}
    };

    localparam logic signed [31:0] layer0_biases [0:127] = '{
        -32'sd2139086, -32'sd61183, -32'sd2716692, 32'sd1491195, -32'sd2025927, 32'sd973610, -32'sd113816, -32'sd1871399, -32'sd2397638, -32'sd1115212, 32'sd21726, -32'sd1225086, -32'sd78274, -32'sd1716191, 32'sd112944, -32'sd101554, 32'sd264733, -32'sd823903, -32'sd744772, 32'sd374569, -32'sd2525431, -32'sd679446, -32'sd601963, -32'sd521449, 32'sd214698, 32'sd143172, -32'sd377562, -32'sd59170, -32'sd2417887, -32'sd737179, -32'sd1493164, 32'sd704328, -32'sd2026122, -32'sd2149869, -32'sd420263, -32'sd1128335, 32'sd1477057, -32'sd1886023, -32'sd458096, -32'sd509175, -32'sd337867, -32'sd1271385, 32'sd110043, 32'sd734814, -32'sd3128944, -32'sd1447739, -32'sd1552562, -32'sd1706958, -32'sd612636, -32'sd680425, -32'sd1356849, -32'sd2690446, -32'sd1732065, -32'sd2634624, -32'sd2090503, -32'sd1423057, 32'sd640393, 32'sd1372582, -32'sd2678528, -32'sd859075, -32'sd1551577, -32'sd1511642, 32'sd775426, -32'sd876349, -32'sd2159295, -32'sd1746623, 32'sd1175956, -32'sd872234, -32'sd868729, -32'sd478563, 32'sd772010, 32'sd1272184, -32'sd740209, -32'sd440004, -32'sd564393, -32'sd117253, -32'sd287076, 32'sd1626306, -32'sd2608846, -32'sd608807, -32'sd1843946, 32'sd2404649, -32'sd3039496, -32'sd791760, -32'sd566307, -32'sd784994, -32'sd1046244, -32'sd183997, -32'sd1976816, -32'sd817898, -32'sd2249845, -32'sd387963, -32'sd4312371, -32'sd67857, -32'sd1846539, -32'sd2529345, -32'sd3750439, -32'sd1761423, -32'sd1856735, -32'sd740413, -32'sd1686855, -32'sd493327, -32'sd1898404, -32'sd53298, -32'sd3958919, -32'sd1078117, 32'sd958036, -32'sd2294904, -32'sd2150007, 32'sd1226028, 32'sd1219076, -32'sd428166, -32'sd754594, 32'sd89263, -32'sd343216, -32'sd1655002, -32'sd765992, -32'sd1122287, -32'sd132881, 32'sd845714, 32'sd1264173, -32'sd1744229, -32'sd4464075, -32'sd1755965, 32'sd1456404, -32'sd87687, -32'sd36186, -32'sd281870
    };

    //Layer 1: 128 inputs, 64 neurons
    localparam logic signed [31:0] layer1_weights [0:63][0:127] = '{
        '{-32'sd2562408, 32'sd4387232, -32'sd1823495, -32'sd3150319, -32'sd1814880, 32'sd852538, 32'sd1545645, -32'sd28787, -32'sd4295431, 32'sd96238, 32'sd972388, -32'sd2523774, 32'sd535334, 32'sd3189803, -32'sd1259025, 32'sd3129232, 32'sd3360, 32'sd508248, 32'sd1695093, 32'sd1138949, -32'sd1803085, 32'sd3041046, -32'sd1247133, -32'sd2697187, 32'sd415668, 32'sd3627218, 32'sd2891178, 32'sd1092796, 32'sd432380, 32'sd2399249, 32'sd4648668, 32'sd2936854, -32'sd1792369, 32'sd159843, -32'sd1114578, 32'sd2343361, -32'sd679969, -32'sd980405, 32'sd679053, -32'sd2642104, 32'sd77654, 32'sd1589644, -32'sd3262600, -32'sd549821, 32'sd866811, -32'sd2068792, -32'sd1823408, -32'sd2663290, 32'sd912021, -32'sd77824, -32'sd1538227, -32'sd1743895, -32'sd325121, -32'sd2843429, 32'sd1295257, -32'sd6019772, -32'sd1335336, 32'sd3300637, 32'sd1904623, 32'sd1362256, -32'sd2975949, 32'sd35051, -32'sd14446, 32'sd620705, 32'sd379851, 32'sd436579, -32'sd1375514, 32'sd2122101, 32'sd336907, 32'sd130123, 32'sd1768457, 32'sd4431225, 32'sd2683938, 32'sd794928, 32'sd3853168, 32'sd552609, -32'sd2302879, 32'sd1848079, -32'sd3728824, 32'sd640510, -32'sd1583278, 32'sd2787903, 32'sd1451212, 32'sd1539332, 32'sd2055969, 32'sd1509716, -32'sd663061, 32'sd2768242, -32'sd236262, 32'sd2147114, 32'sd2433962, 32'sd2494682, -32'sd1204524, -32'sd3061393, 32'sd2971883, -32'sd3425438, 32'sd1901615, -32'sd3743301, 32'sd4363727, 32'sd526495, -32'sd1855342, -32'sd1474664, 32'sd1295784, 32'sd686310, -32'sd83643, 32'sd4429071, -32'sd2883398, 32'sd803125, -32'sd569533, 32'sd2871446, -32'sd160333, -32'sd3528981, 32'sd2105996, 32'sd1277989, -32'sd2056103, -32'sd136128, 32'sd4556952, -32'sd529038, 32'sd4211393, 32'sd580424, 32'sd1111786, -32'sd819812, 32'sd152923, -32'sd1294025, 32'sd3064686, 32'sd2571543, 32'sd2541353, 32'sd2051415},
        '{32'sd1841416, -32'sd2378645, -32'sd2100559, -32'sd1812147, -32'sd2836692, -32'sd2649980, -32'sd1484856, -32'sd3498719, -32'sd3346489, -32'sd1673902, 32'sd2559156, -32'sd2774361, -32'sd776583, 32'sd1094246, 32'sd4682553, -32'sd1536277, 32'sd3502395, -32'sd1366000, 32'sd3437152, 32'sd3359830, -32'sd3219249, 32'sd2419320, 32'sd1149261, -32'sd4447351, 32'sd2962136, 32'sd73283, 32'sd3149597, 32'sd3959134, -32'sd2914227, -32'sd1215219, 32'sd2114788, 32'sd1285567, 32'sd2457643, 32'sd1827177, 32'sd1662604, -32'sd2851184, -32'sd4060611, -32'sd1469614, -32'sd899462, -32'sd679280, -32'sd3489688, -32'sd1742729, 32'sd3312453, 32'sd3678607, -32'sd463374, -32'sd2539297, -32'sd3323916, 32'sd1622853, 32'sd595773, 32'sd1196509, 32'sd2164848, 32'sd5025395, -32'sd528168, -32'sd555163, 32'sd678273, 32'sd377504, -32'sd2769330, -32'sd2240649, 32'sd328358, 32'sd4263496, 32'sd2444833, -32'sd1796867, -32'sd2449190, -32'sd1564336, -32'sd315125, -32'sd406825, -32'sd2644642, 32'sd837975, -32'sd1542680, 32'sd883789, -32'sd3911142, 32'sd64497, 32'sd1828094, 32'sd2302693, -32'sd676526, 32'sd3542308, 32'sd987427, 32'sd712929, 32'sd2928341, -32'sd169558, 32'sd2938223, -32'sd324462, 32'sd213699, -32'sd562824, -32'sd1780365, 32'sd1431725, -32'sd2035281, -32'sd1420782, 32'sd719882, 32'sd757940, 32'sd3122677, 32'sd4182406, 32'sd1945767, 32'sd1948330, -32'sd1933857, 32'sd1017101, -32'sd900720, 32'sd854054, 32'sd2725618, 32'sd1574022, -32'sd633784, 32'sd1559794, -32'sd2312507, 32'sd1282658, -32'sd1757337, 32'sd352443, -32'sd2968460, -32'sd1958009, -32'sd181799, -32'sd73435, -32'sd3248070, -32'sd2745720, 32'sd1118780, 32'sd429919, 32'sd2420389, -32'sd2602154, 32'sd1771245, -32'sd1445179, 32'sd2959292, -32'sd33762, 32'sd80352, 32'sd1421122, 32'sd2375060, -32'sd1613222, 32'sd737644, 32'sd1388982, -32'sd772742, -32'sd4346137},
        '{32'sd1741946, 32'sd1414829, -32'sd631836, -32'sd2284326, -32'sd4775333, 32'sd2800278, 32'sd1615350, -32'sd228826, 32'sd3154497, 32'sd794256, 32'sd367747, -32'sd1922306, 32'sd3674996, 32'sd1068899, -32'sd1051898, -32'sd1597263, 32'sd1586303, -32'sd414651, 32'sd480470, -32'sd116879, -32'sd637367, -32'sd3891274, 32'sd3178972, -32'sd3296533, 32'sd3631792, -32'sd3674428, -32'sd222570, -32'sd408973, -32'sd3131354, 32'sd1051112, -32'sd2579967, -32'sd2943492, 32'sd884199, -32'sd1008096, 32'sd909899, 32'sd2178167, 32'sd170617, 32'sd1241287, -32'sd2432186, 32'sd2555498, 32'sd2381480, -32'sd1637422, -32'sd495739, 32'sd2223506, -32'sd797832, -32'sd682413, -32'sd1207686, 32'sd1470966, 32'sd4770781, 32'sd4058302, 32'sd2417530, 32'sd6233357, 32'sd1482394, -32'sd2345827, -32'sd4457997, -32'sd3919344, 32'sd577086, 32'sd997322, 32'sd920809, -32'sd916802, -32'sd3350901, 32'sd2055264, -32'sd1243826, 32'sd966941, 32'sd1178701, 32'sd1687947, 32'sd183857, -32'sd851784, 32'sd2130327, -32'sd1199263, 32'sd3097463, 32'sd405611, -32'sd4015709, 32'sd2858768, 32'sd1960101, -32'sd1689237, 32'sd2480993, -32'sd849853, -32'sd5050041, -32'sd1587470, 32'sd1595941, 32'sd3902327, 32'sd4790179, 32'sd2718225, -32'sd2261231, 32'sd2987661, -32'sd90370, 32'sd309549, 32'sd288531, -32'sd487861, 32'sd1791586, -32'sd1990790, -32'sd2444978, -32'sd4265552, 32'sd1870085, -32'sd986957, 32'sd1310851, 32'sd2920202, 32'sd4214355, 32'sd1439086, 32'sd798877, -32'sd772384, -32'sd841201, -32'sd4182827, 32'sd721618, 32'sd1232675, -32'sd26502, -32'sd867333, -32'sd1839002, -32'sd1770774, 32'sd2111682, -32'sd437725, -32'sd2068482, 32'sd3317949, 32'sd121528, -32'sd606018, -32'sd1364440, 32'sd868419, 32'sd3219777, 32'sd1338866, 32'sd327614, -32'sd1647187, -32'sd3374938, 32'sd1630895, -32'sd572532, 32'sd3085295, -32'sd3046468, -32'sd2694881},
        '{32'sd827222, -32'sd273151, 32'sd3710924, -32'sd307377, -32'sd2121460, -32'sd1008515, 32'sd2081724, -32'sd845105, -32'sd2573217, 32'sd2501291, 32'sd2052453, 32'sd3994654, 32'sd3233359, -32'sd3619321, -32'sd584296, -32'sd165745, -32'sd6476206, 32'sd287770, 32'sd1195080, -32'sd1466035, -32'sd4296173, -32'sd1502575, -32'sd296937, 32'sd85263, 32'sd2231564, 32'sd4628432, -32'sd171198, 32'sd1912573, 32'sd1867380, -32'sd1346839, -32'sd1081419, 32'sd2525840, 32'sd2092335, -32'sd1804713, -32'sd1347351, 32'sd647870, 32'sd235665, 32'sd3125924, -32'sd808084, 32'sd1403415, 32'sd3858768, 32'sd3158886, -32'sd4224730, -32'sd542091, -32'sd3146739, 32'sd592082, -32'sd813232, 32'sd2491756, 32'sd543839, 32'sd1697326, 32'sd1322132, 32'sd2327633, 32'sd3617340, -32'sd1473012, -32'sd2755603, 32'sd1860519, -32'sd415386, 32'sd1515216, -32'sd1595105, 32'sd672697, -32'sd186414, -32'sd3411980, -32'sd4323048, -32'sd2907428, 32'sd2270980, 32'sd4964603, 32'sd62335, 32'sd331856, 32'sd1386298, 32'sd230701, -32'sd2688979, 32'sd91447, -32'sd2879063, -32'sd1151889, 32'sd723889, 32'sd3752057, -32'sd296541, -32'sd3074962, -32'sd1422429, -32'sd1641642, -32'sd4077, 32'sd2097352, -32'sd187037, -32'sd2413250, 32'sd2216935, 32'sd2079508, -32'sd59225, -32'sd584566, -32'sd1008507, 32'sd2596993, 32'sd260881, -32'sd2622871, 32'sd2875892, 32'sd2230775, -32'sd2672951, 32'sd5626295, 32'sd4717618, -32'sd235800, -32'sd1173454, 32'sd1660046, -32'sd1733458, -32'sd1415946, 32'sd1296164, -32'sd2306097, -32'sd1206509, -32'sd127120, -32'sd2468626, -32'sd1352552, 32'sd173655, -32'sd1147032, -32'sd2848048, 32'sd973794, -32'sd3944826, 32'sd1264159, 32'sd2835860, -32'sd2653206, -32'sd2579403, -32'sd1518312, 32'sd3312258, -32'sd254000, 32'sd3641929, 32'sd1452293, -32'sd957052, 32'sd818491, -32'sd4028191, 32'sd28493, 32'sd1835140, -32'sd1368662},
        '{32'sd1886386, -32'sd1504175, 32'sd3382593, 32'sd2984420, 32'sd1709446, -32'sd1927329, 32'sd1439519, -32'sd1616865, -32'sd264791, 32'sd1735012, 32'sd2084527, -32'sd2047493, 32'sd3246196, 32'sd2074229, -32'sd2740479, -32'sd1986854, -32'sd2255215, 32'sd2453945, 32'sd2330258, 32'sd3928021, 32'sd982739, 32'sd564122, 32'sd2501552, 32'sd3276639, 32'sd401719, -32'sd2241433, 32'sd2338269, 32'sd4002611, -32'sd2595800, -32'sd2799135, -32'sd2434612, 32'sd3936249, -32'sd2250888, -32'sd2062925, -32'sd2431143, -32'sd675198, 32'sd515285, -32'sd114210, 32'sd1402869, -32'sd2339385, -32'sd910914, -32'sd3447601, -32'sd682302, 32'sd898664, -32'sd3075203, -32'sd4772584, -32'sd1809439, -32'sd1449869, 32'sd1248228, 32'sd3884622, -32'sd4986515, 32'sd2070276, -32'sd469663, -32'sd630433, 32'sd2684525, 32'sd654820, -32'sd1156688, -32'sd1955508, 32'sd2900981, -32'sd1962512, -32'sd4236385, -32'sd1915924, -32'sd904699, 32'sd2171244, 32'sd502088, -32'sd717450, -32'sd5518227, 32'sd1862572, 32'sd1650246, -32'sd2880183, 32'sd1928703, 32'sd2725954, -32'sd2825428, -32'sd2344361, -32'sd1544859, -32'sd1710063, -32'sd1192648, 32'sd4338662, -32'sd2323429, -32'sd2512047, 32'sd1316048, 32'sd1560049, -32'sd3525601, -32'sd2964706, -32'sd4948880, 32'sd3235536, 32'sd2429630, -32'sd1898525, -32'sd2247299, 32'sd3537541, 32'sd3769175, -32'sd2982157, -32'sd73843, 32'sd2350957, -32'sd1346244, -32'sd2091808, -32'sd1611416, 32'sd1981161, 32'sd2806722, 32'sd1197359, -32'sd1956907, 32'sd265932, 32'sd4622376, -32'sd2923343, -32'sd1367440, -32'sd1421778, -32'sd1284886, 32'sd1642490, 32'sd3077167, 32'sd585956, -32'sd3549065, 32'sd274578, 32'sd3883178, -32'sd2078950, -32'sd1594846, 32'sd1916997, -32'sd2190875, -32'sd771279, -32'sd60930, -32'sd1018887, 32'sd47679, -32'sd1917740, 32'sd2791, 32'sd858286, 32'sd3269992, -32'sd378963, 32'sd861597, 32'sd500120},
        '{32'sd2865290, 32'sd158667, 32'sd1171791, 32'sd3654500, -32'sd3140909, -32'sd3951672, -32'sd398929, -32'sd685207, -32'sd3192648, 32'sd2109950, -32'sd3644579, -32'sd2513087, -32'sd2684014, 32'sd1007353, -32'sd1080473, -32'sd1301686, -32'sd3155222, 32'sd735853, -32'sd2535486, 32'sd44325, 32'sd305886, -32'sd1842422, 32'sd1508562, 32'sd2250807, -32'sd3198917, -32'sd3273947, 32'sd183152, -32'sd3405588, -32'sd756921, 32'sd2511358, 32'sd640365, -32'sd604980, -32'sd915867, -32'sd3139401, 32'sd860578, 32'sd356879, -32'sd1518261, -32'sd2740043, 32'sd1230064, 32'sd3010816, -32'sd2222926, 32'sd2890896, 32'sd929230, 32'sd1750565, -32'sd688105, -32'sd2109653, -32'sd1937182, 32'sd2647659, 32'sd2796708, 32'sd3424058, 32'sd2740392, 32'sd1784491, 32'sd358175, -32'sd616871, 32'sd96819, 32'sd1642729, 32'sd1199622, -32'sd387679, -32'sd4312057, -32'sd2619176, -32'sd1462130, -32'sd2356018, 32'sd1344481, 32'sd1898852, -32'sd471263, 32'sd5292145, -32'sd4508250, -32'sd1203951, -32'sd3044193, 32'sd4202075, -32'sd2127840, -32'sd4955690, -32'sd1111678, 32'sd103129, 32'sd704929, 32'sd4416004, 32'sd3102671, 32'sd1638174, 32'sd3237315, -32'sd3452225, -32'sd646177, 32'sd3151909, -32'sd579427, -32'sd1167961, 32'sd2436966, 32'sd1057735, 32'sd628886, -32'sd3531531, 32'sd353092, 32'sd5018432, -32'sd197703, 32'sd3152848, 32'sd104944, -32'sd806456, 32'sd2669984, 32'sd2213740, -32'sd625152, 32'sd537198, -32'sd6425261, -32'sd3668882, -32'sd696026, 32'sd3764601, 32'sd849412, 32'sd3223301, 32'sd270122, -32'sd2788221, 32'sd3436641, 32'sd1214129, -32'sd4005439, -32'sd3941935, -32'sd2675291, 32'sd1726493, 32'sd692324, 32'sd2067982, -32'sd181418, -32'sd1545191, 32'sd461781, 32'sd3162966, 32'sd3144788, -32'sd578237, 32'sd1012219, 32'sd1149945, 32'sd3309229, -32'sd12041, -32'sd4085460, -32'sd1291545, 32'sd1896354, -32'sd3025892},
        '{32'sd3473665, 32'sd3923165, 32'sd925130, -32'sd2594916, -32'sd1478843, 32'sd3871690, 32'sd3144866, 32'sd1027734, 32'sd2375409, -32'sd798969, 32'sd1419894, 32'sd918184, 32'sd3207657, 32'sd1935753, -32'sd2102616, 32'sd3474928, -32'sd3750, -32'sd4074035, -32'sd1197616, -32'sd2262080, -32'sd3006256, 32'sd4023552, -32'sd1630243, -32'sd3716403, -32'sd1792336, -32'sd907826, -32'sd966193, -32'sd2260551, -32'sd286444, 32'sd1670511, 32'sd2477997, 32'sd3131488, -32'sd958641, 32'sd411226, 32'sd1044091, 32'sd2609493, -32'sd774139, 32'sd2507612, 32'sd2570272, 32'sd607544, -32'sd315583, 32'sd500872, 32'sd2977135, 32'sd1892441, 32'sd1955390, -32'sd161552, -32'sd2441276, 32'sd2212107, 32'sd886706, 32'sd2526122, -32'sd2063196, 32'sd1362805, -32'sd1256165, 32'sd3121543, -32'sd809298, 32'sd2449200, 32'sd2355296, 32'sd2266667, 32'sd2058545, 32'sd198669, 32'sd408014, 32'sd3057931, -32'sd2017163, 32'sd2603915, -32'sd2095110, 32'sd3706823, 32'sd5027722, -32'sd2171573, 32'sd1097123, -32'sd859245, -32'sd1321057, -32'sd4538328, -32'sd502374, -32'sd1571142, -32'sd1299417, 32'sd2827438, -32'sd272802, -32'sd2105353, 32'sd1425566, 32'sd417269, -32'sd3386635, 32'sd2749030, -32'sd1633011, 32'sd1257245, -32'sd2930979, 32'sd1478812, -32'sd5758951, -32'sd2759662, -32'sd2221134, 32'sd430422, -32'sd3535994, -32'sd2602499, 32'sd3025689, 32'sd2609096, -32'sd778668, 32'sd3529351, -32'sd351555, -32'sd123956, -32'sd1184739, 32'sd3898525, -32'sd1126180, -32'sd5363461, 32'sd49502, 32'sd393376, 32'sd1000970, 32'sd3282911, -32'sd2180362, -32'sd1428127, -32'sd2243346, 32'sd2702693, -32'sd34108, -32'sd1602596, -32'sd2769154, -32'sd227296, 32'sd1521277, -32'sd3153716, -32'sd2627263, -32'sd3225466, -32'sd52750, -32'sd637744, 32'sd3241719, 32'sd1860599, 32'sd283442, -32'sd936494, -32'sd103713, -32'sd1588651, 32'sd1539558, -32'sd2340735},
        '{32'sd4603869, 32'sd3171218, -32'sd696773, -32'sd2513756, -32'sd3151846, 32'sd795629, 32'sd4622300, -32'sd1813182, 32'sd2527299, -32'sd1223331, 32'sd3191718, 32'sd349588, -32'sd1041695, 32'sd1528156, 32'sd442369, 32'sd3839140, -32'sd1433152, -32'sd42801, 32'sd3340470, 32'sd4535968, 32'sd3775698, -32'sd2055434, 32'sd3323265, 32'sd1093789, -32'sd27949, -32'sd1771932, 32'sd1243120, -32'sd1132630, -32'sd1518110, -32'sd2880076, -32'sd1857830, 32'sd1166751, -32'sd1135512, -32'sd383899, 32'sd2232988, -32'sd1440701, -32'sd199891, 32'sd2210049, 32'sd1535440, 32'sd5215644, -32'sd2408608, -32'sd441749, 32'sd3240781, 32'sd3695109, -32'sd3119092, 32'sd2679984, 32'sd1482749, 32'sd2550482, -32'sd2495007, 32'sd4806908, -32'sd4528796, -32'sd1074172, 32'sd472305, 32'sd3075696, 32'sd1713578, 32'sd2391999, -32'sd2228605, -32'sd1906227, -32'sd580075, 32'sd1423619, -32'sd335620, 32'sd627345, -32'sd1343400, 32'sd821939, 32'sd2928639, 32'sd2137760, -32'sd84819, 32'sd1070251, -32'sd2393258, 32'sd197560, -32'sd1162552, -32'sd1242796, 32'sd2082120, -32'sd4219336, 32'sd1081044, -32'sd287940, 32'sd3496585, -32'sd864058, -32'sd1980937, 32'sd734637, 32'sd215406, 32'sd3609829, -32'sd2564875, -32'sd701611, -32'sd4198537, -32'sd2048854, 32'sd562718, -32'sd2833312, 32'sd50796, -32'sd2207652, 32'sd3820040, -32'sd2819495, 32'sd3108120, -32'sd1797064, 32'sd4842376, -32'sd3531798, -32'sd1594946, -32'sd1037891, 32'sd1930511, 32'sd1829640, 32'sd3993661, 32'sd1152259, -32'sd1127233, -32'sd908156, 32'sd2241269, -32'sd361612, -32'sd519107, 32'sd701947, -32'sd4937885, 32'sd4484250, -32'sd1264905, -32'sd1688125, -32'sd2691238, -32'sd1603433, 32'sd1754893, 32'sd3469582, -32'sd1280122, 32'sd1859946, -32'sd1203270, 32'sd1717266, -32'sd3650763, -32'sd1733675, -32'sd5798407, 32'sd2701675, 32'sd2971291, -32'sd2106313, -32'sd2361520, 32'sd94526},
        '{32'sd751570, -32'sd3047704, -32'sd1818626, 32'sd510654, -32'sd3224040, -32'sd3092031, -32'sd442029, -32'sd2392566, 32'sd659250, 32'sd2512054, 32'sd690414, -32'sd2720399, 32'sd2475912, -32'sd256764, -32'sd2982681, -32'sd2514836, -32'sd46477, -32'sd715888, 32'sd1294425, -32'sd1348945, -32'sd3012472, -32'sd1420093, -32'sd2632918, 32'sd315962, -32'sd1122821, 32'sd2117425, -32'sd2633601, -32'sd1854138, -32'sd650322, -32'sd3446950, -32'sd4401137, -32'sd1949991, -32'sd2968311, 32'sd1509624, 32'sd1488257, 32'sd2405243, 32'sd312194, 32'sd1257587, 32'sd1403547, 32'sd1511903, 32'sd1105232, 32'sd1397562, -32'sd4725691, -32'sd1786955, -32'sd2625002, 32'sd689270, 32'sd633786, -32'sd1633661, -32'sd1169849, -32'sd211180, -32'sd1187683, -32'sd3401714, 32'sd2721087, 32'sd1086598, -32'sd2385791, 32'sd2241271, -32'sd2154428, 32'sd2178795, -32'sd1812425, 32'sd2981529, 32'sd315630, 32'sd2388476, 32'sd3116516, 32'sd2073555, -32'sd3803722, -32'sd2202352, 32'sd2783729, 32'sd4243788, -32'sd2520838, -32'sd3306366, 32'sd2580367, -32'sd2327137, -32'sd3105766, -32'sd4390168, -32'sd2543295, 32'sd2015439, 32'sd1068956, 32'sd2043144, -32'sd2562551, 32'sd990574, -32'sd1463104, 32'sd706400, 32'sd635063, 32'sd2236541, 32'sd663223, 32'sd670165, 32'sd896555, 32'sd2948771, 32'sd1121142, -32'sd5448164, -32'sd3035067, 32'sd1453812, -32'sd834272, -32'sd3087277, -32'sd2388927, 32'sd74927, 32'sd2649824, -32'sd2903510, -32'sd527598, -32'sd62020, -32'sd3165218, 32'sd4448573, 32'sd1153992, 32'sd3922050, -32'sd514825, 32'sd3647089, 32'sd379365, 32'sd2111038, -32'sd1181319, 32'sd3431334, 32'sd830497, 32'sd1351783, -32'sd656148, 32'sd4348954, -32'sd891714, -32'sd2457472, 32'sd3958428, -32'sd2726465, 32'sd4317899, -32'sd131774, 32'sd2623866, -32'sd2139653, -32'sd2427864, 32'sd3358565, -32'sd764574, 32'sd1442528, 32'sd1819942, 32'sd1136816},
        '{-32'sd609751, -32'sd278410, -32'sd1740991, 32'sd3923207, 32'sd1258990, -32'sd839176, 32'sd998995, -32'sd2984769, 32'sd790648, -32'sd1844265, -32'sd2833020, -32'sd1593241, 32'sd2687781, 32'sd3871948, 32'sd4424942, 32'sd2235972, 32'sd1797161, 32'sd2106491, 32'sd2787864, 32'sd2893215, -32'sd1939813, 32'sd2399395, -32'sd2360230, 32'sd1608821, -32'sd4950356, -32'sd2697230, 32'sd3799688, -32'sd2514798, -32'sd1335704, -32'sd1978465, 32'sd654673, 32'sd97877, -32'sd419231, 32'sd3227380, 32'sd3920134, 32'sd2274791, 32'sd2736791, -32'sd2119932, 32'sd1601095, -32'sd1931688, 32'sd1061769, 32'sd3577135, 32'sd1915274, -32'sd4736166, 32'sd243737, -32'sd3004943, -32'sd1893769, -32'sd1883141, -32'sd3488143, -32'sd1156743, -32'sd707655, -32'sd45920, -32'sd2661167, 32'sd1063828, -32'sd1472838, -32'sd1095315, -32'sd1275494, -32'sd1374536, 32'sd979626, 32'sd3068068, 32'sd2194527, 32'sd682731, 32'sd2566181, -32'sd689511, 32'sd249992, -32'sd2917958, 32'sd853275, 32'sd4435620, -32'sd591116, 32'sd316360, -32'sd2175896, 32'sd852181, -32'sd1947242, 32'sd1677849, -32'sd731264, -32'sd1152697, -32'sd3158898, -32'sd1349508, -32'sd969722, 32'sd2468720, 32'sd1873672, -32'sd2245048, -32'sd1196456, 32'sd2984457, -32'sd1098663, 32'sd3779230, -32'sd1736650, -32'sd3776796, 32'sd668097, 32'sd2187527, 32'sd486378, 32'sd1798043, 32'sd1339587, 32'sd3709232, -32'sd1537736, -32'sd3350514, -32'sd3610519, 32'sd507469, -32'sd1604430, -32'sd3795064, -32'sd4827385, 32'sd3202071, -32'sd2433796, 32'sd2135159, -32'sd1325928, -32'sd541019, -32'sd2023352, 32'sd3255748, 32'sd1859163, 32'sd2812221, 32'sd1154376, 32'sd1852947, -32'sd925621, -32'sd934981, 32'sd2168035, -32'sd685227, 32'sd1750814, 32'sd162401, 32'sd3082102, 32'sd699411, 32'sd1019021, -32'sd1540919, 32'sd2528348, -32'sd67493, -32'sd724073, -32'sd4284674, 32'sd3060079, 32'sd26923},
        '{32'sd1487412, -32'sd3591943, -32'sd1641854, 32'sd735461, 32'sd2542027, 32'sd647669, -32'sd2745972, -32'sd3732837, 32'sd4360199, -32'sd2137922, 32'sd3816022, 32'sd3675676, 32'sd847903, 32'sd3363106, 32'sd1453059, -32'sd3282124, -32'sd3020346, 32'sd1606252, -32'sd1759117, -32'sd2788298, -32'sd1988078, 32'sd1450857, -32'sd2962209, 32'sd2036249, -32'sd2191135, 32'sd1027148, -32'sd4582145, -32'sd2196833, -32'sd1246163, -32'sd1327991, -32'sd4419714, 32'sd1472493, 32'sd1400691, -32'sd2821756, -32'sd995936, -32'sd1211306, -32'sd3590027, 32'sd2792177, -32'sd2417067, 32'sd2077287, -32'sd1492439, 32'sd134172, -32'sd785688, -32'sd645163, -32'sd1285739, -32'sd2952571, -32'sd689499, -32'sd3421130, -32'sd730072, -32'sd3377476, 32'sd3229183, 32'sd592859, -32'sd4274304, 32'sd2162523, -32'sd767668, 32'sd3303297, 32'sd2048818, 32'sd1490900, 32'sd3285588, 32'sd2724032, 32'sd364962, -32'sd2290385, -32'sd1451898, 32'sd1604686, 32'sd1880250, 32'sd1162088, 32'sd3232434, 32'sd2251891, -32'sd3914618, -32'sd2495861, 32'sd2990755, -32'sd822241, 32'sd3610300, 32'sd690127, 32'sd2886909, -32'sd1105706, -32'sd3442935, 32'sd2526076, 32'sd2638688, 32'sd3462857, -32'sd2716861, -32'sd1361781, -32'sd651662, 32'sd1517983, 32'sd1042523, -32'sd2743587, 32'sd60698, 32'sd588027, 32'sd1669699, 32'sd2975780, 32'sd843689, -32'sd1281685, 32'sd1156931, 32'sd4325262, -32'sd2461577, 32'sd3840089, -32'sd961970, 32'sd1128775, 32'sd3462971, -32'sd2845262, 32'sd2610956, -32'sd999277, -32'sd3199904, -32'sd3105424, -32'sd3570313, 32'sd1996792, 32'sd90543, -32'sd4321398, -32'sd1545345, 32'sd1588966, -32'sd4899724, -32'sd2690653, -32'sd1815506, 32'sd991670, 32'sd3861630, 32'sd4137179, 32'sd2861886, 32'sd4143645, -32'sd2022505, -32'sd64471, 32'sd3878726, 32'sd1098741, -32'sd548476, -32'sd266268, -32'sd2729792, 32'sd1811657, -32'sd4326937, 32'sd2605143},
        '{32'sd2976702, 32'sd3547503, -32'sd2169872, 32'sd1374071, 32'sd1233636, 32'sd2573580, -32'sd1595232, -32'sd3130522, 32'sd1500108, -32'sd1987081, -32'sd340591, -32'sd506506, -32'sd3012695, -32'sd212796, 32'sd2401503, 32'sd2309377, -32'sd1786541, 32'sd1678627, 32'sd1089688, 32'sd561978, -32'sd1170479, 32'sd1555352, 32'sd3348105, 32'sd1283653, 32'sd36217, 32'sd2526822, 32'sd1625862, -32'sd2610766, -32'sd291141, -32'sd1836839, 32'sd2572815, -32'sd429758, -32'sd3622561, 32'sd143318, -32'sd1261012, 32'sd3191718, -32'sd2618904, -32'sd828076, 32'sd1544716, 32'sd5369496, -32'sd1737725, -32'sd69152, -32'sd1133684, -32'sd1123685, 32'sd5016955, -32'sd51876, 32'sd883719, 32'sd2722473, -32'sd2788975, 32'sd207312, -32'sd4217924, 32'sd219215, 32'sd3069446, 32'sd2114499, -32'sd915149, -32'sd3296187, -32'sd2383170, 32'sd217094, 32'sd480818, 32'sd1147738, -32'sd3220166, -32'sd8198, 32'sd1633803, -32'sd249, 32'sd753771, -32'sd2594459, 32'sd2715474, -32'sd4287331, 32'sd2205572, -32'sd1627866, 32'sd3040011, -32'sd169533, -32'sd948396, -32'sd1131528, 32'sd282476, 32'sd100859, 32'sd1275046, -32'sd1608730, -32'sd1314699, 32'sd1978327, -32'sd2485215, -32'sd1863645, 32'sd5320253, -32'sd737915, -32'sd3356885, 32'sd1495749, 32'sd2655346, -32'sd1623997, 32'sd1428128, 32'sd2597417, -32'sd3624055, -32'sd3863848, 32'sd1096255, 32'sd3303203, -32'sd2268625, -32'sd1888441, 32'sd550914, 32'sd123187, -32'sd1663617, 32'sd1485802, 32'sd3150876, 32'sd1099098, 32'sd2404563, -32'sd3520605, 32'sd2628435, 32'sd1599118, -32'sd3633201, 32'sd195095, -32'sd4022528, 32'sd3938524, -32'sd977838, -32'sd288463, -32'sd1450349, 32'sd4148328, 32'sd2668366, -32'sd2987954, -32'sd348521, -32'sd1842169, 32'sd2363785, 32'sd3114097, -32'sd3310889, 32'sd1726641, -32'sd2633769, -32'sd3174985, 32'sd3282545, -32'sd2872315, 32'sd987956, 32'sd159375},
        '{32'sd2866862, 32'sd2251836, -32'sd2624290, -32'sd297667, -32'sd3796498, 32'sd3635489, 32'sd936564, 32'sd3468543, 32'sd1785975, -32'sd2439108, 32'sd346491, 32'sd959696, 32'sd2785677, -32'sd414972, -32'sd333804, 32'sd2325546, 32'sd592348, -32'sd2581175, -32'sd2363366, -32'sd3815653, -32'sd453335, -32'sd751301, -32'sd1968784, 32'sd1387046, -32'sd4438325, -32'sd847708, 32'sd703476, -32'sd2809252, -32'sd221340, 32'sd3642901, -32'sd3428350, 32'sd1188613, 32'sd1222365, 32'sd998781, -32'sd762148, 32'sd1191782, 32'sd3667478, 32'sd2821197, 32'sd425963, -32'sd2893929, -32'sd2031733, 32'sd1215128, 32'sd2804121, -32'sd2326765, 32'sd1894958, 32'sd2070604, 32'sd3849123, -32'sd3142135, 32'sd724364, 32'sd3020758, 32'sd3288137, -32'sd4577184, -32'sd2113781, -32'sd3531631, -32'sd1508492, -32'sd316185, 32'sd2375359, -32'sd547697, -32'sd4615560, 32'sd1316175, 32'sd160611, 32'sd3369572, -32'sd177127, 32'sd4511298, 32'sd731088, -32'sd869165, -32'sd2229044, 32'sd2303883, 32'sd1208744, -32'sd2914577, -32'sd147971, 32'sd2520767, 32'sd1487609, 32'sd1411682, 32'sd3533718, -32'sd2911399, 32'sd647762, 32'sd2038842, 32'sd2246945, -32'sd649662, 32'sd1408566, -32'sd906464, -32'sd1666421, -32'sd3241492, -32'sd886243, 32'sd1310769, -32'sd2476814, -32'sd3456520, 32'sd4189563, -32'sd411359, -32'sd1762144, 32'sd5040171, -32'sd4429975, 32'sd5218876, -32'sd2630390, 32'sd2135751, -32'sd3009006, -32'sd3295607, -32'sd1212959, -32'sd3128181, -32'sd3362096, -32'sd2422704, 32'sd735596, -32'sd356013, -32'sd1957634, 32'sd563538, -32'sd851979, 32'sd1301359, -32'sd2626310, 32'sd4578490, 32'sd1148039, 32'sd1544627, 32'sd3475803, 32'sd638318, 32'sd930100, 32'sd2365481, -32'sd2425020, -32'sd2265769, 32'sd1541827, 32'sd3036500, 32'sd702199, 32'sd1377133, -32'sd533424, 32'sd1332846, 32'sd745447, -32'sd2906638, 32'sd1556972, 32'sd3361777},
        '{32'sd3861493, 32'sd2894947, 32'sd2136487, 32'sd4193496, -32'sd1758985, -32'sd3851208, -32'sd1923210, -32'sd979189, 32'sd418314, 32'sd484804, 32'sd1270559, 32'sd1745747, 32'sd502658, -32'sd1777895, 32'sd648597, -32'sd1195455, -32'sd2494742, -32'sd3664556, -32'sd728502, -32'sd3731555, 32'sd1831831, -32'sd216218, -32'sd3248624, 32'sd3399910, -32'sd1101924, 32'sd2723154, -32'sd2154190, -32'sd5595695, -32'sd1247803, 32'sd435344, -32'sd3742702, 32'sd2488468, 32'sd2790290, -32'sd3085455, 32'sd1900248, -32'sd3433942, -32'sd1365650, -32'sd812079, 32'sd1065725, -32'sd514773, 32'sd338573, 32'sd2725376, -32'sd2796004, -32'sd341138, 32'sd1572220, 32'sd2658928, 32'sd2983485, -32'sd637305, 32'sd301679, -32'sd3619179, 32'sd1651739, -32'sd4365643, 32'sd2645126, -32'sd17553, -32'sd2824425, -32'sd2810344, 32'sd1426993, -32'sd1175365, 32'sd1775940, -32'sd2588391, 32'sd1384918, -32'sd441042, 32'sd584614, 32'sd867831, 32'sd1012440, 32'sd1523034, 32'sd541623, 32'sd1924189, 32'sd176146, 32'sd3072091, 32'sd529213, -32'sd1321840, -32'sd529439, -32'sd548239, 32'sd396184, 32'sd3349003, -32'sd487702, 32'sd5244791, 32'sd2108167, -32'sd3288955, 32'sd2845086, 32'sd4233071, -32'sd2535030, -32'sd2821932, 32'sd476646, -32'sd2377677, 32'sd2104890, 32'sd893982, 32'sd2915113, 32'sd410317, -32'sd1830864, 32'sd4116454, -32'sd988242, -32'sd1774976, 32'sd1996398, -32'sd1345360, -32'sd2363752, 32'sd370869, -32'sd2178562, -32'sd1009734, 32'sd2154325, 32'sd354358, 32'sd5027502, 32'sd3188811, 32'sd1888480, 32'sd2693470, 32'sd499897, -32'sd2226475, -32'sd3484856, 32'sd3286290, 32'sd3468721, -32'sd2621542, -32'sd852229, 32'sd2053240, 32'sd1712827, 32'sd2568903, -32'sd3163051, -32'sd188576, 32'sd2613120, 32'sd1602557, 32'sd2117023, 32'sd1101134, -32'sd3659203, 32'sd952128, 32'sd113588, 32'sd368055, -32'sd1672869, -32'sd1097842},
        '{-32'sd4110200, 32'sd1436701, 32'sd2381429, 32'sd3506336, -32'sd3712536, 32'sd2268550, 32'sd2757973, 32'sd1842431, -32'sd4141733, 32'sd1268724, -32'sd1348752, -32'sd244113, 32'sd3052548, 32'sd851110, -32'sd710191, 32'sd3981119, -32'sd296715, -32'sd2539252, 32'sd1187329, -32'sd5015680, -32'sd2203298, 32'sd3491861, -32'sd1660113, 32'sd444559, -32'sd289021, -32'sd2530404, 32'sd1805082, -32'sd1319172, -32'sd170758, 32'sd940507, -32'sd2377731, 32'sd3310706, 32'sd394300, -32'sd2447547, 32'sd1505545, 32'sd3927076, -32'sd860212, 32'sd3095245, 32'sd1080770, -32'sd2364512, 32'sd143813, 32'sd199174, 32'sd2922194, 32'sd1639974, -32'sd4156798, 32'sd1103195, 32'sd1165021, -32'sd744315, 32'sd717950, 32'sd753032, -32'sd760031, -32'sd365464, 32'sd1793694, -32'sd1021117, -32'sd4473399, 32'sd301976, 32'sd3327791, 32'sd3661592, -32'sd2848045, -32'sd1011571, 32'sd1122870, 32'sd237930, -32'sd2674046, -32'sd211291, -32'sd983835, 32'sd3070900, -32'sd817814, -32'sd1097983, -32'sd1878409, 32'sd1574518, 32'sd2859750, 32'sd530743, -32'sd1426106, -32'sd2572096, -32'sd256823, 32'sd1456641, 32'sd1849715, 32'sd3065862, -32'sd3284966, -32'sd1608277, -32'sd3019346, 32'sd95283, 32'sd2740971, -32'sd435646, 32'sd1270800, 32'sd3126458, -32'sd811642, 32'sd2062541, 32'sd1944377, -32'sd2618918, 32'sd1026256, -32'sd1669509, 32'sd923144, 32'sd864505, -32'sd2672491, 32'sd1594862, 32'sd1116114, 32'sd805859, -32'sd141045, -32'sd2164299, 32'sd2303158, 32'sd1997183, 32'sd2638869, 32'sd2511370, -32'sd2956519, 32'sd353972, 32'sd2700142, 32'sd258585, -32'sd2699113, -32'sd1349041, 32'sd2929138, 32'sd1185878, -32'sd4523066, 32'sd5783193, 32'sd1887124, -32'sd2155109, -32'sd1802084, -32'sd694400, 32'sd1693847, -32'sd2470708, 32'sd2659787, 32'sd68867, -32'sd1223120, 32'sd1147592, 32'sd1533447, 32'sd1121694, -32'sd2079079, -32'sd209216},
        '{32'sd236723, 32'sd2751948, 32'sd1707947, -32'sd3648562, -32'sd709047, 32'sd2041370, -32'sd5387550, -32'sd429682, 32'sd3755630, -32'sd3628424, 32'sd3878431, 32'sd452873, -32'sd2629326, 32'sd1780758, 32'sd2232578, -32'sd551799, 32'sd2667757, 32'sd1072325, 32'sd353676, -32'sd1885702, 32'sd562153, 32'sd517671, 32'sd4324794, 32'sd2263691, -32'sd2529173, -32'sd390401, -32'sd2586740, -32'sd1163520, -32'sd296320, 32'sd3163560, 32'sd1347696, 32'sd1733495, -32'sd2742365, 32'sd1922200, -32'sd3044251, 32'sd1152616, -32'sd3552651, -32'sd2386860, -32'sd1767430, 32'sd2387137, -32'sd1358464, 32'sd246595, 32'sd1389840, 32'sd2740503, -32'sd3416319, 32'sd1026095, -32'sd3209444, -32'sd454625, -32'sd2834037, 32'sd2624154, -32'sd911035, 32'sd1762636, -32'sd1017597, -32'sd980555, 32'sd1294532, 32'sd2463824, -32'sd2965837, 32'sd867116, -32'sd2953695, 32'sd2038999, -32'sd235466, 32'sd346484, -32'sd810800, 32'sd2902388, 32'sd695850, -32'sd474003, -32'sd1391190, -32'sd1962324, -32'sd3310649, -32'sd2379734, -32'sd2931253, -32'sd1387962, 32'sd2361556, -32'sd2464824, 32'sd4194308, -32'sd2460387, -32'sd988505, 32'sd591870, 32'sd1407049, 32'sd1023120, 32'sd2610683, -32'sd2526129, -32'sd438533, 32'sd748521, 32'sd42407, -32'sd343291, -32'sd2946055, -32'sd402979, -32'sd549288, 32'sd3027920, 32'sd1138503, 32'sd548989, 32'sd1866829, 32'sd2166575, 32'sd2162048, 32'sd2723451, 32'sd586981, 32'sd2718077, 32'sd948633, -32'sd932622, -32'sd2331670, -32'sd2635480, -32'sd3751549, 32'sd264396, -32'sd2289342, -32'sd3726144, 32'sd1605840, 32'sd2441708, 32'sd1020646, -32'sd1160060, -32'sd2539253, -32'sd1789250, 32'sd4245880, -32'sd3701267, 32'sd1603128, -32'sd941446, 32'sd1907297, 32'sd930815, -32'sd1037276, -32'sd3844317, 32'sd2419719, 32'sd885359, 32'sd3111817, -32'sd3341965, 32'sd2332714, 32'sd2178379, -32'sd2323318, 32'sd4088451},
        '{-32'sd4686891, 32'sd3100056, -32'sd1953307, -32'sd3899553, -32'sd534245, -32'sd520080, 32'sd1849137, 32'sd2613192, -32'sd3034608, 32'sd1166270, -32'sd1254372, -32'sd2508695, 32'sd168529, 32'sd3653209, 32'sd1147644, 32'sd3427658, -32'sd1512683, 32'sd912693, 32'sd1289017, -32'sd1560813, 32'sd497837, 32'sd490636, 32'sd1303027, 32'sd1978875, 32'sd3634689, 32'sd2481101, 32'sd387483, 32'sd3781532, 32'sd1895001, 32'sd1749951, -32'sd355018, -32'sd3380021, -32'sd2953642, -32'sd733870, -32'sd881470, -32'sd2725718, -32'sd3826724, -32'sd1184646, -32'sd3928876, -32'sd2932367, -32'sd1080859, 32'sd11834, 32'sd130064, 32'sd629893, -32'sd2249903, -32'sd52790, 32'sd2682505, -32'sd392146, -32'sd1405496, 32'sd1843961, 32'sd2213238, 32'sd2452260, 32'sd206523, 32'sd950550, 32'sd1686218, 32'sd2899730, -32'sd1725763, 32'sd1494345, 32'sd5707008, -32'sd85437, -32'sd267232, 32'sd2616396, -32'sd1311781, 32'sd2262640, 32'sd2129038, 32'sd1167470, -32'sd1729355, 32'sd2125418, -32'sd2496125, 32'sd2248296, -32'sd1358512, 32'sd4313895, 32'sd2865052, -32'sd3057684, -32'sd918629, -32'sd1156532, -32'sd1425600, -32'sd1237018, -32'sd1136979, 32'sd3036959, -32'sd2341412, 32'sd2267777, -32'sd1184599, -32'sd1058985, -32'sd1548913, -32'sd594268, -32'sd310710, 32'sd4379571, -32'sd2968869, -32'sd2223986, 32'sd1173968, 32'sd2028797, -32'sd2315585, 32'sd820077, 32'sd63281, -32'sd735651, -32'sd2508464, -32'sd2941183, 32'sd2017987, 32'sd2607130, -32'sd1132642, -32'sd2379444, -32'sd2947784, -32'sd1903975, -32'sd21811, 32'sd4534745, -32'sd3499981, 32'sd132679, 32'sd2613150, -32'sd4988989, -32'sd2861010, -32'sd3810836, -32'sd3030346, 32'sd54670, 32'sd3074960, 32'sd3113327, 32'sd1102969, 32'sd3359349, -32'sd2315515, -32'sd2632711, 32'sd1041696, -32'sd4495555, 32'sd2402699, -32'sd1678326, -32'sd1736129, 32'sd1456797, -32'sd1103239, -32'sd1914238},
        '{32'sd856039, 32'sd3086456, 32'sd2013224, -32'sd1412345, 32'sd1275720, -32'sd2011101, 32'sd4160305, -32'sd831439, -32'sd2821390, -32'sd2924908, -32'sd1312043, -32'sd110936, 32'sd2952856, -32'sd2664543, 32'sd607394, -32'sd479966, 32'sd3062501, -32'sd2050403, 32'sd1191483, -32'sd117447, -32'sd1228625, -32'sd3669145, -32'sd775898, -32'sd1411707, -32'sd1737960, -32'sd3119975, 32'sd538403, 32'sd3182059, 32'sd2023028, -32'sd2629911, -32'sd1754581, 32'sd649292, 32'sd4753079, 32'sd3147025, 32'sd2726763, -32'sd2643625, 32'sd2058962, -32'sd2867038, -32'sd2740293, 32'sd913644, -32'sd1131420, -32'sd2095467, -32'sd2170755, 32'sd1896717, 32'sd939068, 32'sd2382962, 32'sd939887, 32'sd2367744, 32'sd3026608, -32'sd418552, -32'sd2041890, 32'sd1916739, 32'sd1931, -32'sd2199956, -32'sd1214693, 32'sd341428, 32'sd847114, 32'sd2354390, -32'sd90668, -32'sd3123286, -32'sd4016638, -32'sd2606929, 32'sd3696165, 32'sd772762, -32'sd1435502, -32'sd5483555, -32'sd2715288, -32'sd2224385, 32'sd4043255, 32'sd1806584, 32'sd3765248, 32'sd3269768, 32'sd297033, -32'sd2763407, -32'sd61534, 32'sd897418, -32'sd677357, 32'sd873337, -32'sd2030871, 32'sd1489152, 32'sd2161038, 32'sd2149971, -32'sd2587407, 32'sd2325778, -32'sd5343801, -32'sd2293798, 32'sd2503453, -32'sd51735, -32'sd1814661, -32'sd1081715, 32'sd2180598, -32'sd1715556, 32'sd2239265, 32'sd983149, -32'sd587929, -32'sd2667054, 32'sd1758763, -32'sd764451, -32'sd2050031, 32'sd2109038, -32'sd2797305, 32'sd1717921, -32'sd1114266, 32'sd3669241, -32'sd3094904, -32'sd4193058, 32'sd3685219, 32'sd2323883, 32'sd952184, -32'sd278443, -32'sd2929131, 32'sd2430441, 32'sd2165960, -32'sd653940, -32'sd1702963, 32'sd2074811, -32'sd1169214, -32'sd633045, 32'sd2199802, 32'sd1402988, 32'sd1736693, 32'sd1365198, -32'sd3014161, -32'sd2532468, -32'sd700966, -32'sd2240977, 32'sd3114415, 32'sd1075620},
        '{32'sd2044146, -32'sd781724, -32'sd2314524, 32'sd2291887, 32'sd340592, 32'sd1415015, 32'sd146344, 32'sd347698, -32'sd248336, 32'sd3218612, 32'sd2363482, 32'sd2068437, 32'sd359063, 32'sd2787997, 32'sd3613532, -32'sd695046, 32'sd4367543, 32'sd135774, -32'sd195395, 32'sd2246465, -32'sd831185, 32'sd1088708, -32'sd1480664, -32'sd1695847, -32'sd1238195, 32'sd1350572, 32'sd2887261, 32'sd1016811, 32'sd403827, 32'sd1082012, 32'sd771989, 32'sd2179942, 32'sd577734, -32'sd950620, -32'sd2882284, 32'sd2399972, -32'sd1325547, -32'sd2659253, 32'sd1428300, 32'sd544580, -32'sd1979338, -32'sd2398119, 32'sd1029411, 32'sd2610761, -32'sd3192318, -32'sd4280073, 32'sd2763169, -32'sd1246253, -32'sd2026569, 32'sd1207851, -32'sd3632608, 32'sd4269961, -32'sd2337636, -32'sd3487337, 32'sd1948133, 32'sd1013198, -32'sd934125, -32'sd2221335, 32'sd613724, 32'sd2054946, -32'sd5164099, -32'sd3407774, -32'sd1063318, -32'sd1185667, -32'sd213894, -32'sd3357078, 32'sd3243720, 32'sd1101961, 32'sd2379722, 32'sd1532818, -32'sd1171663, 32'sd4186593, 32'sd70931, -32'sd788755, -32'sd1582399, 32'sd2297773, -32'sd502350, 32'sd2589191, -32'sd39071, 32'sd1596407, 32'sd245624, 32'sd190075, 32'sd2015089, 32'sd4573870, 32'sd2972452, -32'sd367684, 32'sd3927459, 32'sd487522, -32'sd1924794, -32'sd548432, -32'sd3151616, 32'sd944777, 32'sd3008716, 32'sd2177179, -32'sd1436617, 32'sd1033968, 32'sd1642238, -32'sd2028805, -32'sd777812, -32'sd3656592, -32'sd2867256, -32'sd2705758, -32'sd2481773, -32'sd3400312, -32'sd1445924, 32'sd1203830, 32'sd3419625, -32'sd1764766, -32'sd4064755, 32'sd997107, 32'sd2256511, 32'sd2843376, 32'sd1494022, 32'sd1451754, 32'sd602769, -32'sd1245712, 32'sd3136271, 32'sd1387193, -32'sd1153663, -32'sd1496112, 32'sd2161770, -32'sd2439938, -32'sd919107, -32'sd3919113, -32'sd863800, -32'sd1386204, -32'sd1017385, 32'sd1344746},
        '{-32'sd818907, 32'sd5086282, 32'sd1019487, -32'sd1276451, -32'sd2549549, 32'sd1905882, 32'sd1344262, 32'sd1555037, -32'sd2762358, 32'sd1467958, 32'sd725596, 32'sd779577, 32'sd1907553, 32'sd4508762, 32'sd166793, 32'sd2201260, 32'sd2964558, 32'sd2973414, 32'sd3078099, 32'sd3978871, 32'sd94370, 32'sd5074820, 32'sd315848, -32'sd3513453, 32'sd2691140, 32'sd397698, 32'sd3113415, 32'sd1663817, -32'sd2981340, -32'sd185092, 32'sd3257569, 32'sd2957433, -32'sd1057847, 32'sd1249327, -32'sd390216, 32'sd2542947, 32'sd241900, -32'sd313754, 32'sd2623940, -32'sd1927940, -32'sd2186381, 32'sd2297790, 32'sd964739, 32'sd3744625, 32'sd2945254, -32'sd1143856, -32'sd1720357, -32'sd1892210, -32'sd1247871, -32'sd490835, 32'sd1623260, 32'sd2132468, -32'sd1980577, -32'sd3000564, 32'sd538200, -32'sd9094, -32'sd311291, 32'sd2026667, 32'sd2174968, 32'sd3481560, -32'sd1199263, 32'sd597021, 32'sd255400, -32'sd3516594, 32'sd329763, -32'sd168603, 32'sd1502681, -32'sd2707640, 32'sd3990458, 32'sd1866863, 32'sd929869, 32'sd2857332, -32'sd139511, 32'sd3725769, 32'sd1653122, -32'sd1295378, -32'sd271, 32'sd1576990, -32'sd2496805, 32'sd3418115, -32'sd552520, 32'sd180216, 32'sd5428879, -32'sd1163054, 32'sd37011, -32'sd685286, -32'sd546700, 32'sd2384998, -32'sd2418550, 32'sd1548801, -32'sd2960214, 32'sd615626, -32'sd1349753, -32'sd2013787, 32'sd642363, 32'sd2725127, 32'sd948527, -32'sd1674527, 32'sd1789051, 32'sd4337370, -32'sd3263805, -32'sd4191294, -32'sd3019337, 32'sd1569518, -32'sd2939930, 32'sd4099822, -32'sd704533, 32'sd1372141, 32'sd2529271, -32'sd59054, -32'sd2500622, -32'sd1004002, 32'sd684882, 32'sd3570278, -32'sd496364, -32'sd3705034, 32'sd3177859, 32'sd944274, 32'sd2687481, 32'sd1797786, -32'sd914845, -32'sd3577429, 32'sd1296717, 32'sd2130495, 32'sd1789841, 32'sd2711854, 32'sd1943575, 32'sd1418427},
        '{-32'sd744142, -32'sd418175, -32'sd1547522, -32'sd5056806, -32'sd1919296, -32'sd1222357, 32'sd2648257, -32'sd1543061, -32'sd3895866, -32'sd2427027, -32'sd1381, -32'sd96131, -32'sd5143463, -32'sd626803, 32'sd1148618, 32'sd689620, 32'sd5107296, 32'sd62161, 32'sd635041, 32'sd1844871, -32'sd2915852, 32'sd180507, -32'sd5178585, 32'sd2500781, -32'sd2323185, 32'sd1869701, -32'sd2153090, -32'sd285683, 32'sd1058523, 32'sd619070, -32'sd651358, -32'sd1499276, -32'sd4399342, -32'sd651835, 32'sd3555040, -32'sd1353332, -32'sd3837005, -32'sd1689128, -32'sd460583, -32'sd876954, -32'sd3208593, 32'sd1136954, 32'sd216070, -32'sd809819, 32'sd4471554, -32'sd46081, -32'sd6532448, -32'sd261993, -32'sd4033177, -32'sd2494236, 32'sd3618183, -32'sd4103318, -32'sd2291305, 32'sd680698, 32'sd1934576, -32'sd2820920, -32'sd892461, 32'sd2727666, 32'sd230354, -32'sd1168460, 32'sd3842557, 32'sd2126696, -32'sd4086559, -32'sd613448, 32'sd3164468, -32'sd1530098, 32'sd1453500, 32'sd299642, -32'sd639212, -32'sd1718325, 32'sd1087379, -32'sd297675, 32'sd194528, 32'sd2716245, -32'sd1445246, 32'sd1563641, -32'sd603521, -32'sd2611747, -32'sd652583, 32'sd946271, -32'sd93385, -32'sd328237, 32'sd1966357, -32'sd1799555, -32'sd337674, 32'sd3304905, 32'sd1805536, 32'sd3721014, -32'sd1954315, -32'sd2420821, 32'sd2337628, -32'sd515450, -32'sd3618884, -32'sd2487025, -32'sd317340, 32'sd742077, 32'sd632885, -32'sd3515372, -32'sd83520, 32'sd3120187, -32'sd4466006, 32'sd22190, -32'sd3916077, 32'sd544585, -32'sd1519005, -32'sd412449, -32'sd3390627, 32'sd937501, 32'sd434174, -32'sd80042, -32'sd1781015, -32'sd2662612, 32'sd3458009, 32'sd3187653, -32'sd1146864, -32'sd2182350, 32'sd1336405, 32'sd1354308, 32'sd2131959, 32'sd317239, 32'sd248385, -32'sd533094, 32'sd1989032, -32'sd1242863, -32'sd2655631, 32'sd403305, 32'sd1462884, 32'sd2329149},
        '{32'sd1262403, -32'sd656556, 32'sd780695, 32'sd464560, -32'sd1368946, -32'sd1542272, -32'sd1588900, -32'sd1452449, -32'sd2820199, 32'sd2471082, -32'sd297101, 32'sd1649386, 32'sd2894095, -32'sd2386686, -32'sd2490223, 32'sd1925876, 32'sd2745637, -32'sd4536795, -32'sd669340, 32'sd588016, -32'sd3793914, -32'sd980356, -32'sd2693137, 32'sd223754, -32'sd2369581, -32'sd2126604, 32'sd3386940, 32'sd137525, -32'sd3854117, 32'sd1762935, 32'sd315591, -32'sd3599170, -32'sd1105630, -32'sd830858, 32'sd3397812, -32'sd2400252, 32'sd3507352, -32'sd2052650, 32'sd2128757, 32'sd460989, 32'sd2664124, 32'sd2784094, 32'sd3487558, 32'sd685857, 32'sd3185026, 32'sd2299545, 32'sd4065617, 32'sd23894, 32'sd1528386, 32'sd2028628, 32'sd6437, -32'sd1337604, 32'sd895319, 32'sd2691642, -32'sd292988, -32'sd2595011, 32'sd4015861, -32'sd2084922, -32'sd3240516, -32'sd321682, -32'sd1364530, -32'sd1805410, 32'sd1941117, 32'sd1012210, 32'sd2402930, 32'sd1311176, 32'sd211123, 32'sd3326466, -32'sd1046508, -32'sd3891717, 32'sd1048184, 32'sd1490391, 32'sd501819, 32'sd1579569, 32'sd1903773, 32'sd2688861, 32'sd1803988, 32'sd4212474, -32'sd1464501, 32'sd1868087, -32'sd3686235, -32'sd293003, 32'sd1551927, 32'sd3001948, 32'sd1776754, -32'sd3128993, -32'sd1859416, -32'sd4215064, -32'sd1675397, 32'sd1054019, 32'sd1553877, -32'sd1739960, 32'sd786978, 32'sd960093, 32'sd1121174, -32'sd3610524, -32'sd390455, 32'sd2318243, 32'sd1636909, 32'sd2142510, 32'sd961794, 32'sd1747, -32'sd2082103, -32'sd1505227, -32'sd2981132, -32'sd1305903, -32'sd3492805, 32'sd1874151, 32'sd1805082, -32'sd841641, 32'sd3238512, -32'sd2403566, -32'sd730890, 32'sd1101631, 32'sd3240286, 32'sd2309406, -32'sd2982721, 32'sd2845309, 32'sd49579, 32'sd547823, 32'sd2960877, 32'sd2479623, 32'sd791597, -32'sd3901134, 32'sd3572327, -32'sd2053221, 32'sd4364843, 32'sd857504},
        '{-32'sd1662026, -32'sd1302138, -32'sd3278951, 32'sd2525857, 32'sd727245, -32'sd1007591, -32'sd3508332, 32'sd2814534, 32'sd2284593, 32'sd403859, -32'sd1771607, -32'sd875899, -32'sd767798, -32'sd1688123, -32'sd3785662, -32'sd3037192, 32'sd2852215, -32'sd3911584, 32'sd461148, -32'sd249957, -32'sd688511, 32'sd935203, 32'sd1911736, 32'sd1489550, -32'sd4353181, 32'sd2872849, 32'sd640734, -32'sd4776267, 32'sd2058505, 32'sd2687403, -32'sd1478361, -32'sd87910, 32'sd2033266, 32'sd227318, -32'sd1074137, -32'sd2425667, 32'sd706761, 32'sd1296114, 32'sd718703, 32'sd1406402, 32'sd864595, 32'sd2379093, 32'sd3009950, 32'sd1411309, -32'sd156281, 32'sd5074629, -32'sd1193440, -32'sd387974, -32'sd1363473, -32'sd2100339, 32'sd942329, -32'sd403351, -32'sd1771964, 32'sd2588821, -32'sd2058471, 32'sd136735, -32'sd2608767, 32'sd396278, 32'sd1294389, 32'sd3983861, -32'sd1838359, 32'sd2658418, 32'sd2306808, 32'sd1599331, 32'sd899334, 32'sd71083, 32'sd1413482, -32'sd496221, -32'sd1658031, -32'sd1427909, -32'sd4535682, -32'sd5111516, -32'sd2807604, 32'sd3061319, -32'sd1510585, 32'sd4037208, 32'sd2964887, -32'sd5168358, 32'sd3712917, -32'sd1250552, -32'sd310778, 32'sd3068737, 32'sd2817715, 32'sd2072913, 32'sd5326658, 32'sd2641801, -32'sd1517853, -32'sd1964521, 32'sd1017650, 32'sd1945977, -32'sd841566, 32'sd2131997, -32'sd642970, 32'sd1081217, 32'sd921367, -32'sd2065071, -32'sd716594, -32'sd132861, 32'sd2507887, 32'sd3459938, -32'sd2082244, -32'sd3163713, 32'sd1621202, 32'sd2826827, -32'sd1199056, -32'sd2416372, -32'sd1843947, -32'sd2841609, 32'sd1724912, 32'sd1894991, 32'sd1482076, -32'sd5503295, -32'sd3980780, 32'sd3127916, -32'sd627315, -32'sd3301478, 32'sd1511851, 32'sd908565, 32'sd815492, 32'sd312107, -32'sd5120451, 32'sd1384589, -32'sd515603, -32'sd2090200, -32'sd3366295, -32'sd3612831, -32'sd1314353, 32'sd885478},
        '{32'sd1243339, -32'sd6204614, -32'sd336172, 32'sd3429327, 32'sd2486078, -32'sd4616010, -32'sd762550, 32'sd659552, 32'sd2532024, -32'sd253089, -32'sd1255089, 32'sd837192, 32'sd456857, 32'sd1961258, 32'sd593038, 32'sd191291, 32'sd358961, 32'sd2514136, -32'sd509296, 32'sd3936192, 32'sd2415432, -32'sd1185111, -32'sd331466, 32'sd1912789, -32'sd7024205, -32'sd1502850, -32'sd4636978, -32'sd1779233, -32'sd3101473, 32'sd486790, -32'sd2885902, 32'sd1428367, -32'sd1260081, 32'sd2973084, 32'sd4115998, -32'sd1450925, -32'sd1266164, -32'sd4491492, 32'sd2389884, 32'sd4862487, 32'sd1002996, 32'sd965222, 32'sd3049459, -32'sd4590905, 32'sd1773973, -32'sd1086710, -32'sd2352877, -32'sd2050361, -32'sd1213083, 32'sd1981764, -32'sd2609615, -32'sd3339290, -32'sd2829713, -32'sd275854, 32'sd1650008, 32'sd2549961, -32'sd2487380, 32'sd109459, -32'sd3024331, -32'sd2570185, 32'sd3585417, 32'sd2431513, -32'sd607407, 32'sd3920189, -32'sd366832, -32'sd3550680, 32'sd95696, 32'sd2571575, -32'sd3341310, -32'sd670963, -32'sd1757665, 32'sd2022771, 32'sd4802687, 32'sd920847, -32'sd2311452, -32'sd5755403, -32'sd1131953, 32'sd1547760, 32'sd2184522, 32'sd262383, -32'sd72191, -32'sd3784453, -32'sd916630, 32'sd1106324, 32'sd740016, -32'sd756203, -32'sd351463, -32'sd1687104, -32'sd1220479, -32'sd3286081, -32'sd2322772, -32'sd1201940, 32'sd2662523, -32'sd2448383, 32'sd3086968, 32'sd2153964, -32'sd778609, 32'sd2801704, 32'sd2368486, -32'sd4133566, -32'sd2520776, 32'sd2461967, -32'sd3062481, -32'sd3126995, -32'sd1501769, -32'sd3573622, -32'sd497832, -32'sd4225905, 32'sd1338192, 32'sd4197582, 32'sd788212, 32'sd287692, 32'sd5258069, -32'sd1196984, -32'sd1219782, -32'sd2377418, 32'sd2973358, -32'sd2294302, 32'sd1197852, 32'sd1554150, -32'sd1236338, 32'sd1648571, 32'sd1834898, 32'sd74344, 32'sd453143, 32'sd40371, 32'sd1622586, 32'sd2533240},
        '{32'sd2932242, -32'sd2534414, 32'sd356217, 32'sd2444400, -32'sd2372073, -32'sd1709524, 32'sd2502426, -32'sd327754, -32'sd2783805, -32'sd2398474, -32'sd512656, -32'sd818325, -32'sd3684497, 32'sd1621718, 32'sd2163466, -32'sd5929405, 32'sd2756878, -32'sd2707006, 32'sd161296, 32'sd2510426, 32'sd1949055, 32'sd390738, -32'sd1134658, -32'sd137537, -32'sd2921965, 32'sd456048, -32'sd2571572, -32'sd940456, -32'sd3742310, -32'sd4996117, 32'sd353389, -32'sd2633631, -32'sd1724461, 32'sd68202, 32'sd845408, -32'sd5442308, 32'sd2813711, -32'sd698761, 32'sd775414, 32'sd4885847, -32'sd1708769, 32'sd2177735, -32'sd2719102, -32'sd1166930, 32'sd3236584, 32'sd2910537, -32'sd5492460, -32'sd4550370, -32'sd2437879, -32'sd3556267, -32'sd3381396, -32'sd1676416, -32'sd560357, 32'sd1339542, 32'sd5292945, -32'sd1957703, 32'sd342988, 32'sd1053816, 32'sd2659864, 32'sd3538394, 32'sd137136, 32'sd3281397, 32'sd1692429, 32'sd4384318, -32'sd414031, -32'sd174441, -32'sd2484332, -32'sd1424171, -32'sd2043902, 32'sd1107866, 32'sd3231083, -32'sd3041706, -32'sd1738833, -32'sd3222872, -32'sd1257463, -32'sd588529, -32'sd314161, 32'sd669036, 32'sd1397612, 32'sd780199, -32'sd952049, 32'sd1889476, 32'sd3586252, -32'sd1975816, 32'sd2096184, 32'sd719605, 32'sd1856648, 32'sd102347, 32'sd1749318, -32'sd2797527, 32'sd3539086, 32'sd567454, -32'sd3611036, -32'sd2751741, -32'sd1323866, -32'sd85293, -32'sd3251602, 32'sd340306, -32'sd1306985, 32'sd2946598, 32'sd537040, -32'sd722055, -32'sd2382584, 32'sd1094518, -32'sd1057244, -32'sd2416827, -32'sd1940833, 32'sd1726669, 32'sd1857718, -32'sd1462805, 32'sd3068838, -32'sd2965048, 32'sd1490361, 32'sd2959219, -32'sd1228472, 32'sd885882, 32'sd532513, 32'sd4381139, 32'sd1430311, 32'sd359186, -32'sd2128667, -32'sd141675, 32'sd549752, -32'sd2658378, -32'sd2305015, -32'sd1553190, -32'sd1736175, -32'sd162654},
        '{-32'sd298057, 32'sd1837286, -32'sd3301189, 32'sd2356918, -32'sd3925241, -32'sd957659, -32'sd255778, -32'sd4220911, -32'sd1513870, 32'sd3318859, 32'sd1769915, 32'sd969616, 32'sd309133, -32'sd108352, 32'sd2035279, 32'sd3307638, 32'sd865361, -32'sd1665050, -32'sd945731, -32'sd4157103, -32'sd652965, -32'sd3643287, 32'sd1445244, -32'sd575125, 32'sd4081942, 32'sd2432508, -32'sd1152623, 32'sd2448669, -32'sd1354306, -32'sd1176524, 32'sd1011990, -32'sd3236771, 32'sd3307511, -32'sd2077892, 32'sd3917842, -32'sd1975192, 32'sd3561074, 32'sd1890535, 32'sd1824963, 32'sd2848873, 32'sd1426295, -32'sd1252097, 32'sd1322394, -32'sd760955, -32'sd5059791, 32'sd2805361, 32'sd1427612, 32'sd1381942, 32'sd1928498, -32'sd3412610, -32'sd108197, -32'sd598000, 32'sd1828703, -32'sd2197885, 32'sd126373, -32'sd2280885, 32'sd1755763, 32'sd774721, 32'sd985146, -32'sd4293491, -32'sd18762, 32'sd1431589, 32'sd994746, -32'sd1848042, -32'sd1291481, 32'sd265851, 32'sd475343, 32'sd3418934, -32'sd3161582, 32'sd669473, -32'sd1055649, 32'sd4602195, 32'sd5206364, -32'sd3041232, 32'sd2628809, -32'sd943798, 32'sd2931559, -32'sd384618, 32'sd1069114, -32'sd2206429, -32'sd3905686, 32'sd615264, -32'sd3408867, -32'sd3265922, -32'sd2368140, 32'sd191885, 32'sd1312346, -32'sd492708, 32'sd1974079, 32'sd3295699, 32'sd590862, 32'sd1450869, 32'sd4066960, -32'sd2550267, 32'sd2101999, 32'sd1015133, 32'sd1463803, 32'sd1541074, 32'sd440836, -32'sd3232978, -32'sd44802, -32'sd1286798, -32'sd1385680, -32'sd77853, 32'sd951944, -32'sd1940311, 32'sd187043, -32'sd2764149, 32'sd71950, 32'sd905012, 32'sd2017699, -32'sd2038890, -32'sd4509869, -32'sd3920099, 32'sd89226, 32'sd405542, -32'sd88469, -32'sd470496, -32'sd1908988, 32'sd1275491, -32'sd1332978, -32'sd2658510, 32'sd1811255, -32'sd2068143, 32'sd3274646, 32'sd2743941, -32'sd1877049, 32'sd2296254},
        '{32'sd1956486, 32'sd514575, 32'sd543032, 32'sd1109142, -32'sd635780, 32'sd2852430, -32'sd303422, 32'sd4310796, 32'sd339595, -32'sd2199872, -32'sd2489977, 32'sd1957863, 32'sd2795695, -32'sd3008108, -32'sd940464, -32'sd1203392, -32'sd259474, 32'sd3421471, 32'sd1082754, 32'sd571143, 32'sd4882519, 32'sd4064069, -32'sd1236863, 32'sd808951, 32'sd2237791, -32'sd2382081, -32'sd3565875, 32'sd2744840, -32'sd2521927, -32'sd3167202, -32'sd94522, -32'sd993594, -32'sd2759706, -32'sd2917177, -32'sd225508, 32'sd3106857, -32'sd78951, 32'sd2739703, -32'sd2014495, -32'sd1480361, 32'sd1641281, 32'sd1437739, -32'sd969882, 32'sd133975, -32'sd431745, -32'sd822493, 32'sd3415095, -32'sd2640705, -32'sd232368, 32'sd2272544, -32'sd1621219, -32'sd2471352, 32'sd14271, 32'sd2355120, -32'sd1036909, -32'sd1548093, 32'sd3630969, 32'sd1235942, 32'sd613902, -32'sd3609414, -32'sd1696739, -32'sd2251865, -32'sd3438807, 32'sd1656135, 32'sd5168932, 32'sd670305, -32'sd2184626, 32'sd688934, -32'sd3859661, 32'sd757978, -32'sd1339637, 32'sd2365892, 32'sd1302538, 32'sd3228626, 32'sd1044400, 32'sd996843, -32'sd490105, 32'sd2918777, 32'sd1850146, -32'sd3101350, 32'sd2091183, -32'sd633846, 32'sd194728, -32'sd1715216, -32'sd2796456, -32'sd2483588, 32'sd673088, 32'sd4104696, -32'sd1280771, -32'sd1769348, -32'sd1711207, -32'sd3412417, -32'sd4046201, 32'sd2876860, 32'sd2123999, -32'sd2160091, 32'sd508945, 32'sd3477693, 32'sd2180239, -32'sd1369228, 32'sd1659933, -32'sd1116586, 32'sd119385, 32'sd3635030, -32'sd5104853, -32'sd1936831, 32'sd2152083, 32'sd921492, -32'sd1808498, 32'sd1430493, -32'sd5148333, -32'sd767006, 32'sd2979172, -32'sd83417, -32'sd2011379, 32'sd3582330, 32'sd2364265, -32'sd298599, 32'sd1464811, -32'sd4196426, 32'sd4349053, 32'sd2703500, 32'sd1221786, 32'sd695622, -32'sd927704, 32'sd1817984, -32'sd1226668, -32'sd861831},
        '{-32'sd1660505, -32'sd1020730, -32'sd1017928, -32'sd1453928, -32'sd1193490, 32'sd1613574, -32'sd2545565, -32'sd2243745, -32'sd559191, 32'sd3579785, 32'sd2850001, 32'sd862731, 32'sd343819, 32'sd873651, -32'sd901205, 32'sd1621472, -32'sd743143, -32'sd2214171, -32'sd3186192, 32'sd1334168, -32'sd2049694, 32'sd3030609, -32'sd3133757, 32'sd755032, -32'sd2743013, 32'sd2112724, 32'sd1697218, -32'sd2340001, 32'sd2794306, -32'sd2930358, -32'sd68876, 32'sd4171332, -32'sd1384587, -32'sd3333368, -32'sd2491152, -32'sd779145, 32'sd1241694, -32'sd143218, -32'sd2982887, -32'sd2392791, 32'sd2245260, -32'sd2618941, -32'sd4896328, 32'sd756284, 32'sd1597033, 32'sd1009774, 32'sd4853987, -32'sd1921520, -32'sd4317693, -32'sd2483846, 32'sd4599566, 32'sd2434740, -32'sd4115669, -32'sd2548878, 32'sd3395781, 32'sd14932, 32'sd1589544, 32'sd3350123, 32'sd916329, -32'sd3431017, 32'sd3047082, -32'sd106740, -32'sd2600544, -32'sd97012, -32'sd450784, -32'sd955611, 32'sd941851, 32'sd2892852, -32'sd5541443, -32'sd969387, -32'sd1901787, 32'sd2031724, 32'sd5149860, -32'sd494267, 32'sd107346, -32'sd713384, 32'sd2327875, -32'sd74274, 32'sd2779886, 32'sd3276441, -32'sd4429402, -32'sd2055226, -32'sd2461488, -32'sd2003821, -32'sd951753, 32'sd3168359, -32'sd3063949, 32'sd2960554, 32'sd1635378, -32'sd492852, 32'sd1876020, 32'sd1458568, -32'sd2206262, 32'sd801409, 32'sd78076, 32'sd869587, -32'sd914218, -32'sd3204183, 32'sd1615816, 32'sd384328, 32'sd452116, -32'sd542328, -32'sd2631974, -32'sd3904334, 32'sd1384463, -32'sd1442607, -32'sd91237, 32'sd2203913, -32'sd969443, 32'sd2690729, -32'sd2597253, -32'sd3816493, -32'sd1458240, -32'sd3141101, 32'sd855304, 32'sd3173109, 32'sd2414401, 32'sd1723163, 32'sd254435, 32'sd2324830, -32'sd1704914, 32'sd1878625, -32'sd574003, 32'sd278800, 32'sd571077, 32'sd5103485, 32'sd156093, 32'sd2326240},
        '{32'sd547074, 32'sd2121431, -32'sd35895, 32'sd1756838, -32'sd2651276, -32'sd3199056, -32'sd226874, -32'sd3982781, -32'sd2851179, -32'sd1766145, 32'sd3767161, -32'sd366147, -32'sd307252, -32'sd196123, 32'sd1490680, -32'sd2259491, -32'sd1365194, -32'sd77652, 32'sd467265, -32'sd820441, -32'sd5700057, 32'sd2192165, 32'sd410934, -32'sd2230573, 32'sd658974, 32'sd4555244, 32'sd4060323, 32'sd3571431, 32'sd3201545, -32'sd3999490, -32'sd5266452, 32'sd876438, -32'sd1605157, -32'sd1714571, -32'sd1384678, 32'sd3164093, -32'sd4228083, -32'sd1681849, 32'sd735981, 32'sd825706, 32'sd782956, -32'sd190193, -32'sd715756, 32'sd2957952, 32'sd481081, 32'sd3761136, -32'sd50849, 32'sd1614995, 32'sd2163107, -32'sd708573, 32'sd854804, 32'sd2271667, -32'sd354733, 32'sd3720019, -32'sd106279, 32'sd681909, -32'sd1631058, 32'sd130794, -32'sd432519, 32'sd3624686, 32'sd171020, -32'sd2418513, -32'sd2654918, 32'sd2149939, 32'sd922323, 32'sd2203436, -32'sd1048363, 32'sd61995, -32'sd1534842, 32'sd886939, 32'sd1971605, -32'sd3085607, -32'sd3382743, -32'sd2805691, -32'sd3129483, 32'sd3311323, -32'sd2420585, 32'sd1885128, -32'sd633571, 32'sd468684, -32'sd355547, -32'sd621687, 32'sd607758, -32'sd1642507, 32'sd578607, -32'sd329082, 32'sd513286, -32'sd2355252, -32'sd1611763, -32'sd2267100, 32'sd81627, -32'sd2342004, 32'sd4790466, 32'sd2214458, -32'sd3099256, 32'sd1569410, 32'sd1962749, -32'sd461990, -32'sd84928, -32'sd2747179, 32'sd978657, 32'sd3089483, 32'sd2667373, -32'sd36461, -32'sd2875525, -32'sd2508883, 32'sd1827272, -32'sd1239554, 32'sd2846674, -32'sd881547, -32'sd3880388, -32'sd1100796, -32'sd313358, 32'sd1092622, 32'sd559369, -32'sd1214244, 32'sd774622, -32'sd2956429, -32'sd330681, 32'sd1140290, 32'sd3896467, -32'sd418240, 32'sd1083776, 32'sd648113, -32'sd2583629, 32'sd3251886, 32'sd1044785, 32'sd980955},
        '{-32'sd3597172, -32'sd1479135, 32'sd2270429, 32'sd238125, 32'sd1296525, 32'sd654648, -32'sd3395551, -32'sd169184, 32'sd2497873, -32'sd724921, -32'sd3146235, 32'sd146451, -32'sd3123026, 32'sd3413335, 32'sd1579957, -32'sd2173211, 32'sd730853, 32'sd3984290, -32'sd64649, 32'sd2376272, -32'sd1708996, -32'sd651942, 32'sd5472415, -32'sd480237, 32'sd67243, -32'sd2939907, 32'sd3113272, 32'sd3679620, -32'sd2383293, -32'sd2890608, 32'sd415791, 32'sd1902813, -32'sd1075710, 32'sd175737, -32'sd1979186, -32'sd2992098, -32'sd1024858, -32'sd669391, 32'sd3409193, 32'sd1337898, -32'sd4549288, 32'sd249104, -32'sd3117078, -32'sd4209162, -32'sd1317987, -32'sd321218, 32'sd469229, -32'sd3283204, -32'sd3890094, -32'sd405481, 32'sd208239, 32'sd108513, -32'sd3270449, -32'sd1654144, 32'sd5462041, -32'sd2359717, -32'sd1261287, 32'sd1962859, -32'sd4368995, 32'sd268475, -32'sd1817202, 32'sd409766, -32'sd3511317, 32'sd4481629, -32'sd1891772, -32'sd2742629, 32'sd373877, 32'sd1973998, -32'sd2678321, -32'sd213489, -32'sd3352647, -32'sd2321934, -32'sd574729, -32'sd2261453, 32'sd1852805, -32'sd59110, 32'sd3417755, -32'sd2779374, 32'sd2512091, 32'sd1352773, 32'sd3285673, -32'sd1963498, 32'sd23782, -32'sd4105776, -32'sd93463, 32'sd960915, -32'sd3724898, 32'sd1336174, 32'sd1518603, -32'sd270076, 32'sd2067082, 32'sd1940451, 32'sd413213, 32'sd2417891, 32'sd420938, 32'sd1958128, 32'sd2389911, 32'sd86549, -32'sd926285, 32'sd2046824, -32'sd2169195, 32'sd265576, -32'sd2129444, 32'sd4043185, -32'sd741199, -32'sd3843635, 32'sd2589919, -32'sd28195, 32'sd920829, -32'sd3996343, 32'sd1603724, 32'sd836381, -32'sd168352, 32'sd1513007, -32'sd2118698, 32'sd2225130, 32'sd1704821, 32'sd631889, 32'sd1324556, 32'sd275379, 32'sd2581827, -32'sd1643353, 32'sd738462, 32'sd1098796, -32'sd2616440, 32'sd1836774, -32'sd52022, 32'sd3074535},
        '{32'sd2923896, -32'sd793624, -32'sd2374613, 32'sd90764, -32'sd689791, -32'sd2118077, 32'sd2272848, 32'sd3091693, -32'sd2046694, 32'sd4314503, 32'sd2338583, 32'sd742903, 32'sd1334370, -32'sd2920794, 32'sd385866, 32'sd1010914, 32'sd1361122, -32'sd2293894, 32'sd719200, -32'sd3187385, 32'sd2199470, -32'sd1542765, -32'sd1099069, -32'sd2597445, -32'sd2048297, 32'sd3888408, 32'sd48427, -32'sd2628332, 32'sd1023028, 32'sd3435157, -32'sd2817614, 32'sd562342, 32'sd4872446, 32'sd1305501, 32'sd3263841, -32'sd2155772, -32'sd40375, 32'sd379953, 32'sd1677673, 32'sd820620, 32'sd1302265, -32'sd4715712, -32'sd1545343, -32'sd1813050, -32'sd4604142, 32'sd1688111, 32'sd5105521, -32'sd2597933, 32'sd2430531, -32'sd929299, 32'sd337568, 32'sd157946, -32'sd2814614, -32'sd3291658, -32'sd1229050, 32'sd906121, 32'sd2569859, 32'sd3688900, -32'sd2032504, 32'sd51261, -32'sd1727593, -32'sd3353499, -32'sd121832, 32'sd3209898, -32'sd1178815, 32'sd2232937, 32'sd1324470, 32'sd1297864, 32'sd2851220, -32'sd429159, 32'sd3490740, 32'sd1241446, -32'sd527165, -32'sd611202, -32'sd2329766, 32'sd2554240, 32'sd1725632, 32'sd2410162, 32'sd466877, 32'sd1459643, 32'sd376563, 32'sd2466886, 32'sd1057914, 32'sd1608964, 32'sd1879553, -32'sd2416200, 32'sd744936, 32'sd2230018, 32'sd2557181, -32'sd3326781, 32'sd454953, 32'sd2268675, -32'sd619200, -32'sd3750022, 32'sd3312915, -32'sd2821556, -32'sd2529120, -32'sd518239, -32'sd2792763, 32'sd2480634, -32'sd2996986, -32'sd97596, 32'sd1277890, 32'sd251346, -32'sd877263, 32'sd3574343, -32'sd498953, -32'sd1521105, -32'sd1184343, 32'sd549301, 32'sd2915878, -32'sd442684, 32'sd1986684, 32'sd619764, 32'sd1829869, 32'sd2326926, 32'sd649222, 32'sd327288, -32'sd2074574, 32'sd209257, -32'sd3190021, 32'sd366890, -32'sd2350461, -32'sd551423, -32'sd543040, 32'sd2694658, -32'sd2836549, 32'sd1226481},
        '{32'sd2254963, -32'sd4709810, -32'sd2503828, -32'sd750952, -32'sd3573134, 32'sd346527, -32'sd45169, 32'sd2355603, 32'sd217201, -32'sd3165683, 32'sd3005175, 32'sd4847468, -32'sd1915074, -32'sd384511, -32'sd717086, -32'sd2630614, 32'sd1135627, 32'sd565379, -32'sd2969841, 32'sd905397, -32'sd2104823, 32'sd3785508, -32'sd683101, 32'sd3115730, 32'sd2214332, -32'sd466412, -32'sd3984640, 32'sd273471, -32'sd447149, 32'sd644202, 32'sd3362662, 32'sd3556840, -32'sd5487191, 32'sd2316624, -32'sd1553962, -32'sd967878, -32'sd858158, 32'sd1625162, -32'sd2293247, -32'sd304005, 32'sd328580, 32'sd2602405, -32'sd4635565, -32'sd2587465, 32'sd882828, -32'sd3232606, 32'sd1450952, -32'sd4785370, -32'sd3192558, -32'sd1875625, 32'sd2469974, -32'sd4961184, 32'sd1347701, -32'sd1575329, 32'sd303949, -32'sd912572, -32'sd737411, 32'sd2461077, -32'sd1815831, -32'sd118975, 32'sd105928, 32'sd3033288, -32'sd275735, 32'sd151928, -32'sd2280802, -32'sd2416180, 32'sd4006475, -32'sd2576722, -32'sd5615824, -32'sd151509, -32'sd534202, -32'sd1348049, 32'sd3492083, -32'sd859320, 32'sd4699622, -32'sd2045581, -32'sd1931071, -32'sd664410, -32'sd338001, -32'sd649722, 32'sd3500216, -32'sd4513, -32'sd1372693, 32'sd1964490, 32'sd2179809, 32'sd903991, 32'sd2596407, 32'sd142407, 32'sd434249, 32'sd310024, -32'sd690609, 32'sd2589455, -32'sd4516787, -32'sd1260833, 32'sd1955491, 32'sd4325930, 32'sd5448498, 32'sd3643936, 32'sd3002097, -32'sd2438073, 32'sd642080, -32'sd922563, -32'sd5109818, -32'sd2851200, -32'sd3926663, -32'sd1339421, -32'sd1366491, 32'sd3904919, 32'sd499443, -32'sd136871, -32'sd2794973, 32'sd1129322, -32'sd1044619, 32'sd605455, -32'sd2790731, -32'sd1612808, -32'sd285251, -32'sd3554327, -32'sd238691, 32'sd1981629, 32'sd2625439, 32'sd5245372, 32'sd2345469, 32'sd1974960, 32'sd261699, 32'sd3486133, 32'sd979068, -32'sd1908139},
        '{32'sd556956, -32'sd419213, -32'sd2779913, 32'sd1425410, 32'sd2157280, 32'sd86734, 32'sd3036698, 32'sd376563, 32'sd3027002, -32'sd1059979, 32'sd881289, 32'sd2710148, 32'sd540416, 32'sd2019915, 32'sd1102927, -32'sd1850374, -32'sd2888463, -32'sd1599601, 32'sd972682, -32'sd1967255, 32'sd1393152, -32'sd2641163, 32'sd708474, 32'sd2235253, -32'sd254234, -32'sd381759, -32'sd2292127, -32'sd2009638, -32'sd4045561, 32'sd2953176, 32'sd1907543, 32'sd706065, -32'sd3603750, 32'sd2667144, -32'sd378600, -32'sd4744804, -32'sd838450, -32'sd3738125, -32'sd4261469, -32'sd2278232, 32'sd899658, 32'sd1528321, -32'sd3169950, -32'sd15110, 32'sd4087582, 32'sd1502976, 32'sd737547, -32'sd2227144, 32'sd2533746, 32'sd225519, 32'sd3271741, -32'sd689498, -32'sd228533, -32'sd2971505, 32'sd1139641, 32'sd4249097, 32'sd559089, 32'sd2732510, 32'sd296517, -32'sd1954562, 32'sd1510179, -32'sd1817207, 32'sd2331640, 32'sd4116063, -32'sd1453794, -32'sd4055490, -32'sd1907432, 32'sd1369730, -32'sd5031857, -32'sd122151, 32'sd1364809, 32'sd3507462, -32'sd3001439, -32'sd4117892, 32'sd797231, -32'sd1449500, -32'sd3758212, 32'sd354232, 32'sd1064763, -32'sd546932, 32'sd64710, -32'sd3805065, -32'sd4796, -32'sd894227, 32'sd1473799, -32'sd3436742, -32'sd351774, -32'sd1854049, 32'sd1920707, 32'sd1450847, 32'sd3642129, -32'sd767957, -32'sd3884070, 32'sd1788108, 32'sd3406393, 32'sd523607, 32'sd1048635, -32'sd709790, -32'sd291935, -32'sd1284343, 32'sd579413, 32'sd2220081, 32'sd314208, -32'sd194064, -32'sd2217019, -32'sd981819, 32'sd1642549, 32'sd1477043, -32'sd1427857, -32'sd2985096, -32'sd2842681, 32'sd1824139, 32'sd2792980, -32'sd3195285, -32'sd3427537, 32'sd1313053, 32'sd1540554, 32'sd2058842, 32'sd1764072, 32'sd222549, 32'sd2330932, 32'sd2241410, -32'sd1455205, -32'sd1778170, -32'sd292893, -32'sd2208422, -32'sd2748558, 32'sd450901},
        '{32'sd67071, -32'sd4002845, -32'sd666248, 32'sd3989555, 32'sd2515680, -32'sd229517, 32'sd618109, -32'sd2322424, 32'sd2675838, -32'sd1392160, 32'sd2800169, 32'sd136880, 32'sd4547544, -32'sd2748373, -32'sd441666, -32'sd2334828, -32'sd2813112, 32'sd3108053, 32'sd1170250, 32'sd1008796, 32'sd2657780, -32'sd1246789, -32'sd1681257, 32'sd1524991, -32'sd1065729, -32'sd1929484, -32'sd48662, 32'sd561959, -32'sd861594, 32'sd161342, -32'sd1906679, 32'sd3864447, -32'sd588213, 32'sd1912080, -32'sd2158396, 32'sd1958091, 32'sd2924359, 32'sd1676643, -32'sd1672293, 32'sd1505424, -32'sd2079830, 32'sd4854928, 32'sd1613263, 32'sd587531, -32'sd1384113, -32'sd651549, 32'sd5179523, -32'sd2898514, 32'sd166998, 32'sd587261, 32'sd4898019, -32'sd2163553, -32'sd2320295, 32'sd524708, 32'sd3839823, 32'sd439886, 32'sd2594340, -32'sd2570170, -32'sd3942154, 32'sd1308062, 32'sd3435025, -32'sd1462627, 32'sd1524957, 32'sd603115, -32'sd329237, 32'sd959383, 32'sd1489919, 32'sd1786869, -32'sd2916386, -32'sd3655410, -32'sd516903, 32'sd2685350, -32'sd1529107, 32'sd3611462, -32'sd2611420, -32'sd1439948, 32'sd1871213, 32'sd1600523, 32'sd1847706, 32'sd3036458, -32'sd1877932, -32'sd2046780, 32'sd588073, -32'sd495323, 32'sd1926267, -32'sd545573, -32'sd6090727, -32'sd574310, 32'sd353314, 32'sd2238542, 32'sd2330461, -32'sd463901, -32'sd1354223, 32'sd2285856, -32'sd1606040, -32'sd2178603, -32'sd1863217, -32'sd1234548, -32'sd3360836, -32'sd58248, -32'sd2241410, 32'sd342638, 32'sd1917469, 32'sd3232533, -32'sd2125099, 32'sd1490619, 32'sd3812098, 32'sd3526875, -32'sd1747872, -32'sd2757199, -32'sd553282, 32'sd2240961, 32'sd605900, 32'sd1899518, 32'sd1834602, -32'sd1799866, -32'sd2217539, 32'sd642219, 32'sd3186979, -32'sd654709, -32'sd1415870, -32'sd2749411, -32'sd489023, -32'sd1372671, 32'sd3353676, 32'sd2014641, -32'sd3079028, 32'sd4432370},
        '{32'sd2594797, -32'sd648562, -32'sd1823144, -32'sd1726344, -32'sd2350243, -32'sd1883529, -32'sd1412706, -32'sd1472821, 32'sd2367030, 32'sd2656245, -32'sd914541, -32'sd1149677, 32'sd1656694, 32'sd2372891, -32'sd3354971, -32'sd2298390, 32'sd2027386, -32'sd585518, 32'sd655532, 32'sd1531246, -32'sd2003834, -32'sd2005073, 32'sd2282460, -32'sd3157269, 32'sd3347418, 32'sd4401387, -32'sd1549766, 32'sd3440325, -32'sd1299448, 32'sd1404291, -32'sd1085018, -32'sd1352131, -32'sd939376, 32'sd1706682, 32'sd2124632, 32'sd1362644, 32'sd3349822, -32'sd278216, 32'sd380233, -32'sd2251945, 32'sd2692646, -32'sd1257841, 32'sd2732021, -32'sd59319, -32'sd2357291, 32'sd94221, 32'sd2829994, -32'sd1968569, 32'sd1071627, -32'sd3013303, 32'sd3784729, -32'sd1832887, -32'sd3450695, 32'sd2451113, -32'sd2740324, 32'sd4006544, 32'sd3105938, -32'sd175114, -32'sd2901945, -32'sd2527711, 32'sd1903451, -32'sd576593, 32'sd1696966, 32'sd4137133, -32'sd2564208, 32'sd368455, -32'sd322281, 32'sd4680119, -32'sd352591, -32'sd1989388, 32'sd3636706, 32'sd1850022, 32'sd6930, 32'sd1091666, 32'sd461439, 32'sd3522184, -32'sd824816, 32'sd4953981, -32'sd52639, 32'sd3323344, -32'sd4392504, -32'sd2744404, -32'sd419091, 32'sd755456, -32'sd764872, -32'sd2266811, -32'sd4935613, 32'sd4486919, 32'sd632805, -32'sd2715516, 32'sd2591882, -32'sd1090908, 32'sd2223976, 32'sd87453, -32'sd3258463, 32'sd2435721, -32'sd1591164, -32'sd2611899, -32'sd1149062, -32'sd384887, 32'sd1928998, 32'sd3457388, 32'sd316686, 32'sd2187517, 32'sd1537786, 32'sd3331942, 32'sd1342925, 32'sd1528397, -32'sd1312443, -32'sd909591, -32'sd1500781, -32'sd3527486, 32'sd331680, -32'sd42633, 32'sd3048375, -32'sd815765, -32'sd3725756, 32'sd402917, 32'sd203248, -32'sd3970410, 32'sd1834592, 32'sd1227337, 32'sd2689186, 32'sd1912394, 32'sd3856670, -32'sd3089827, -32'sd4150648, -32'sd780118},
        '{-32'sd1456131, -32'sd5399158, -32'sd3174859, 32'sd1107317, -32'sd2916194, -32'sd3408405, 32'sd2316778, -32'sd1482312, -32'sd1708057, 32'sd481909, 32'sd520726, -32'sd3100617, 32'sd2852338, -32'sd2263245, 32'sd1369747, 32'sd726108, 32'sd68867, -32'sd3178931, 32'sd2713873, -32'sd2246997, -32'sd2193896, -32'sd1077506, 32'sd2388293, 32'sd688257, -32'sd2712520, 32'sd277283, 32'sd2732136, -32'sd635338, -32'sd2362369, 32'sd194303, 32'sd1464414, -32'sd1348925, -32'sd38520, 32'sd4040875, -32'sd1143971, 32'sd497659, 32'sd1622793, 32'sd2810664, 32'sd2943412, 32'sd1010770, -32'sd3898079, 32'sd2915956, -32'sd2229014, -32'sd2836999, -32'sd1651067, 32'sd3105468, 32'sd618651, -32'sd3568787, -32'sd4892308, 32'sd81, 32'sd1538414, 32'sd3331576, -32'sd1442842, 32'sd2269009, 32'sd902131, 32'sd2059815, 32'sd971307, -32'sd1362625, -32'sd1754702, 32'sd2074158, 32'sd708205, -32'sd281225, -32'sd1287282, -32'sd293204, 32'sd1436755, 32'sd2844688, 32'sd1417272, -32'sd191696, -32'sd3593999, 32'sd2117267, -32'sd2084321, 32'sd1430183, 32'sd2425506, 32'sd3348286, -32'sd2505565, -32'sd4620402, 32'sd1301059, 32'sd367654, 32'sd571250, 32'sd2818466, -32'sd1546131, -32'sd3977201, -32'sd2552129, 32'sd2014686, -32'sd1052140, -32'sd849994, 32'sd3492617, 32'sd144947, -32'sd571213, -32'sd731393, 32'sd3498781, 32'sd3425221, 32'sd1262118, -32'sd462784, -32'sd1702441, 32'sd2158510, -32'sd3202529, -32'sd2087210, -32'sd558746, -32'sd1706870, -32'sd2145360, -32'sd111800, 32'sd3291014, -32'sd2450358, 32'sd1228673, -32'sd6412929, 32'sd1608074, 32'sd2365636, -32'sd289326, -32'sd39527, 32'sd264123, 32'sd2143584, 32'sd478529, 32'sd657142, -32'sd1060147, -32'sd1677434, 32'sd2955071, -32'sd1057870, -32'sd314393, -32'sd206925, 32'sd3753462, -32'sd1076869, 32'sd494230, 32'sd2077355, 32'sd897698, 32'sd2165368, -32'sd1922394, 32'sd2365532},
        '{-32'sd279114, -32'sd777376, 32'sd365915, -32'sd1400593, -32'sd2228617, 32'sd1571423, -32'sd1154290, 32'sd3471490, 32'sd904870, -32'sd2191290, 32'sd784262, 32'sd286788, 32'sd1383992, -32'sd2494520, -32'sd4097368, 32'sd239288, -32'sd2381509, 32'sd2459976, 32'sd326773, -32'sd3146028, 32'sd16115, -32'sd374613, -32'sd1860547, -32'sd2735523, 32'sd3375498, 32'sd2181175, -32'sd1157981, 32'sd2367941, -32'sd1774194, -32'sd76095, -32'sd3618122, 32'sd3711722, 32'sd465316, -32'sd852974, 32'sd322431, 32'sd752699, -32'sd995821, 32'sd2416567, 32'sd2194062, -32'sd2512130, 32'sd2358426, 32'sd376111, -32'sd2393948, -32'sd3640479, 32'sd1171537, -32'sd3284949, -32'sd2804877, 32'sd1824499, 32'sd1403579, -32'sd345655, -32'sd2113374, 32'sd2698041, -32'sd2254944, 32'sd2092543, 32'sd384308, 32'sd600786, -32'sd3695881, -32'sd3639501, -32'sd271332, -32'sd1964112, -32'sd239767, 32'sd3401019, -32'sd2040433, -32'sd868567, 32'sd109263, 32'sd2747951, 32'sd3747334, 32'sd490564, -32'sd1115806, 32'sd1520178, -32'sd748295, -32'sd592995, -32'sd20540, 32'sd2250912, -32'sd1331544, 32'sd511419, 32'sd2162195, -32'sd203264, -32'sd138268, -32'sd2173978, 32'sd2078591, 32'sd2608507, 32'sd62481, -32'sd567447, -32'sd4537336, 32'sd3197714, -32'sd2530879, 32'sd3529826, 32'sd1277224, 32'sd345003, 32'sd1286256, 32'sd1423426, -32'sd1229924, 32'sd3906903, 32'sd703658, 32'sd342082, -32'sd359069, 32'sd856960, -32'sd3134785, 32'sd2073053, 32'sd1951688, 32'sd2218952, 32'sd412296, -32'sd9047, -32'sd3368805, -32'sd600343, 32'sd1225457, 32'sd1504664, 32'sd1807801, 32'sd691922, -32'sd4789445, 32'sd1226986, -32'sd909785, 32'sd120771, 32'sd2473511, 32'sd181071, -32'sd1503814, -32'sd2095821, -32'sd293653, -32'sd2009490, -32'sd1979493, 32'sd1516811, 32'sd3033322, 32'sd3200168, -32'sd1248993, 32'sd3613244, -32'sd1274455, 32'sd35481},
        '{-32'sd3703127, 32'sd513887, 32'sd670421, 32'sd418385, -32'sd2429005, 32'sd1295134, 32'sd3591659, 32'sd2096589, 32'sd2080421, -32'sd100042, 32'sd2170024, -32'sd1248721, 32'sd728115, 32'sd986369, 32'sd385677, 32'sd3144007, 32'sd608566, -32'sd4078717, 32'sd248078, 32'sd381998, -32'sd286948, -32'sd3230477, -32'sd4647302, 32'sd2484602, -32'sd472368, -32'sd70044, -32'sd2308886, -32'sd85044, -32'sd259732, 32'sd2544602, 32'sd3256874, -32'sd1007282, -32'sd1335947, 32'sd1490057, -32'sd1108268, -32'sd821783, 32'sd975646, -32'sd1903412, 32'sd3255491, 32'sd2220704, 32'sd1311648, -32'sd3147953, 32'sd3795993, 32'sd744586, 32'sd1317451, 32'sd2488524, 32'sd4276318, 32'sd670028, 32'sd3339150, 32'sd743326, 32'sd435235, -32'sd2965135, 32'sd399226, -32'sd4166860, 32'sd441814, -32'sd465777, -32'sd2200260, -32'sd3376611, -32'sd1293509, -32'sd1873835, 32'sd2462652, -32'sd1527018, -32'sd2747974, 32'sd1870154, 32'sd440352, -32'sd155368, 32'sd1030243, 32'sd1582583, 32'sd679387, 32'sd2884091, -32'sd3989293, -32'sd1127648, 32'sd3147809, 32'sd1505677, -32'sd2788294, 32'sd3016242, 32'sd2333644, 32'sd2841218, 32'sd3026572, -32'sd4434452, -32'sd506821, 32'sd1137153, 32'sd1238843, -32'sd550867, 32'sd2754387, -32'sd989775, -32'sd146173, -32'sd3942349, 32'sd2893811, 32'sd3651226, 32'sd2112855, 32'sd3852046, 32'sd1459162, -32'sd2486320, 32'sd3072630, -32'sd4652627, -32'sd2269205, -32'sd275565, -32'sd2149465, 32'sd1970615, -32'sd1774885, -32'sd2151517, 32'sd978368, -32'sd2764571, 32'sd850983, -32'sd2382470, 32'sd1042417, -32'sd1128480, 32'sd2359218, -32'sd2088008, -32'sd1145551, 32'sd1875292, -32'sd3195072, 32'sd438510, -32'sd328267, 32'sd4405480, -32'sd1577923, 32'sd2650636, -32'sd3995802, 32'sd4303052, -32'sd3364268, -32'sd1416036, 32'sd2550655, -32'sd1520041, -32'sd1951523, -32'sd5371883, 32'sd3075946, 32'sd3752621},
        '{-32'sd2631911, 32'sd2880116, -32'sd4733292, 32'sd2831281, 32'sd2004, -32'sd2487103, -32'sd2228390, 32'sd1647812, -32'sd1155545, -32'sd3697416, -32'sd754046, 32'sd769083, 32'sd1255348, -32'sd1434378, -32'sd880295, -32'sd93782, 32'sd2156940, 32'sd551501, -32'sd2683237, -32'sd1540492, -32'sd1136631, -32'sd500237, -32'sd4895253, -32'sd754852, -32'sd1548142, 32'sd2781504, 32'sd2998410, -32'sd2386755, -32'sd2738501, 32'sd4542363, -32'sd672132, -32'sd2430652, -32'sd1710972, 32'sd511916, 32'sd270833, -32'sd1418101, 32'sd804808, 32'sd2133064, -32'sd3024678, 32'sd1923052, -32'sd1610573, 32'sd2382503, 32'sd1829544, -32'sd2955255, -32'sd2545002, 32'sd2121635, 32'sd3621921, 32'sd3342060, 32'sd363343, 32'sd1225543, 32'sd4167633, -32'sd608459, -32'sd366704, -32'sd1232336, -32'sd2031689, -32'sd2203418, -32'sd1830267, -32'sd2104, 32'sd1057417, 32'sd1079663, 32'sd2363762, -32'sd1464246, 32'sd4319528, 32'sd806578, -32'sd3812555, -32'sd1652103, 32'sd4420387, 32'sd2844803, 32'sd325263, 32'sd626192, -32'sd2683865, -32'sd5360954, -32'sd2215656, -32'sd2906635, 32'sd2105794, 32'sd4487197, 32'sd3960241, -32'sd1654889, -32'sd2030020, -32'sd278856, 32'sd4526679, 32'sd592812, 32'sd787269, 32'sd737100, 32'sd565275, -32'sd1450572, -32'sd722569, 32'sd2013321, -32'sd2168321, -32'sd3884194, -32'sd1026780, 32'sd414839, -32'sd868000, -32'sd2701438, -32'sd4257407, -32'sd1888530, 32'sd1468981, 32'sd3283472, -32'sd982027, 32'sd1360913, -32'sd1773495, 32'sd2880770, 32'sd1136061, -32'sd1815700, -32'sd4755934, 32'sd84759, -32'sd386560, 32'sd507963, -32'sd2741047, 32'sd2353880, 32'sd884835, 32'sd2868537, 32'sd4383258, -32'sd109043, -32'sd209756, 32'sd438490, 32'sd1290234, -32'sd2208160, 32'sd2960496, 32'sd1706033, -32'sd1474992, -32'sd1317124, -32'sd2816815, -32'sd2770725, -32'sd3831977, 32'sd845122, 32'sd1987308, -32'sd1778966},
        '{-32'sd3432586, 32'sd618544, -32'sd668290, 32'sd223308, 32'sd3464124, 32'sd3115763, -32'sd3417622, 32'sd2918566, -32'sd1409157, 32'sd24515, 32'sd293872, 32'sd400476, 32'sd606334, -32'sd528052, -32'sd1356509, 32'sd2395779, 32'sd2643995, -32'sd1870258, -32'sd3118235, 32'sd402523, 32'sd1378548, 32'sd366728, 32'sd1587179, 32'sd2795910, 32'sd2579906, 32'sd2687953, 32'sd2690206, -32'sd1098175, 32'sd1181131, -32'sd3349980, -32'sd4537312, -32'sd1883542, -32'sd11590, -32'sd3318727, -32'sd21994, 32'sd2198858, 32'sd32553, -32'sd1339214, -32'sd87999, 32'sd3171257, -32'sd982353, 32'sd1250571, -32'sd1434170, -32'sd3168068, -32'sd1861644, 32'sd208325, 32'sd3311380, 32'sd1427364, -32'sd2796358, 32'sd890016, 32'sd897745, 32'sd3222975, -32'sd4413655, 32'sd2917795, -32'sd4341441, -32'sd1172000, -32'sd2089233, -32'sd804281, -32'sd690305, -32'sd1192461, 32'sd4043300, 32'sd769577, 32'sd603984, 32'sd3341234, 32'sd1482476, 32'sd3988371, -32'sd2195459, -32'sd526892, 32'sd333659, -32'sd4020891, 32'sd3756998, 32'sd217708, -32'sd1802699, 32'sd2588393, -32'sd5579955, -32'sd2671566, -32'sd2153564, 32'sd181661, 32'sd2931098, -32'sd564307, -32'sd2523476, 32'sd602748, 32'sd2950152, -32'sd397017, -32'sd51200, -32'sd4810823, 32'sd42665, -32'sd512514, 32'sd1323107, -32'sd988004, -32'sd2145640, -32'sd2854942, 32'sd490887, -32'sd671953, 32'sd1272744, 32'sd1141243, -32'sd4065384, -32'sd1071730, 32'sd2294018, -32'sd479268, -32'sd1441835, -32'sd1989181, 32'sd3712926, -32'sd3007009, -32'sd774799, -32'sd3214882, 32'sd3017044, -32'sd379873, 32'sd530401, -32'sd1948101, 32'sd273162, 32'sd115993, -32'sd2152872, -32'sd1635125, 32'sd1770354, 32'sd3646577, -32'sd2406408, -32'sd1911909, 32'sd2292012, -32'sd1716061, 32'sd1989248, -32'sd2414535, 32'sd1635121, -32'sd2826880, 32'sd1771029, 32'sd1517803, -32'sd1039505, -32'sd216377},
        '{32'sd391831, -32'sd2776229, -32'sd4087902, 32'sd3835332, 32'sd2363710, 32'sd2752218, -32'sd1287369, 32'sd2161528, -32'sd1088905, 32'sd1310257, 32'sd2390794, 32'sd3394942, 32'sd1088437, -32'sd350159, -32'sd894377, -32'sd3323145, -32'sd1357357, -32'sd1879486, -32'sd460707, -32'sd1960094, -32'sd1793794, 32'sd2131651, -32'sd4077355, -32'sd392253, -32'sd670233, 32'sd3186343, -32'sd4582262, 32'sd403378, 32'sd1584249, 32'sd2127140, -32'sd420781, 32'sd134419, -32'sd3518835, -32'sd252001, 32'sd1914649, 32'sd40027, 32'sd1022440, 32'sd1201448, -32'sd4859155, -32'sd1970750, 32'sd4811674, 32'sd1505966, 32'sd1756882, 32'sd2705805, 32'sd2968378, -32'sd2549215, -32'sd599570, -32'sd465589, 32'sd86045, -32'sd2650643, 32'sd3550203, 32'sd904198, 32'sd1673731, 32'sd2785214, 32'sd3710308, 32'sd697452, -32'sd2242246, 32'sd2353637, -32'sd1155570, 32'sd989372, 32'sd2706590, 32'sd1366408, -32'sd57535, 32'sd2293344, 32'sd454916, -32'sd3905411, 32'sd840445, 32'sd1700882, -32'sd3748896, 32'sd1544196, 32'sd359475, 32'sd3418887, 32'sd1168610, -32'sd1753996, 32'sd3452959, 32'sd3395531, 32'sd323908, -32'sd1601973, 32'sd2996336, 32'sd1911057, -32'sd1370441, -32'sd2450149, 32'sd1134768, -32'sd774748, 32'sd3172463, -32'sd3100776, 32'sd850692, -32'sd815498, 32'sd1845096, -32'sd899364, 32'sd473206, 32'sd2626846, 32'sd249610, 32'sd2874870, 32'sd141329, -32'sd2210328, 32'sd664402, 32'sd3744201, -32'sd2276722, 32'sd1511135, 32'sd112154, -32'sd1052116, -32'sd2988972, 32'sd1211680, -32'sd1235957, -32'sd1703031, 32'sd538186, 32'sd1494264, -32'sd2329213, 32'sd2405972, -32'sd3890632, 32'sd464004, 32'sd1364526, 32'sd61483, 32'sd1357853, 32'sd1130830, -32'sd2643661, 32'sd279367, 32'sd2903729, -32'sd4777912, 32'sd4013479, 32'sd885130, -32'sd13934, -32'sd1037633, 32'sd3329756, 32'sd1901106, -32'sd912914, 32'sd3897204},
        '{32'sd3348377, 32'sd3163746, 32'sd306902, -32'sd1783629, -32'sd3919111, -32'sd475206, 32'sd1502575, 32'sd2924255, -32'sd3282933, 32'sd1596800, -32'sd2276960, 32'sd533845, -32'sd659443, 32'sd1577697, -32'sd2200367, -32'sd3558620, 32'sd3732567, -32'sd2408322, 32'sd1191945, 32'sd737849, -32'sd1258722, -32'sd843531, 32'sd2668968, 32'sd1472858, 32'sd1742875, 32'sd3505245, -32'sd1595383, -32'sd40730, -32'sd563510, 32'sd2121214, -32'sd2266015, -32'sd2940451, 32'sd1186053, -32'sd1565960, 32'sd532681, -32'sd1340397, 32'sd3434501, -32'sd1368616, 32'sd869641, 32'sd1326753, 32'sd2351324, 32'sd1562389, 32'sd999114, 32'sd2812175, -32'sd3849238, -32'sd122570, -32'sd478229, -32'sd215937, -32'sd724606, -32'sd1748145, 32'sd2652593, 32'sd1276014, 32'sd129947, 32'sd1027865, -32'sd2806023, -32'sd2334249, 32'sd3620935, 32'sd123659, -32'sd3474709, 32'sd2001822, 32'sd2375154, 32'sd92082, 32'sd1469922, 32'sd2056982, 32'sd1052860, -32'sd2285259, -32'sd375089, -32'sd1522825, 32'sd2660000, -32'sd675577, 32'sd3157767, 32'sd314753, 32'sd1083674, 32'sd3421586, -32'sd4180510, 32'sd2888284, -32'sd2272001, -32'sd708748, 32'sd1519275, 32'sd1101217, 32'sd406607, 32'sd1238099, 32'sd3330183, 32'sd1665131, -32'sd1310981, 32'sd3577664, 32'sd693936, 32'sd3160800, 32'sd4332371, -32'sd2880920, -32'sd2984213, -32'sd788392, -32'sd1141463, 32'sd798061, -32'sd2093092, -32'sd2689664, -32'sd994126, -32'sd3084339, 32'sd3979100, 32'sd356190, 32'sd2675887, 32'sd2609196, -32'sd1725792, -32'sd857328, -32'sd615325, 32'sd2400984, 32'sd3308862, -32'sd1614900, -32'sd2905450, 32'sd3288259, 32'sd2616285, -32'sd2726664, 32'sd706642, 32'sd4521351, 32'sd207215, 32'sd1237866, 32'sd923092, 32'sd757627, 32'sd355492, 32'sd3811365, -32'sd837261, -32'sd4188773, -32'sd1435300, 32'sd598817, 32'sd1737847, 32'sd1814605, -32'sd852683, -32'sd2008594},
        '{32'sd753163, 32'sd1060514, 32'sd617649, 32'sd2541689, 32'sd691094, -32'sd2650924, 32'sd2362528, -32'sd3710976, 32'sd1922833, -32'sd266247, -32'sd2979375, -32'sd1322513, -32'sd2878244, -32'sd3920371, 32'sd4032242, 32'sd120847, 32'sd1703927, 32'sd847754, -32'sd1415319, 32'sd608575, 32'sd1817775, -32'sd2985999, 32'sd677378, 32'sd2268450, 32'sd1385893, -32'sd128967, -32'sd2461704, -32'sd1717037, 32'sd712140, 32'sd3192837, -32'sd1983034, -32'sd4249334, 32'sd2860285, 32'sd2760420, 32'sd2659887, 32'sd313841, 32'sd1311827, -32'sd576563, -32'sd1054507, -32'sd2442574, -32'sd3086913, -32'sd1407444, 32'sd570127, 32'sd2378298, -32'sd650738, -32'sd2081109, 32'sd3011485, -32'sd3139637, 32'sd2049965, 32'sd2431381, -32'sd1698723, -32'sd2291243, 32'sd1586983, 32'sd1835603, -32'sd3870443, -32'sd2619128, 32'sd2900304, -32'sd2595228, 32'sd1003501, -32'sd3142644, 32'sd4592014, 32'sd349631, -32'sd4079532, 32'sd1606258, -32'sd697158, -32'sd729980, 32'sd851131, 32'sd1354980, 32'sd2411152, 32'sd390599, -32'sd2558091, 32'sd321317, 32'sd1744771, 32'sd3039563, -32'sd4623104, -32'sd1314618, 32'sd1775846, -32'sd668911, 32'sd2119904, 32'sd2774353, 32'sd1255385, -32'sd1768078, 32'sd1701303, -32'sd2018146, 32'sd1446146, 32'sd1705405, 32'sd10252, -32'sd1514694, 32'sd2816067, 32'sd4955689, 32'sd2149251, 32'sd3528299, 32'sd3226763, -32'sd1175321, 32'sd3160254, -32'sd3409086, -32'sd901082, -32'sd4329223, -32'sd984623, -32'sd547917, 32'sd680083, -32'sd1783601, 32'sd2827555, -32'sd46578, 32'sd2786483, 32'sd263934, 32'sd2694206, -32'sd2617235, 32'sd780246, -32'sd1543302, 32'sd2012593, -32'sd2930324, -32'sd5479865, 32'sd587270, 32'sd3125223, 32'sd998423, -32'sd3591449, 32'sd975771, -32'sd1948949, 32'sd1096488, -32'sd1661859, 32'sd883536, 32'sd2271987, 32'sd212037, -32'sd1520686, -32'sd5458401, 32'sd4877214, 32'sd4032536},
        '{32'sd1333463, 32'sd595433, -32'sd1090471, 32'sd1384502, 32'sd2470612, -32'sd336395, 32'sd1718644, 32'sd793733, 32'sd405918, -32'sd1808908, 32'sd1847534, 32'sd3240073, -32'sd1135983, 32'sd2779267, 32'sd1487160, -32'sd3495707, -32'sd3461433, -32'sd269650, 32'sd1157454, -32'sd3082354, -32'sd87603, -32'sd539115, 32'sd3057913, -32'sd1104875, 32'sd2771339, 32'sd2882353, -32'sd289800, -32'sd335544, 32'sd358709, 32'sd1581526, -32'sd1359464, -32'sd2774755, 32'sd1228797, -32'sd285040, 32'sd122831, 32'sd107447, -32'sd152840, 32'sd1151454, 32'sd2226143, 32'sd2646739, 32'sd336897, 32'sd2152333, 32'sd1429601, 32'sd3777039, 32'sd4959029, -32'sd2970879, -32'sd2246809, 32'sd2132666, 32'sd3691619, -32'sd2852198, -32'sd3283652, 32'sd5010947, -32'sd2783807, -32'sd3636411, 32'sd593960, -32'sd35041, -32'sd1527127, 32'sd1622669, 32'sd1139157, 32'sd1942404, -32'sd3733992, -32'sd3904648, -32'sd2680187, 32'sd1520439, -32'sd743189, -32'sd550267, -32'sd430283, -32'sd883282, 32'sd3771569, 32'sd444289, -32'sd2508992, 32'sd446548, -32'sd1267604, -32'sd3478528, -32'sd4058729, 32'sd436629, -32'sd2549293, -32'sd1400046, -32'sd136004, -32'sd2040061, -32'sd563779, 32'sd592979, -32'sd1106799, 32'sd3086341, 32'sd2173644, -32'sd3537536, -32'sd2049322, 32'sd2732418, -32'sd3782423, 32'sd4214904, -32'sd4159404, -32'sd1612111, 32'sd423303, 32'sd3296779, 32'sd1031820, 32'sd1737230, 32'sd1811421, -32'sd1783523, 32'sd2582022, 32'sd4158252, 32'sd3420263, -32'sd652348, -32'sd1786406, -32'sd1597738, 32'sd2529716, -32'sd2190647, -32'sd1264497, -32'sd2530319, 32'sd2647882, -32'sd106525, -32'sd2179934, -32'sd3810017, 32'sd3326552, -32'sd4440177, 32'sd3142187, -32'sd1959172, 32'sd3633889, 32'sd2687404, -32'sd716938, 32'sd3503291, 32'sd2278281, -32'sd2230365, -32'sd4344156, -32'sd4414600, 32'sd174384, -32'sd1525914, 32'sd4744910, 32'sd827991},
        '{32'sd2015772, 32'sd827597, -32'sd2530438, -32'sd1203621, 32'sd3438291, -32'sd1119394, -32'sd2570621, 32'sd2149605, 32'sd1904158, -32'sd2620254, 32'sd20968, 32'sd2783904, 32'sd1423201, 32'sd1541066, -32'sd45919, 32'sd1805494, 32'sd1826606, -32'sd1227732, -32'sd3990604, 32'sd1205429, -32'sd459848, 32'sd896227, 32'sd4052997, 32'sd3228656, 32'sd1677803, 32'sd1453830, -32'sd4314599, 32'sd1519775, -32'sd500102, -32'sd151961, -32'sd3024007, 32'sd838747, -32'sd4809869, -32'sd1979986, -32'sd300830, 32'sd2879379, -32'sd2528006, -32'sd2319627, -32'sd1000440, 32'sd3852353, -32'sd2032714, 32'sd3517871, 32'sd2384897, 32'sd4107739, 32'sd3940454, 32'sd2164533, -32'sd3242377, 32'sd2285248, 32'sd1450784, -32'sd2447065, -32'sd411235, -32'sd931391, 32'sd1672843, 32'sd1041484, 32'sd1902480, 32'sd162196, -32'sd2810695, 32'sd323713, 32'sd1201025, 32'sd1508292, -32'sd3555467, -32'sd1775384, 32'sd2349349, 32'sd91038, 32'sd3848932, 32'sd1438957, 32'sd2725307, -32'sd2931515, 32'sd2086835, -32'sd3292309, 32'sd1147723, -32'sd3002283, 32'sd102060, -32'sd1278928, 32'sd273152, 32'sd2894257, -32'sd282878, 32'sd428790, 32'sd3020127, -32'sd1180334, -32'sd2099204, -32'sd2191475, 32'sd1558012, 32'sd1035492, -32'sd1116293, -32'sd931484, -32'sd3755063, -32'sd388487, -32'sd1264153, 32'sd1105874, -32'sd3223839, -32'sd3076917, -32'sd42122, 32'sd367319, -32'sd1621617, -32'sd1958836, 32'sd1735140, -32'sd2662112, -32'sd969332, 32'sd696178, 32'sd1492238, -32'sd1445603, -32'sd9796, 32'sd188447, -32'sd1706652, -32'sd1000685, -32'sd3040937, 32'sd1300198, -32'sd2979087, 32'sd2545267, -32'sd5376987, -32'sd3818129, -32'sd1714740, -32'sd1003763, 32'sd252782, -32'sd1277377, -32'sd1064362, -32'sd3470827, -32'sd702412, -32'sd1243631, 32'sd1296247, 32'sd3232707, 32'sd2693766, -32'sd2736125, 32'sd280468, -32'sd1376926, -32'sd3010180, -32'sd1128257},
        '{32'sd632068, 32'sd2314140, -32'sd2172393, 32'sd3188451, 32'sd1529367, -32'sd2277099, 32'sd2828787, 32'sd2049270, -32'sd1107991, 32'sd1292393, -32'sd134976, -32'sd1150803, 32'sd1041142, -32'sd1777548, -32'sd711106, 32'sd2536620, 32'sd2092659, 32'sd1178944, 32'sd2334183, 32'sd527960, 32'sd434978, -32'sd2237219, 32'sd865294, 32'sd263346, 32'sd98545, 32'sd1453007, 32'sd4425262, -32'sd395798, 32'sd1213950, -32'sd4214486, -32'sd496235, -32'sd483490, 32'sd1421895, -32'sd2000001, 32'sd2204990, 32'sd1285308, -32'sd1845600, 32'sd380766, 32'sd1663296, -32'sd2021403, 32'sd2432130, -32'sd2687473, -32'sd2400371, 32'sd1908145, -32'sd2225184, -32'sd1035357, -32'sd42602, -32'sd2892894, -32'sd3342717, 32'sd1676651, -32'sd208892, 32'sd2427430, 32'sd378384, 32'sd2967952, -32'sd3161990, -32'sd159829, 32'sd1171845, 32'sd1136179, 32'sd1893391, 32'sd297802, 32'sd840327, -32'sd1890513, -32'sd862791, -32'sd1091072, -32'sd2416231, -32'sd1743763, 32'sd596262, 32'sd2174103, -32'sd2323916, 32'sd3875236, 32'sd42034, 32'sd2119047, 32'sd1833394, 32'sd1940841, 32'sd2016458, 32'sd1784227, -32'sd433722, 32'sd4525643, -32'sd2745152, -32'sd1548031, 32'sd39984, 32'sd3244562, -32'sd681830, 32'sd2959018, 32'sd602540, -32'sd2349435, 32'sd4211789, -32'sd1063750, -32'sd1395479, -32'sd3340311, -32'sd411500, -32'sd144597, 32'sd2833625, -32'sd5792030, 32'sd3772109, -32'sd2200365, 32'sd449182, -32'sd1043862, -32'sd611734, -32'sd3442786, 32'sd2546808, -32'sd557858, 32'sd3641586, -32'sd743288, -32'sd1956769, 32'sd997049, -32'sd362042, -32'sd4992999, -32'sd1005560, 32'sd312934, 32'sd2536339, 32'sd2117900, 32'sd1761629, -32'sd1244533, 32'sd3168356, 32'sd1475200, 32'sd506572, -32'sd83812, 32'sd71809, -32'sd115370, 32'sd2106867, 32'sd3843741, -32'sd1092515, 32'sd1302377, -32'sd2778292, 32'sd3461137, -32'sd2026458, 32'sd455675},
        '{-32'sd1031593, 32'sd3461084, 32'sd1992823, -32'sd277042, 32'sd917736, -32'sd2560555, -32'sd2767859, -32'sd613385, 32'sd1466804, -32'sd989492, -32'sd1998758, -32'sd2048192, -32'sd2086171, 32'sd167732, 32'sd3422369, -32'sd669963, -32'sd2940131, 32'sd2118697, 32'sd4541858, 32'sd1723650, -32'sd333337, -32'sd3998961, 32'sd259072, 32'sd1465931, -32'sd3096664, -32'sd2187267, 32'sd330715, 32'sd1047197, -32'sd1412867, -32'sd3434625, -32'sd3851, -32'sd692721, 32'sd2742862, -32'sd1130274, -32'sd350732, 32'sd193875, 32'sd1685844, -32'sd1220241, 32'sd1796580, 32'sd1216325, -32'sd4920686, -32'sd428436, 32'sd3189761, 32'sd1418151, 32'sd2693329, 32'sd1632079, -32'sd1401371, -32'sd1871823, 32'sd2864037, 32'sd3022907, -32'sd2508427, 32'sd80614, -32'sd2026149, -32'sd253888, -32'sd76805, -32'sd3070506, -32'sd1884478, -32'sd4386444, 32'sd2278224, 32'sd2170343, 32'sd3321205, 32'sd4446209, 32'sd2267217, 32'sd2370415, 32'sd306937, 32'sd1988007, -32'sd1144690, 32'sd107536, 32'sd2205342, -32'sd105505, 32'sd760476, 32'sd2377065, -32'sd2750074, -32'sd1565965, 32'sd586797, 32'sd3336371, 32'sd1055602, -32'sd276914, 32'sd2677530, -32'sd2895350, -32'sd2976704, -32'sd1132706, 32'sd465873, -32'sd1233584, 32'sd2639404, 32'sd1014254, 32'sd2546917, -32'sd2915258, 32'sd418816, 32'sd3119434, 32'sd1191684, -32'sd774737, 32'sd2569603, 32'sd1023439, -32'sd3215127, 32'sd2406337, -32'sd2997110, -32'sd2784557, -32'sd1719509, 32'sd598249, 32'sd2082976, -32'sd35437, 32'sd644043, 32'sd493352, 32'sd2650513, 32'sd580868, -32'sd889242, 32'sd2790254, 32'sd1558447, -32'sd2250269, 32'sd2388474, 32'sd1463985, -32'sd3862567, 32'sd808402, 32'sd1446196, 32'sd719710, -32'sd2301020, 32'sd4957927, -32'sd3047139, 32'sd3157799, -32'sd1953096, -32'sd601819, 32'sd2654995, 32'sd2276780, 32'sd866973, -32'sd3153395, 32'sd2091818, 32'sd1816978},
        '{-32'sd635163, -32'sd295472, -32'sd1729628, 32'sd1524348, -32'sd3332413, 32'sd150767, 32'sd1416306, 32'sd345267, -32'sd1251876, 32'sd3408803, 32'sd1216769, 32'sd2050003, 32'sd2304089, -32'sd1675636, -32'sd376923, 32'sd981070, 32'sd2433271, 32'sd3143694, 32'sd1530102, -32'sd1331608, -32'sd5319831, 32'sd102222, -32'sd2127542, 32'sd1643325, 32'sd1245107, 32'sd264700, 32'sd216256, -32'sd1036191, -32'sd2238581, 32'sd1636756, 32'sd2955152, 32'sd3153778, -32'sd518594, 32'sd2733718, 32'sd1726873, 32'sd2325289, -32'sd2347880, -32'sd4706004, 32'sd2925738, -32'sd1062355, 32'sd1219154, -32'sd4027383, 32'sd272805, -32'sd927804, 32'sd2629389, -32'sd3929109, -32'sd308803, 32'sd935601, -32'sd4469067, 32'sd188820, 32'sd1135056, -32'sd788995, 32'sd3092812, -32'sd2828952, -32'sd3603393, -32'sd588495, -32'sd3687671, -32'sd45133, 32'sd1371200, 32'sd4786531, 32'sd1632254, 32'sd2395552, 32'sd1184092, -32'sd4304922, -32'sd5030205, -32'sd3032692, 32'sd1704147, 32'sd721806, -32'sd592767, -32'sd2530320, 32'sd1965136, -32'sd4060300, -32'sd1634205, -32'sd2925204, 32'sd1417931, -32'sd3244357, -32'sd520961, -32'sd1355418, -32'sd5135015, 32'sd360582, -32'sd2672644, 32'sd1614682, 32'sd5042955, -32'sd1279042, 32'sd1620997, 32'sd1171667, 32'sd3006070, -32'sd1994933, 32'sd1987246, -32'sd2857985, 32'sd1347157, -32'sd1484325, 32'sd1378915, -32'sd2776249, -32'sd2827766, -32'sd1529921, 32'sd3189878, 32'sd3251339, -32'sd3213409, -32'sd1643025, -32'sd387924, -32'sd3002570, 32'sd793879, 32'sd698391, 32'sd1849521, 32'sd3520289, 32'sd4681362, 32'sd550338, -32'sd3440225, 32'sd1888400, 32'sd2004574, 32'sd850649, 32'sd3336700, 32'sd383924, -32'sd417344, 32'sd2098876, -32'sd1617349, 32'sd2225577, -32'sd1916065, 32'sd1122229, -32'sd487050, 32'sd1344182, -32'sd183343, 32'sd2126630, 32'sd628902, -32'sd1397444, -32'sd2494636, -32'sd754463},
        '{32'sd709624, -32'sd1726232, -32'sd2065602, 32'sd1206211, -32'sd2712316, -32'sd1044100, -32'sd2106866, 32'sd3102643, 32'sd884975, 32'sd2290590, 32'sd544859, -32'sd1533447, 32'sd4069696, 32'sd2529266, -32'sd1635720, 32'sd1288452, -32'sd3483150, -32'sd2016080, -32'sd4470058, 32'sd751778, -32'sd2139672, 32'sd2019870, -32'sd2535504, -32'sd341124, -32'sd3041633, -32'sd1018347, 32'sd1243614, 32'sd2523643, -32'sd3529241, -32'sd2158039, -32'sd2003072, -32'sd2793282, 32'sd2516595, -32'sd345946, 32'sd2342501, -32'sd3815008, 32'sd113917, -32'sd452231, 32'sd1013027, -32'sd2005576, 32'sd2799008, -32'sd1536401, 32'sd3306963, 32'sd2628868, -32'sd633868, 32'sd1524392, 32'sd2016658, 32'sd221213, 32'sd344036, -32'sd1418223, 32'sd3568884, 32'sd944426, -32'sd1143658, -32'sd1547152, 32'sd872257, 32'sd297619, 32'sd1693360, 32'sd2260302, -32'sd1459873, 32'sd2178485, -32'sd1424270, 32'sd1821302, -32'sd1513862, 32'sd1517349, -32'sd137206, 32'sd60890, 32'sd1937960, -32'sd546146, -32'sd144578, -32'sd2842565, -32'sd594905, 32'sd67918, -32'sd66029, 32'sd868661, -32'sd2401190, -32'sd3034299, -32'sd1122793, 32'sd4233717, -32'sd940021, 32'sd3625513, -32'sd261718, -32'sd4246999, -32'sd2605652, 32'sd15535, 32'sd2518725, -32'sd2436699, -32'sd3812474, 32'sd131145, -32'sd1757529, 32'sd1537447, 32'sd2730727, 32'sd366997, -32'sd750780, 32'sd726842, -32'sd963892, 32'sd3438877, -32'sd2488436, 32'sd983338, 32'sd2907302, -32'sd880738, 32'sd3023887, -32'sd456163, -32'sd1796033, 32'sd105234, 32'sd2380062, -32'sd3732175, -32'sd747511, -32'sd918036, 32'sd3230826, 32'sd2318081, 32'sd784138, 32'sd3255215, 32'sd2328124, -32'sd823170, 32'sd2558788, 32'sd626551, -32'sd1480046, 32'sd2844616, -32'sd2142593, -32'sd2329411, 32'sd3468025, 32'sd859215, -32'sd1070660, -32'sd1313803, 32'sd3935414, 32'sd2467362, 32'sd4101903, -32'sd1371750},
        '{32'sd3435478, -32'sd3595763, -32'sd2059916, -32'sd356375, 32'sd1106733, -32'sd393641, 32'sd875496, 32'sd160952, -32'sd4110023, -32'sd535124, 32'sd1098053, -32'sd3289966, 32'sd2571186, -32'sd2343706, -32'sd1302613, 32'sd1956904, -32'sd616043, -32'sd2585434, -32'sd3896974, 32'sd410927, 32'sd1764318, 32'sd1651854, -32'sd932367, 32'sd1790240, -32'sd1872634, 32'sd2070976, 32'sd2125544, -32'sd2069484, -32'sd2206790, -32'sd3609806, -32'sd2809817, -32'sd2671408, 32'sd1892398, 32'sd2725699, -32'sd1994762, 32'sd2645791, 32'sd3826395, 32'sd3171782, -32'sd2007821, -32'sd32364, 32'sd3458260, 32'sd1292663, 32'sd1428094, -32'sd4928320, -32'sd1749114, 32'sd3753865, -32'sd731529, 32'sd2910491, 32'sd1554379, 32'sd668163, 32'sd1912379, -32'sd775907, 32'sd1349595, 32'sd1557663, -32'sd556487, 32'sd590643, -32'sd517972, -32'sd3053363, -32'sd668543, 32'sd1804844, -32'sd2148512, 32'sd2852911, 32'sd1913928, 32'sd2573273, -32'sd2613186, 32'sd867213, -32'sd1399064, 32'sd1023923, -32'sd361331, -32'sd1141900, 32'sd2830855, 32'sd1141501, 32'sd2846363, -32'sd1478141, 32'sd1333994, 32'sd465297, -32'sd2261473, -32'sd639045, -32'sd1135188, -32'sd2262637, 32'sd820317, -32'sd2341009, -32'sd175638, 32'sd2387680, 32'sd1784981, -32'sd369896, -32'sd3997748, 32'sd2364696, 32'sd3070895, -32'sd3685896, 32'sd2983590, 32'sd3808562, -32'sd2323758, -32'sd2210207, -32'sd2182464, -32'sd888466, 32'sd452201, 32'sd869440, -32'sd869117, 32'sd926942, -32'sd815665, 32'sd2261249, 32'sd448017, 32'sd2481244, -32'sd660615, -32'sd1448488, 32'sd1714525, -32'sd1737280, 32'sd2723439, -32'sd514839, 32'sd3287465, 32'sd3209632, -32'sd4105023, 32'sd2668244, 32'sd1667860, -32'sd1880662, 32'sd842744, 32'sd1585709, 32'sd754328, 32'sd2172481, 32'sd2382382, 32'sd1542790, -32'sd1976090, 32'sd4049466, 32'sd3880305, 32'sd2869332, 32'sd754954, -32'sd303326},
        '{32'sd3708218, 32'sd1835148, -32'sd1582531, -32'sd3223251, -32'sd2006689, 32'sd1834103, 32'sd116836, 32'sd343840, -32'sd1510025, 32'sd848144, 32'sd319080, 32'sd2440606, 32'sd90294, -32'sd994248, -32'sd817996, -32'sd3375866, 32'sd2333176, -32'sd169663, 32'sd1196377, 32'sd2910378, 32'sd3957472, -32'sd1013452, 32'sd2421755, -32'sd2564864, -32'sd3352474, -32'sd1557458, 32'sd3017951, 32'sd3438700, 32'sd446807, -32'sd575529, 32'sd2499592, -32'sd971495, 32'sd1722139, -32'sd3115283, -32'sd3615666, -32'sd306466, -32'sd838027, 32'sd285120, 32'sd2374580, -32'sd1233763, 32'sd489558, 32'sd1259183, 32'sd2651032, -32'sd4118009, 32'sd1264298, -32'sd284892, -32'sd1675826, 32'sd2266545, 32'sd1997583, 32'sd1219411, -32'sd3690097, -32'sd1656465, -32'sd927333, 32'sd1146322, -32'sd1567516, -32'sd3050554, -32'sd1652189, -32'sd2203685, -32'sd1307547, 32'sd3458717, -32'sd451281, -32'sd1646676, 32'sd2027009, 32'sd2298067, 32'sd3592998, -32'sd4083344, -32'sd1088878, -32'sd1288776, 32'sd3021352, 32'sd2016971, -32'sd2325096, 32'sd1219482, -32'sd7584408, 32'sd1449134, -32'sd3231348, -32'sd3940246, -32'sd2471159, 32'sd557561, -32'sd3454018, -32'sd3105504, -32'sd1728238, 32'sd3049343, -32'sd1940921, -32'sd2801796, -32'sd1535733, -32'sd585618, 32'sd4103706, 32'sd744090, -32'sd372684, -32'sd1485185, 32'sd1526949, -32'sd2822330, -32'sd3652637, 32'sd1247236, 32'sd420228, -32'sd1246069, -32'sd3762904, 32'sd3650113, 32'sd2799571, 32'sd2214248, 32'sd2407288, -32'sd1551669, -32'sd1708571, 32'sd1595657, 32'sd3077969, -32'sd960001, 32'sd668835, 32'sd1351199, 32'sd2990182, -32'sd373387, -32'sd2424828, 32'sd4517219, 32'sd391329, -32'sd1134834, -32'sd3380723, 32'sd267486, 32'sd2032648, -32'sd2377626, 32'sd4785235, 32'sd2044091, 32'sd3685779, 32'sd2447194, 32'sd100889, -32'sd3458967, -32'sd5257307, 32'sd6535, 32'sd3578144, -32'sd1811133},
        '{32'sd1271810, 32'sd910530, -32'sd1369561, -32'sd727529, 32'sd3026236, 32'sd2957774, -32'sd100072, -32'sd1464845, -32'sd2386885, -32'sd2557769, -32'sd909662, 32'sd2818972, -32'sd3820743, 32'sd1795977, 32'sd2009369, 32'sd277465, -32'sd928731, -32'sd1863150, 32'sd939222, 32'sd3372942, 32'sd592843, -32'sd1059325, 32'sd2082080, 32'sd384151, 32'sd2595662, -32'sd514364, -32'sd3465491, -32'sd2624801, 32'sd4140670, -32'sd1402766, 32'sd2402819, -32'sd1460185, -32'sd4386703, -32'sd248893, 32'sd3118630, -32'sd893446, -32'sd384237, -32'sd53861, -32'sd2096520, 32'sd3201948, -32'sd1598508, -32'sd803981, 32'sd2998233, -32'sd257562, -32'sd2928206, 32'sd2276065, -32'sd3559964, 32'sd4485852, -32'sd3586081, -32'sd1142611, -32'sd577264, 32'sd85019, 32'sd2958603, -32'sd684808, 32'sd2356383, -32'sd2630599, 32'sd1440970, -32'sd1809462, 32'sd2117348, 32'sd1029676, 32'sd2049666, -32'sd177877, -32'sd3083825, -32'sd2829887, 32'sd1238546, 32'sd3294674, 32'sd1771812, -32'sd867470, 32'sd2304387, 32'sd1759685, 32'sd250981, -32'sd2170521, -32'sd1262477, -32'sd1986701, 32'sd2736331, 32'sd3447969, 32'sd2932725, -32'sd662445, -32'sd30590, -32'sd3413668, 32'sd23326, 32'sd661994, -32'sd46905, -32'sd2003882, 32'sd2807946, 32'sd2360904, 32'sd2897349, 32'sd430660, -32'sd634988, -32'sd1046402, -32'sd3442630, -32'sd2881568, -32'sd1716771, 32'sd1637721, 32'sd2053555, 32'sd115714, 32'sd1088211, 32'sd2113894, -32'sd1436534, -32'sd340147, 32'sd2685521, 32'sd957879, -32'sd1447904, 32'sd895636, 32'sd1501678, -32'sd2872195, -32'sd1439049, 32'sd749027, 32'sd1768367, 32'sd2990783, 32'sd394989, -32'sd4020960, -32'sd99953, 32'sd1404871, 32'sd3284076, 32'sd1653783, -32'sd90923, 32'sd5037513, 32'sd3318142, -32'sd863630, -32'sd837794, 32'sd2669527, -32'sd2576206, -32'sd404894, -32'sd1620900, -32'sd783462, -32'sd1145800, 32'sd2858971},
        '{32'sd1966760, -32'sd2747398, 32'sd1672447, -32'sd2257432, 32'sd3633785, -32'sd4663888, -32'sd2716633, -32'sd985473, -32'sd2017753, -32'sd3722655, -32'sd1386970, 32'sd1791277, -32'sd1932157, -32'sd473932, -32'sd1113048, -32'sd710303, -32'sd1178052, 32'sd2489089, -32'sd842104, -32'sd199473, 32'sd106115, 32'sd2152938, 32'sd1627688, -32'sd356478, 32'sd448806, -32'sd2417664, -32'sd2701345, -32'sd1764610, -32'sd236821, 32'sd481477, 32'sd1956032, 32'sd4012941, -32'sd913455, 32'sd1207923, -32'sd671325, 32'sd801106, -32'sd4086276, -32'sd2024149, -32'sd2836106, 32'sd3051099, 32'sd2524517, 32'sd1017882, -32'sd1529770, -32'sd579197, -32'sd3604432, 32'sd2254863, -32'sd1623489, -32'sd594173, 32'sd4103830, 32'sd2263566, -32'sd2256491, -32'sd2399926, -32'sd1634102, 32'sd1408882, -32'sd727342, -32'sd4106560, -32'sd2106617, -32'sd4050000, 32'sd3018571, -32'sd1735535, -32'sd3954496, 32'sd224863, -32'sd1132885, -32'sd841214, -32'sd997580, 32'sd1152246, 32'sd1916942, -32'sd1043653, 32'sd1598426, -32'sd258209, 32'sd1686677, 32'sd841953, -32'sd566815, -32'sd1903664, -32'sd180921, 32'sd1548381, 32'sd2229269, 32'sd379471, 32'sd2400349, 32'sd2536315, 32'sd2660508, -32'sd1053420, 32'sd1683298, 32'sd824583, -32'sd2956513, 32'sd2711478, -32'sd2922743, -32'sd3583701, -32'sd2024478, 32'sd1515261, -32'sd1560338, -32'sd2803752, -32'sd1502041, -32'sd2019828, -32'sd1298946, -32'sd2977491, -32'sd557230, 32'sd2049350, 32'sd168847, 32'sd397975, -32'sd635625, -32'sd2384459, 32'sd2318497, -32'sd1073243, 32'sd837103, 32'sd2472072, 32'sd10299, 32'sd1198592, -32'sd1889133, -32'sd1877758, -32'sd26720, -32'sd1154854, 32'sd4952239, -32'sd771294, 32'sd387023, -32'sd2285153, -32'sd1282780, -32'sd1029210, 32'sd1686123, -32'sd5535511, -32'sd2259376, 32'sd1378878, -32'sd3207318, -32'sd4205276, -32'sd1724171, -32'sd1540905, 32'sd1513275, 32'sd2323969},
        '{32'sd1196991, 32'sd3459353, 32'sd66721, -32'sd1892331, -32'sd274895, -32'sd3760628, 32'sd2621665, 32'sd2345232, -32'sd2146018, -32'sd3788818, -32'sd1697993, 32'sd1573987, 32'sd1226120, 32'sd3162456, 32'sd2161991, 32'sd313430, -32'sd321567, 32'sd367717, -32'sd3294812, 32'sd1072495, 32'sd706315, 32'sd1804700, 32'sd389461, 32'sd2019285, -32'sd3139823, -32'sd2660649, 32'sd1986459, -32'sd936369, -32'sd6396252, -32'sd1440266, 32'sd974712, -32'sd1838628, 32'sd637416, -32'sd1614439, -32'sd2327092, -32'sd3007492, 32'sd3951156, -32'sd3052510, 32'sd1896043, 32'sd1987125, 32'sd31777, 32'sd1396821, -32'sd2356747, 32'sd1334969, -32'sd583357, 32'sd3149852, 32'sd925657, 32'sd1026185, -32'sd1365455, -32'sd2414615, 32'sd4531042, -32'sd842632, -32'sd2316867, -32'sd3218185, 32'sd26985, 32'sd749887, -32'sd2087560, -32'sd291665, -32'sd1392624, -32'sd1999088, 32'sd1351666, -32'sd454738, 32'sd48112, -32'sd456841, 32'sd1751271, -32'sd2421705, -32'sd1878706, -32'sd4075894, 32'sd2599181, 32'sd32109, 32'sd1890239, 32'sd2510905, 32'sd2581516, 32'sd2637933, -32'sd248905, -32'sd3063378, 32'sd2669360, 32'sd1146843, 32'sd363371, -32'sd2438808, -32'sd921997, 32'sd1866104, 32'sd2282051, 32'sd1363346, 32'sd2813847, -32'sd210481, -32'sd738116, -32'sd370000, 32'sd3240378, -32'sd2051256, 32'sd2159690, 32'sd2723393, -32'sd3517730, 32'sd1911729, 32'sd132123, 32'sd832336, -32'sd2603323, 32'sd1362099, -32'sd3752086, 32'sd2902100, -32'sd2159453, 32'sd409706, -32'sd1948500, 32'sd1590234, -32'sd2684795, 32'sd2641490, 32'sd4024928, 32'sd2819507, 32'sd1571005, 32'sd583914, 32'sd1175929, 32'sd1360445, 32'sd2613090, -32'sd1441861, 32'sd46364, 32'sd1126285, 32'sd1287933, -32'sd4099147, 32'sd1105268, 32'sd4160493, 32'sd2400651, 32'sd1338515, -32'sd4325349, -32'sd358255, 32'sd799729, -32'sd194989, 32'sd2087099, 32'sd751589},
        '{-32'sd2409028, 32'sd2517374, -32'sd1817096, 32'sd1301828, -32'sd3341464, -32'sd3108929, -32'sd2732493, -32'sd3636939, 32'sd1132211, 32'sd4015096, 32'sd1354368, 32'sd3189404, 32'sd2314459, 32'sd35259, 32'sd750890, 32'sd2267957, -32'sd3443629, -32'sd3354533, -32'sd267096, -32'sd2920066, 32'sd3231831, -32'sd2368228, 32'sd301602, 32'sd2587615, -32'sd1643619, -32'sd2560790, 32'sd1600082, -32'sd1568113, 32'sd3887139, 32'sd2462887, -32'sd631267, 32'sd552142, -32'sd1996878, -32'sd4552730, 32'sd598044, -32'sd425145, -32'sd1547951, 32'sd4163831, 32'sd2601579, -32'sd764760, -32'sd723984, -32'sd2949549, -32'sd2176884, -32'sd14602, -32'sd14635, 32'sd2615641, 32'sd6471337, -32'sd2487513, 32'sd1253820, 32'sd1301150, 32'sd1478022, -32'sd3859439, -32'sd2967853, -32'sd737856, -32'sd2923185, -32'sd2801123, 32'sd2995814, 32'sd748379, 32'sd1860208, -32'sd708891, -32'sd1457267, 32'sd1041680, 32'sd615628, 32'sd2078992, -32'sd1159825, 32'sd3817127, -32'sd485079, -32'sd720434, -32'sd1459412, 32'sd3017218, 32'sd580169, -32'sd869869, 32'sd3393196, -32'sd586089, 32'sd1367590, -32'sd1721752, -32'sd1640214, 32'sd401000, 32'sd2244389, 32'sd1612712, 32'sd2028508, 32'sd75471, 32'sd848462, -32'sd4889571, -32'sd2085323, 32'sd140968, -32'sd603388, 32'sd885456, -32'sd341156, 32'sd3530125, 32'sd522828, 32'sd25960, -32'sd1152803, -32'sd2693428, 32'sd3895061, -32'sd809848, 32'sd2184379, -32'sd2930435, 32'sd268905, 32'sd2455934, 32'sd3153570, 32'sd48495, 32'sd1732879, -32'sd1003173, 32'sd3546896, -32'sd1981408, 32'sd1968278, 32'sd1442533, -32'sd3917033, 32'sd1940087, 32'sd2440581, -32'sd1393616, -32'sd327364, -32'sd4284943, 32'sd3869168, 32'sd2480986, -32'sd3705435, 32'sd3423241, 32'sd115232, -32'sd605840, 32'sd934705, -32'sd3192715, -32'sd2126677, 32'sd3179837, 32'sd4164209, 32'sd3304688, 32'sd561290, 32'sd2802092},
        '{-32'sd4707746, 32'sd2083386, -32'sd2131988, 32'sd2497611, -32'sd1886705, 32'sd2317397, 32'sd1187911, -32'sd1516499, -32'sd4553725, 32'sd3197390, 32'sd2038826, 32'sd1925632, 32'sd362705, -32'sd1971620, 32'sd570998, -32'sd1313784, 32'sd3861184, 32'sd599432, 32'sd60048, -32'sd2643896, -32'sd3231108, -32'sd2097677, -32'sd4367923, 32'sd93999, 32'sd2895783, 32'sd2401093, 32'sd910562, -32'sd113123, 32'sd2769266, 32'sd89937, -32'sd1521085, 32'sd2382131, -32'sd3283076, -32'sd252927, 32'sd1748820, -32'sd2162997, -32'sd4051504, 32'sd2297390, -32'sd415053, -32'sd3583553, 32'sd83843, -32'sd1990570, 32'sd2165133, -32'sd1709571, -32'sd111665, 32'sd1756163, -32'sd3480740, -32'sd3748748, 32'sd2182892, 32'sd1910428, 32'sd2859850, -32'sd2652863, 32'sd1559266, 32'sd673178, 32'sd2219650, -32'sd928434, 32'sd1120442, 32'sd278963, 32'sd1709060, 32'sd2560600, 32'sd657161, 32'sd1127311, 32'sd95085, -32'sd1219894, 32'sd277370, -32'sd1747472, -32'sd2394544, 32'sd541499, 32'sd837963, 32'sd2318507, 32'sd2514808, -32'sd368716, -32'sd1345862, -32'sd2613396, -32'sd858548, 32'sd1885072, -32'sd1397301, 32'sd2724731, 32'sd3337068, -32'sd843766, -32'sd4721869, 32'sd2622647, 32'sd1501571, -32'sd4248496, 32'sd3357511, -32'sd1100937, 32'sd391054, -32'sd408116, 32'sd267768, -32'sd940013, -32'sd2200103, 32'sd1053784, -32'sd1140705, 32'sd1261822, -32'sd514913, -32'sd1780157, -32'sd2534331, -32'sd850249, -32'sd561474, -32'sd2038301, 32'sd3547180, 32'sd4006011, 32'sd1590, -32'sd4083831, -32'sd1470709, 32'sd82142, -32'sd939137, -32'sd2483319, -32'sd1961316, -32'sd2522052, 32'sd2475553, -32'sd2382752, -32'sd2615195, -32'sd2097069, 32'sd4943868, 32'sd447047, -32'sd1457582, -32'sd2102514, 32'sd1015258, -32'sd1566419, 32'sd3207349, 32'sd2268799, 32'sd502382, 32'sd968847, -32'sd201695, 32'sd801776, 32'sd1060979, 32'sd1530678},
        '{32'sd1179737, 32'sd3068269, 32'sd167987, -32'sd411043, 32'sd3914803, 32'sd4374420, -32'sd4074653, 32'sd2114128, -32'sd1632583, 32'sd1764625, 32'sd885093, -32'sd619619, 32'sd498852, -32'sd409655, -32'sd1336622, -32'sd523900, -32'sd1287421, -32'sd992457, 32'sd3325009, 32'sd2852916, 32'sd2559680, 32'sd5803942, -32'sd1545868, 32'sd2541079, -32'sd699139, -32'sd1114845, -32'sd3738942, -32'sd3835758, -32'sd414995, -32'sd39182, 32'sd2744946, -32'sd1952988, -32'sd5026146, -32'sd847395, 32'sd1272155, 32'sd2749871, 32'sd1216804, -32'sd1027477, -32'sd4178061, -32'sd480989, 32'sd3516116, 32'sd297622, -32'sd2786853, 32'sd6777, 32'sd2422079, 32'sd468449, -32'sd2114347, 32'sd1841418, 32'sd57560, 32'sd2543666, 32'sd3499771, -32'sd1081946, -32'sd542693, -32'sd1762149, 32'sd3450578, -32'sd2224944, -32'sd3457316, 32'sd481796, -32'sd317422, 32'sd2690511, -32'sd398785, -32'sd13437, 32'sd1540886, 32'sd923597, 32'sd2601842, -32'sd2448036, -32'sd1596734, 32'sd1561268, -32'sd1442815, 32'sd1692275, -32'sd1188799, -32'sd2197312, 32'sd1455678, -32'sd377022, -32'sd940354, -32'sd863671, -32'sd2910911, -32'sd541819, 32'sd2654682, 32'sd842132, -32'sd2752559, 32'sd3476470, 32'sd704966, -32'sd668706, 32'sd316936, 32'sd499014, -32'sd2523861, 32'sd2436390, -32'sd1418283, -32'sd698047, 32'sd131298, 32'sd1571502, 32'sd199412, 32'sd2114526, 32'sd1055550, 32'sd789139, 32'sd2795001, 32'sd122191, 32'sd460247, -32'sd2609767, 32'sd3197226, 32'sd1760636, -32'sd186683, 32'sd2567582, -32'sd1870412, 32'sd2776170, 32'sd1677536, -32'sd2225724, -32'sd573434, 32'sd1375716, 32'sd1520714, -32'sd2866314, 32'sd2627982, 32'sd1480838, 32'sd257166, -32'sd3616908, 32'sd3899464, 32'sd215986, 32'sd342807, -32'sd4142301, -32'sd1233480, 32'sd2071621, 32'sd2004563, 32'sd1185750, 32'sd1907334, 32'sd4085153, -32'sd3646786, 32'sd3376423},
        '{32'sd1614350, 32'sd1659293, 32'sd459818, 32'sd2932076, 32'sd3237698, 32'sd1374200, -32'sd3146872, 32'sd345767, -32'sd1758967, 32'sd1663999, -32'sd1581920, 32'sd1171380, 32'sd882124, 32'sd2510863, 32'sd2557672, -32'sd1994733, -32'sd770918, -32'sd118761, 32'sd3558515, 32'sd1630689, 32'sd135607, 32'sd3353355, 32'sd2163476, 32'sd1914241, -32'sd2916754, 32'sd193724, 32'sd1516187, 32'sd2326198, 32'sd35863, -32'sd3882627, -32'sd2787094, -32'sd1021878, 32'sd1559740, -32'sd390095, 32'sd529781, 32'sd2649230, 32'sd2151332, 32'sd145334, 32'sd33659, 32'sd3293542, 32'sd1214542, 32'sd4832876, 32'sd2641721, -32'sd1835935, 32'sd1896077, 32'sd2835233, -32'sd6186247, 32'sd3694167, -32'sd4070174, -32'sd2690051, -32'sd1329632, 32'sd1893876, 32'sd3633324, 32'sd3372078, -32'sd978527, -32'sd4517441, -32'sd1169347, -32'sd1586189, 32'sd445856, 32'sd1842872, 32'sd292728, -32'sd356627, 32'sd913219, 32'sd887911, 32'sd1524776, -32'sd824671, -32'sd3080134, 32'sd712406, 32'sd2313747, 32'sd3642940, -32'sd2590451, -32'sd4827122, -32'sd5719630, 32'sd3587857, -32'sd4394487, -32'sd2491284, -32'sd3930076, -32'sd5588742, 32'sd1609665, -32'sd1955885, 32'sd718711, 32'sd60361, 32'sd3753736, 32'sd2961509, 32'sd1363385, 32'sd49658, 32'sd470388, -32'sd2041468, 32'sd1835486, 32'sd150296, -32'sd1940095, 32'sd2003446, -32'sd2994469, 32'sd4065882, -32'sd2869794, 32'sd334163, -32'sd1070066, 32'sd1985858, -32'sd1125418, 32'sd1256778, 32'sd1907348, 32'sd2908176, -32'sd1136643, 32'sd2529637, -32'sd627140, 32'sd1515862, 32'sd2028820, -32'sd2388118, -32'sd1685511, 32'sd1664051, 32'sd598020, 32'sd753388, 32'sd1967854, 32'sd2882668, -32'sd296538, -32'sd2650351, 32'sd2274164, -32'sd798071, -32'sd1632381, 32'sd1995528, 32'sd676551, -32'sd1863321, -32'sd1570596, -32'sd122573, -32'sd1189717, 32'sd3133352, 32'sd3361182, -32'sd4688286},
        '{-32'sd3539054, 32'sd1898410, 32'sd1362396, -32'sd1497378, -32'sd1764536, 32'sd2580399, 32'sd823283, 32'sd3129595, -32'sd1686626, 32'sd542041, -32'sd3467197, -32'sd96029, -32'sd1709977, -32'sd1275589, 32'sd414811, 32'sd2267622, -32'sd2729015, 32'sd577196, 32'sd2027607, -32'sd7352, 32'sd1038508, -32'sd327629, 32'sd1751302, -32'sd350179, 32'sd4795358, 32'sd3298249, 32'sd593022, -32'sd2086939, -32'sd835162, 32'sd1741570, 32'sd472834, -32'sd3489705, -32'sd1167665, -32'sd2376860, -32'sd4324118, -32'sd677137, -32'sd475247, -32'sd3239962, 32'sd1697097, -32'sd1526691, -32'sd666031, -32'sd2383160, 32'sd378776, 32'sd1847918, 32'sd1838644, 32'sd859897, 32'sd193555, 32'sd3497148, 32'sd805259, 32'sd866459, -32'sd2175909, 32'sd3284085, -32'sd985791, -32'sd4675189, 32'sd41523, 32'sd4565454, -32'sd295321, -32'sd847437, 32'sd2562443, -32'sd1243912, 32'sd775281, 32'sd627131, -32'sd3724982, -32'sd764067, -32'sd1653706, 32'sd123019, -32'sd2229021, -32'sd4066586, -32'sd2461949, -32'sd3848258, 32'sd1424139, 32'sd761865, -32'sd3833310, 32'sd1376471, 32'sd1556500, 32'sd553511, 32'sd2112382, 32'sd2452643, -32'sd2202261, 32'sd620321, -32'sd4670156, 32'sd516264, 32'sd2111746, 32'sd1157971, 32'sd856164, -32'sd1738996, 32'sd2079918, 32'sd1460335, -32'sd3614775, 32'sd2690127, -32'sd2483039, -32'sd483679, 32'sd898504, -32'sd2143244, -32'sd3838233, -32'sd1083450, 32'sd350218, 32'sd796682, 32'sd2197709, 32'sd3685358, -32'sd1453479, -32'sd3499964, 32'sd91777, 32'sd1757272, 32'sd2238250, -32'sd1803147, 32'sd2354333, 32'sd1986420, 32'sd818107, -32'sd7161, 32'sd1262580, 32'sd3013170, 32'sd2450174, -32'sd1268311, -32'sd3449491, -32'sd3132368, 32'sd355942, 32'sd751038, -32'sd71207, 32'sd4055567, 32'sd1824719, 32'sd3409581, -32'sd220364, -32'sd2557358, -32'sd2151512, -32'sd2325983, 32'sd2478429, 32'sd1515131},
        '{-32'sd1337164, -32'sd5537475, -32'sd1049831, 32'sd3614389, 32'sd1471246, 32'sd1097504, -32'sd4888980, 32'sd531124, 32'sd3480524, -32'sd2662192, 32'sd3374708, 32'sd1528612, 32'sd940563, 32'sd1116412, 32'sd3890226, -32'sd452063, 32'sd3780529, 32'sd2204015, 32'sd342705, 32'sd2826929, 32'sd400038, 32'sd1946591, 32'sd951459, -32'sd1926941, -32'sd343528, -32'sd283703, -32'sd522898, -32'sd1879728, -32'sd2583525, 32'sd1478843, 32'sd4896670, 32'sd700982, -32'sd1684657, 32'sd1055459, 32'sd3043192, 32'sd946937, -32'sd2969933, -32'sd1809778, -32'sd3309331, 32'sd3187375, 32'sd891791, 32'sd1135504, -32'sd3489144, -32'sd437311, -32'sd4524494, 32'sd138193, -32'sd1175801, -32'sd1771721, -32'sd2212503, -32'sd2719388, -32'sd1355601, -32'sd738837, -32'sd3476523, 32'sd479615, 32'sd1653689, 32'sd142710, -32'sd2620812, -32'sd1874656, -32'sd3698086, 32'sd2063322, -32'sd1179962, -32'sd2826255, 32'sd1949791, 32'sd2398965, -32'sd1698936, -32'sd1438023, 32'sd3562690, -32'sd1484608, 32'sd1046197, 32'sd634542, 32'sd629676, 32'sd2730313, 32'sd2080302, -32'sd917301, 32'sd3140852, 32'sd1123698, -32'sd3686656, -32'sd216698, -32'sd1140901, 32'sd1606749, -32'sd1800205, -32'sd309576, 32'sd695885, 32'sd1081787, 32'sd3390200, -32'sd4233917, -32'sd925808, -32'sd2412834, -32'sd1239591, 32'sd239612, -32'sd2048774, 32'sd989567, 32'sd371630, 32'sd2333246, -32'sd1122492, -32'sd2740491, 32'sd306864, 32'sd2346944, 32'sd2980697, -32'sd2281337, 32'sd822315, 32'sd1718245, -32'sd2714536, -32'sd333322, -32'sd120222, -32'sd5475303, -32'sd1812835, 32'sd371582, 32'sd2032518, 32'sd1203440, -32'sd2615747, -32'sd347250, 32'sd4938850, -32'sd5208393, -32'sd1432367, -32'sd1719799, 32'sd2271603, -32'sd1311887, -32'sd179044, 32'sd1949699, 32'sd1874331, 32'sd2359190, 32'sd2445670, -32'sd2534942, 32'sd1787836, -32'sd1115157, -32'sd1336400, -32'sd42738},
        '{32'sd2314719, -32'sd279401, -32'sd2664536, 32'sd5067452, 32'sd4791119, -32'sd712595, -32'sd2022998, -32'sd567124, 32'sd875452, 32'sd1026294, -32'sd367256, -32'sd3371273, -32'sd1259865, -32'sd1733190, -32'sd3314740, -32'sd4893142, -32'sd4431334, 32'sd351393, -32'sd108769, -32'sd2334046, 32'sd2850266, 32'sd1134316, 32'sd3758081, -32'sd510138, 32'sd2186507, 32'sd2847226, 32'sd1814256, -32'sd769179, 32'sd1757360, -32'sd7012496, -32'sd982960, 32'sd2023984, -32'sd3139103, -32'sd673233, -32'sd1563328, -32'sd1938676, 32'sd3635046, -32'sd3537425, 32'sd75241, 32'sd1051559, 32'sd465694, -32'sd451994, -32'sd412264, -32'sd6555955, -32'sd1804530, -32'sd1412101, -32'sd4490377, 32'sd793865, 32'sd583761, 32'sd3062033, -32'sd1559121, 32'sd3116944, -32'sd728984, 32'sd3642417, -32'sd2679323, -32'sd1185809, -32'sd2934978, -32'sd3068702, -32'sd3809734, 32'sd2744019, 32'sd326400, -32'sd148573, -32'sd274996, 32'sd1426903, 32'sd699628, 32'sd513687, 32'sd1650082, -32'sd227993, -32'sd3057319, -32'sd384611, -32'sd1681133, 32'sd791094, -32'sd3793208, -32'sd2956838, -32'sd4202596, 32'sd4376983, 32'sd44438, -32'sd2024551, 32'sd1420501, -32'sd612300, -32'sd226902, 32'sd2226602, -32'sd1691186, -32'sd1438719, 32'sd1407314, 32'sd784708, -32'sd3109255, -32'sd525017, 32'sd895117, -32'sd5453825, 32'sd1713933, -32'sd3660876, 32'sd2552044, 32'sd3402251, -32'sd1093940, 32'sd1680515, 32'sd232280, 32'sd2417015, 32'sd569056, -32'sd2491901, 32'sd3041506, 32'sd1794594, 32'sd1517549, 32'sd2093542, 32'sd3309560, -32'sd1057759, -32'sd109341, 32'sd689548, 32'sd2071190, 32'sd433582, 32'sd3641724, 32'sd2554536, 32'sd399550, 32'sd2474634, -32'sd3784590, 32'sd1098691, 32'sd674738, 32'sd2242481, -32'sd2943835, -32'sd1591322, -32'sd1797434, -32'sd1292260, -32'sd3925997, 32'sd1611782, -32'sd580303, 32'sd1556519, -32'sd2763228, -32'sd3691535},
        '{-32'sd237331, 32'sd3498577, -32'sd719679, -32'sd2887165, -32'sd3128858, -32'sd2405176, 32'sd1762346, 32'sd3604008, 32'sd1119933, 32'sd622325, -32'sd644329, -32'sd1287511, -32'sd1074773, 32'sd2734064, 32'sd2262548, -32'sd494227, -32'sd455330, 32'sd3003086, -32'sd1173728, 32'sd1598691, -32'sd850119, 32'sd2330241, 32'sd3939276, 32'sd2740877, 32'sd2754922, 32'sd2514839, -32'sd1237044, 32'sd1847274, 32'sd677456, -32'sd72571, 32'sd1425365, 32'sd2122060, -32'sd558689, 32'sd408709, -32'sd1197262, 32'sd640605, -32'sd1216004, 32'sd3421708, 32'sd1940243, 32'sd1537316, -32'sd3831364, -32'sd5178174, -32'sd2709625, -32'sd1439425, -32'sd5274711, -32'sd1963396, 32'sd2785395, 32'sd1943512, -32'sd1949216, -32'sd2491058, 32'sd2006080, -32'sd1656312, -32'sd2601557, 32'sd1125289, 32'sd6381007, -32'sd231057, 32'sd2083800, -32'sd388738, 32'sd1843198, 32'sd1219558, 32'sd832971, -32'sd4781359, -32'sd731616, -32'sd3103377, -32'sd2117605, 32'sd114080, -32'sd3640061, -32'sd1963800, 32'sd2264897, -32'sd3629037, -32'sd2857387, -32'sd405330, 32'sd1817153, -32'sd3403575, 32'sd177653, 32'sd619565, 32'sd1365991, 32'sd732557, -32'sd3583462, 32'sd3315587, -32'sd1563985, 32'sd3102597, 32'sd748200, -32'sd2953344, -32'sd1929089, 32'sd890769, 32'sd1637310, 32'sd4312388, -32'sd3383835, 32'sd2306294, 32'sd2361892, -32'sd790269, 32'sd3614419, -32'sd3015648, 32'sd1731607, -32'sd2392812, 32'sd2200104, -32'sd2784657, 32'sd4024181, -32'sd754277, 32'sd11771, 32'sd2914464, -32'sd3657537, -32'sd3043394, 32'sd1199853, 32'sd611576, -32'sd1579364, 32'sd1945918, 32'sd37850, -32'sd3944078, -32'sd1457501, -32'sd4988428, 32'sd507224, 32'sd239820, -32'sd1661896, 32'sd3377896, -32'sd408396, 32'sd3640757, 32'sd1415711, 32'sd1908867, -32'sd1542795, -32'sd316343, -32'sd861370, 32'sd1890742, 32'sd719602, -32'sd2239313, -32'sd2008426, -32'sd50919},
        '{32'sd1868481, 32'sd3177886, -32'sd2993848, -32'sd1961902, 32'sd523273, -32'sd1503471, -32'sd4466171, 32'sd805136, 32'sd531587, 32'sd2602961, 32'sd1004992, -32'sd2052589, 32'sd4155590, 32'sd1283827, 32'sd2792790, -32'sd4507658, 32'sd4457260, 32'sd55089, 32'sd217228, 32'sd328604, -32'sd341688, -32'sd2510587, 32'sd1668983, -32'sd2761540, 32'sd1611501, -32'sd2818947, 32'sd2227841, -32'sd715449, -32'sd1342562, 32'sd3364180, 32'sd2043772, -32'sd437481, -32'sd2582459, -32'sd371557, 32'sd1214052, -32'sd3651035, 32'sd3280217, 32'sd1218468, 32'sd2628821, -32'sd3473806, -32'sd2675559, -32'sd2694237, -32'sd2431155, 32'sd3949119, -32'sd1657622, -32'sd2465443, 32'sd3361835, 32'sd1153135, -32'sd3183552, 32'sd446323, -32'sd2228816, 32'sd1284122, 32'sd4023181, -32'sd3565963, -32'sd4236603, -32'sd1598887, -32'sd1202025, 32'sd1937303, -32'sd2863149, -32'sd2861453, 32'sd3012164, 32'sd1627227, -32'sd1538171, 32'sd1805054, -32'sd952255, 32'sd2247164, 32'sd2024201, -32'sd2971861, -32'sd544877, 32'sd1364162, 32'sd1056538, -32'sd830066, 32'sd161120, 32'sd3324717, 32'sd1938078, 32'sd2877224, -32'sd203227, 32'sd134992, -32'sd2595006, -32'sd2668494, -32'sd1434979, -32'sd855439, 32'sd1538164, 32'sd65582, -32'sd679004, -32'sd823451, 32'sd2655836, 32'sd2048598, -32'sd1975278, -32'sd3704330, 32'sd3761417, 32'sd80800, -32'sd1370715, -32'sd2946569, -32'sd3271843, 32'sd491580, -32'sd6050526, 32'sd2425252, -32'sd1686609, 32'sd2202683, 32'sd2624401, 32'sd3656301, -32'sd611440, -32'sd340574, -32'sd3650312, 32'sd1065233, 32'sd1178845, -32'sd748723, -32'sd647819, 32'sd674060, -32'sd1981125, 32'sd2261873, -32'sd2341785, 32'sd1044105, -32'sd2268270, 32'sd1843567, -32'sd1001754, -32'sd2116343, 32'sd1718155, -32'sd2133126, 32'sd1063281, -32'sd1649419, 32'sd621521, -32'sd1480599, -32'sd3659333, -32'sd311871, 32'sd1668296, 32'sd1989411},
        '{32'sd89262, -32'sd3458129, 32'sd1104819, -32'sd2319616, 32'sd1485371, -32'sd125622, 32'sd3869222, -32'sd1085559, 32'sd1996673, 32'sd714481, 32'sd1182245, 32'sd3092581, -32'sd2999596, 32'sd2267027, -32'sd611272, -32'sd2689287, 32'sd2516746, 32'sd2613773, -32'sd426428, -32'sd2395323, 32'sd465675, -32'sd2521758, 32'sd1242502, 32'sd1288152, 32'sd2773498, -32'sd1007502, 32'sd792402, 32'sd2454172, -32'sd14854, -32'sd110324, 32'sd1436261, 32'sd312885, -32'sd1426164, -32'sd2600936, -32'sd1749363, 32'sd671834, -32'sd2241453, 32'sd2205505, -32'sd1224685, -32'sd13877, 32'sd2880231, -32'sd3040952, 32'sd762297, 32'sd3005982, -32'sd4905380, 32'sd2391286, 32'sd1372169, 32'sd1538847, 32'sd179575, -32'sd1634113, 32'sd2705124, 32'sd695724, -32'sd3155031, 32'sd2054360, 32'sd412163, 32'sd2858967, -32'sd1968829, 32'sd3425954, 32'sd2649356, -32'sd1068187, -32'sd1216204, -32'sd4784930, -32'sd991298, 32'sd2782139, -32'sd1611029, 32'sd913072, 32'sd2996084, 32'sd3665727, -32'sd1354262, 32'sd816445, 32'sd1616773, -32'sd640210, -32'sd1125280, 32'sd1084391, 32'sd3502603, 32'sd3139594, -32'sd3008688, -32'sd616895, -32'sd1948708, -32'sd141655, 32'sd2840754, 32'sd879049, -32'sd3527209, 32'sd1128775, -32'sd3561312, 32'sd2132490, 32'sd1706386, 32'sd109767, -32'sd3081890, 32'sd1306175, 32'sd3545090, -32'sd353947, 32'sd2040001, -32'sd3320551, 32'sd3175769, 32'sd978152, 32'sd577208, 32'sd3155847, 32'sd1515955, -32'sd288798, 32'sd53318, 32'sd3416606, -32'sd3246394, 32'sd327390, 32'sd1187249, 32'sd2703039, -32'sd579444, -32'sd1022650, 32'sd1715752, 32'sd267922, -32'sd674128, 32'sd1622904, 32'sd4103803, -32'sd1232485, -32'sd781226, 32'sd1618329, -32'sd893067, -32'sd3089564, 32'sd3669112, -32'sd464701, 32'sd2759889, 32'sd972612, -32'sd2073378, 32'sd232160, -32'sd270568, 32'sd1210633, -32'sd428391, -32'sd3219530}
    };

    localparam logic signed [31:0] layer1_biases [0:63] = '{
        32'sd1323763, 32'sd283564, -32'sd2519065, -32'sd633071, -32'sd391775, -32'sd484931, 32'sd2334649, 32'sd2841104, -32'sd444368, 32'sd1029247, -32'sd1998424, -32'sd3279888, 32'sd1688242, -32'sd1073175, 32'sd2327013, -32'sd502605, -32'sd1762486, 32'sd14818, -32'sd496505, 32'sd3344483, -32'sd503506, -32'sd1534096, 32'sd3159614, -32'sd631470, -32'sd3136928, 32'sd1291038, 32'sd3042584, -32'sd34918, -32'sd1340647, -32'sd1337915, 32'sd37384, -32'sd1656521, -32'sd2592211, 32'sd919961, 32'sd2499197, -32'sd1525807, 32'sd1157333, 32'sd3217006, 32'sd3725416, -32'sd2732652, 32'sd188411, 32'sd3080427, 32'sd1099557, -32'sd2646309, 32'sd2640901, 32'sd2878705, -32'sd3846477, 32'sd717378, 32'sd3815551, 32'sd708646, -32'sd7867, 32'sd2525834, -32'sd2071826, 32'sd1314560, 32'sd1228529, -32'sd588072, 32'sd3091701, 32'sd202229, 32'sd172533, -32'sd1576308, 32'sd2341765, 32'sd1020744, 32'sd3712642, -32'sd1400503
    };

    //Layer 2: 64 inputs, 10 neurons
    localparam logic signed [31:0] layer2_weights [0:9][0:63] = '{
        '{32'sd3211402, -32'sd918263, -32'sd637125, 32'sd5749780, -32'sd2272214, 32'sd1724238, -32'sd8310484, 32'sd3837882, 32'sd5260417, 32'sd3882587, -32'sd5411538, -32'sd648262, -32'sd7778050, 32'sd1642367, -32'sd2781014, -32'sd2933147, -32'sd5791443, -32'sd6445594, -32'sd6301890, -32'sd6849037, 32'sd4002711, -32'sd2206384, 32'sd2597414, 32'sd3568370, 32'sd1408406, -32'sd5776981, -32'sd661685, -32'sd2269318, 32'sd2079065, -32'sd5615581, -32'sd5805745, 32'sd3780187, -32'sd5241979, -32'sd5736268, -32'sd7050747, -32'sd5049094, -32'sd3674121, -32'sd5661537, 32'sd2613493, -32'sd3937388, 32'sd1919265, 32'sd3910816, 32'sd2091297, 32'sd1307680, -32'sd6236716, 32'sd3562641, -32'sd4936586, -32'sd6947352, -32'sd2105314, 32'sd5298115, 32'sd4264337, 32'sd6022847, -32'sd6376370, 32'sd42755, -32'sd2667035, 32'sd4420418, 32'sd5752855, 32'sd4742742, -32'sd3073993, 32'sd3120951, 32'sd5801117, -32'sd8156892, -32'sd6254310, 32'sd613947},
        '{32'sd2339677, 32'sd1750189, -32'sd3202453, 32'sd4315454, 32'sd3921228, 32'sd46725, -32'sd889183, -32'sd1424455, -32'sd871892, -32'sd6023627, -32'sd5667044, 32'sd2119383, -32'sd359010, -32'sd6985869, -32'sd5599634, 32'sd4920397, 32'sd5438179, -32'sd5365109, -32'sd4073943, 32'sd4501074, 32'sd6250426, -32'sd4631023, 32'sd177721, 32'sd5274888, 32'sd6403575, 32'sd814343, -32'sd5555555, 32'sd376865, -32'sd5665440, 32'sd5644475, -32'sd6613032, 32'sd3273425, 32'sd1375972, -32'sd2376675, -32'sd4321941, -32'sd8663346, -32'sd5449530, 32'sd2228917, -32'sd6420015, -32'sd4545873, 32'sd2480016, -32'sd4939864, 32'sd5276795, -32'sd959785, -32'sd2508200, -32'sd7220185, 32'sd3797791, -32'sd3230647, -32'sd8095569, -32'sd1663179, -32'sd432561, 32'sd3611746, -32'sd1395200, -32'sd3228687, 32'sd1907912, 32'sd2012640, 32'sd2216428, -32'sd4918087, 32'sd5925115, 32'sd1062780, -32'sd4894889, 32'sd6862252, -32'sd4597497, -32'sd2187926},
        '{32'sd507804, -32'sd2131416, 32'sd6167205, 32'sd3251093, 32'sd2660912, -32'sd5886828, 32'sd3932161, 32'sd4048981, -32'sd1349063, -32'sd3441475, -32'sd3810868, 32'sd4814447, -32'sd2396608, -32'sd116110, 32'sd1545028, 32'sd714710, -32'sd4628251, 32'sd1724219, 32'sd2742277, 32'sd5160206, -32'sd2127877, -32'sd2789247, -32'sd2916097, -32'sd2361206, -32'sd2834933, -32'sd4659853, -32'sd166907, -32'sd7836883, 32'sd1951147, -32'sd2850510, 32'sd478926, 32'sd3295204, -32'sd2726296, -32'sd4859964, -32'sd5276595, 32'sd517454, 32'sd1438294, -32'sd2774592, -32'sd1510070, 32'sd3615313, -32'sd6123629, 32'sd39878, -32'sd5428253, 32'sd4503279, 32'sd176868, 32'sd2185429, -32'sd2753549, 32'sd6100743, 32'sd3998108, -32'sd193114, 32'sd6189518, -32'sd136092, 32'sd894524, 32'sd5652080, -32'sd3253750, -32'sd5346435, -32'sd74814, 32'sd628996, 32'sd3229039, -32'sd1503070, -32'sd5903732, -32'sd2235151, 32'sd3347884, -32'sd1195116},
        '{32'sd964606, 32'sd445973, 32'sd3475807, 32'sd1905330, -32'sd7613995, 32'sd2129979, -32'sd5273047, 32'sd4706797, 32'sd2339730, -32'sd1363140, 32'sd1520399, -32'sd2229863, -32'sd5359574, 32'sd608093, -32'sd86810, -32'sd4874664, 32'sd4822016, 32'sd2631835, 32'sd5208573, -32'sd1521243, -32'sd6006070, -32'sd3486906, -32'sd6471186, 32'sd568491, -32'sd1010023, 32'sd5591604, -32'sd4281732, 32'sd3663993, 32'sd4260472, 32'sd4187581, 32'sd4972687, -32'sd5311008, -32'sd2061072, -32'sd4134793, 32'sd4716142, 32'sd3106203, -32'sd6298070, -32'sd136636, 32'sd432352, -32'sd2199311, -32'sd2760398, 32'sd5401595, 32'sd492155, 32'sd3364044, -32'sd2878290, 32'sd5606945, -32'sd5036140, -32'sd1698951, 32'sd3059383, -32'sd2086727, -32'sd5779590, 32'sd1909311, -32'sd4263972, -32'sd1788153, 32'sd620499, 32'sd2662489, -32'sd3348403, -32'sd6608742, -32'sd3049031, 32'sd695672, -32'sd4079013, 32'sd6175680, -32'sd1767598, 32'sd5481755},
        '{-32'sd964633, -32'sd1161822, -32'sd1139450, -32'sd9551696, 32'sd4173732, -32'sd2132354, -32'sd6898512, -32'sd8559887, 32'sd721789, 32'sd1335604, 32'sd3526719, -32'sd2157622, 32'sd5626385, -32'sd5751050, -32'sd7424080, 32'sd3401972, -32'sd4666025, 32'sd752649, 32'sd2647020, -32'sd185065, 32'sd4888393, -32'sd2026005, -32'sd3531561, 32'sd6074230, -32'sd1074370, -32'sd7504783, 32'sd710568, 32'sd5524019, -32'sd4827139, 32'sd2829700, 32'sd670684, 32'sd3128330, 32'sd3566901, 32'sd5517839, 32'sd870774, 32'sd963738, -32'sd350003, 32'sd326727, 32'sd5233665, -32'sd3535325, 32'sd3917653, -32'sd7981911, -32'sd1119996, 32'sd2381634, -32'sd8153498, -32'sd3111085, -32'sd6287022, 32'sd1962843, 32'sd4391315, 32'sd1504785, 32'sd3276431, -32'sd6969290, 32'sd628864, 32'sd4685037, -32'sd4075120, -32'sd6897220, -32'sd457053, -32'sd2516122, -32'sd309361, 32'sd5932700, -32'sd1115896, -32'sd216007, 32'sd3415395, 32'sd2006947},
        '{-32'sd6463844, 32'sd500834, -32'sd1360766, -32'sd550130, 32'sd851928, 32'sd2184343, 32'sd4099301, 32'sd2094673, -32'sd3437500, -32'sd820938, 32'sd2390100, 32'sd988280, 32'sd2776396, 32'sd5701704, -32'sd1335420, -32'sd5586667, -32'sd6750293, -32'sd39310, -32'sd6551592, -32'sd5590397, -32'sd205702, 32'sd4914486, 32'sd645390, 32'sd3718102, 32'sd456205, 32'sd3821658, -32'sd8312929, -32'sd1324732, -32'sd1270904, -32'sd7673190, 32'sd4078614, -32'sd3659712, 32'sd3192888, 32'sd1274482, 32'sd984436, 32'sd2262245, -32'sd1419001, 32'sd6287804, -32'sd9443360, 32'sd6040793, -32'sd583278, -32'sd1149860, 32'sd6326869, 32'sd4213376, -32'sd1565777, 32'sd1284224, 32'sd2916930, -32'sd6700072, 32'sd4377739, 32'sd3919357, -32'sd6920305, 32'sd1766385, -32'sd1590812, 32'sd174030, 32'sd3964586, -32'sd3181114, -32'sd6632481, -32'sd3580769, 32'sd4090958, -32'sd5394375, 32'sd2502496, -32'sd4292347, 32'sd4391970, -32'sd4483957},
        '{-32'sd5730425, 32'sd4163815, 32'sd714377, 32'sd606314, 32'sd4170100, 32'sd3223878, -32'sd1658919, -32'sd3098376, 32'sd5003937, 32'sd6150612, -32'sd4148025, 32'sd73893, 32'sd2604021, 32'sd4505690, 32'sd924720, -32'sd355042, -32'sd3450907, -32'sd1248164, -32'sd5844275, -32'sd658197, -32'sd464092, -32'sd5262932, 32'sd1883339, 32'sd1956036, 32'sd7411898, -32'sd794649, -32'sd5092163, -32'sd174532, 32'sd5055252, 32'sd4167668, 32'sd2352003, -32'sd3308753, -32'sd4419115, 32'sd4046475, -32'sd6872386, 32'sd4940869, 32'sd4637947, -32'sd1508843, 32'sd1199270, -32'sd5334197, -32'sd5521041, 32'sd4063479, 32'sd1877324, 32'sd3584381, -32'sd6144827, -32'sd3176764, 32'sd3493400, -32'sd2509539, -32'sd5964828, 32'sd2680145, 32'sd4241616, -32'sd3968024, 32'sd2945183, 32'sd2811199, -32'sd4884431, -32'sd1921994, -32'sd5320674, 32'sd5192635, -32'sd4676995, -32'sd4797685, -32'sd255927, 32'sd2299271, 32'sd693012, -32'sd1422184},
        '{-32'sd1381858, 32'sd4413231, 32'sd2487408, 32'sd3291666, 32'sd172156, -32'sd6448941, 32'sd4321087, -32'sd4654433, -32'sd5815665, 32'sd672592, 32'sd5729803, 32'sd732187, -32'sd3860031, -32'sd4403653, -32'sd5386107, 32'sd3410327, 32'sd4849602, -32'sd2097586, 32'sd3878168, 32'sd2690671, -32'sd1336349, -32'sd278413, -32'sd5413975, 32'sd2600049, -32'sd4793693, -32'sd1643689, -32'sd1570512, 32'sd972923, 32'sd3888483, -32'sd5223998, -32'sd5571532, 32'sd491066, -32'sd2443785, 32'sd2882914, 32'sd1157362, -32'sd290048, -32'sd1142147, -32'sd5305623, -32'sd515094, 32'sd5061132, 32'sd4971782, -32'sd2109781, 32'sd2894266, 32'sd6313805, 32'sd4871887, -32'sd1445513, 32'sd1723221, -32'sd3998885, -32'sd3842606, -32'sd4589240, -32'sd4293299, 32'sd475675, 32'sd4053528, -32'sd7106497, -32'sd4465435, -32'sd3158158, 32'sd263901, -32'sd2969532, -32'sd2993129, 32'sd3612011, 32'sd887800, 32'sd301096, -32'sd2102143, 32'sd1858371},
        '{32'sd3527100, -32'sd621809, -32'sd752447, -32'sd6623311, 32'sd6019406, -32'sd7152330, 32'sd3457698, -32'sd6962257, 32'sd4765811, 32'sd5355623, -32'sd7635840, -32'sd3815805, 32'sd5969896, 32'sd1946469, 32'sd1900058, -32'sd5772300, -32'sd3918771, -32'sd3018064, 32'sd5337061, 32'sd3016758, 32'sd3298498, 32'sd4013995, 32'sd3703933, -32'sd7460029, -32'sd4874362, -32'sd2329536, 32'sd603816, -32'sd2868384, -32'sd1503621, -32'sd5580956, 32'sd3410231, -32'sd7904340, -32'sd6048638, 32'sd3882380, 32'sd1027045, -32'sd1917507, -32'sd2892522, 32'sd932830, 32'sd4616600, 32'sd230266, 32'sd3447936, 32'sd5566602, 32'sd2715766, -32'sd7997875, -32'sd617397, -32'sd961126, -32'sd3800818, 32'sd5725404, 32'sd776042, 32'sd3207070, -32'sd3705696, -32'sd659699, -32'sd1824950, 32'sd3116999, -32'sd2640655, 32'sd276619, 32'sd2673791, -32'sd1810700, -32'sd7501195, 32'sd1099069, -32'sd1618885, -32'sd2244373, 32'sd7617273, -32'sd5312032},
        '{-32'sd1513344, -32'sd6218759, -32'sd7844244, 32'sd4975122, 32'sd3805345, 32'sd2387404, 32'sd3460036, -32'sd1576503, 32'sd4609779, -32'sd7988867, 32'sd4039194, -32'sd5158646, 32'sd4890584, 32'sd3546268, 32'sd4205380, -32'sd3421032, 32'sd1271546, -32'sd1203579, -32'sd4695495, -32'sd3087555, -32'sd487430, -32'sd2258846, -32'sd106236, -32'sd5508852, -32'sd3708761, 32'sd6111069, 32'sd4599934, 32'sd6207765, 32'sd3576413, -32'sd4103299, 32'sd1407341, 32'sd1127294, 32'sd953775, 32'sd4736510, 32'sd3193405, -32'sd5856808, 32'sd5178943, -32'sd3462708, 32'sd4737509, 32'sd2230356, 32'sd2200629, -32'sd5183642, -32'sd3827320, -32'sd6698454, -32'sd1885713, -32'sd20239, -32'sd4025901, -32'sd5675548, 32'sd415168, 32'sd5063125, -32'sd2648186, -32'sd2309977, -32'sd1747562, -32'sd794411, 32'sd3609824, 32'sd74052, 32'sd513572, -32'sd5864061, -32'sd752141, -32'sd4730420, 32'sd3807618, -32'sd1295541, -32'sd10538617, 32'sd2288457}
    };

    localparam logic signed [31:0] layer2_biases [0:9] = '{
        32'sd2500701, 32'sd173921, 32'sd1628997, -32'sd4294093, -32'sd2750769, -32'sd630976, -32'sd4443872, -32'sd5495012, 32'sd3519044, -32'sd3498747
    };


    //Intermediate outputs
    logic signed [31:0] layer0_out [0:127];
    logic signed [31:0] layer1_out [0:63];


    //Instantiate Layers
    //Layer 0
    layer #(
        .NEURONS(128),
        .PREV_LAYER_OUTPUTS(784)
    ) layer0 (
        .data_inputs(data_inputs),
        .weights(layer0_weights),
        .biases(layer0_biases),
        .data_outputs(layer0_out)
    );

    //Layer 1
    layer #(
        .NEURONS(64),
        .PREV_LAYER_OUTPUTS(128)
    ) layer1 (
        .data_inputs(layer0_out),
        .weights(layer1_weights),
        .biases(layer1_biases),
        .data_outputs(layer1_out)
    );

    //Layer 2
    layer #(
        .NEURONS(10),
        .PREV_LAYER_OUTPUTS(64)
    ) layer2 (
        .data_inputs(layer1_out),
        .weights(layer2_weights),
        .biases(layer2_biases),
        .data_outputs(data_outputs)
    );



    // Predicted class logic
    always_comb begin
        logic signed [31:0] max_val;
        max_val = data_outputs[0];
        predicted_class = '0;

        for (int i = 1; i < OUTPUTS; i++) begin
            if (data_outputs[i] > max_val) begin
                max_val = data_outputs[i];
                predicted_class = i[OUTPUT_IDX_BITS-1:0];
            end
        end
    end
endmodule
