module mlp_neural_net #(
    parameter int INPUTS           = 784,
    parameter int OUTPUTS          = 10,
    parameter int OUTPUT_IDX_BITS  = 4
) (
    input  logic signed [31:0] data_inputs  [0:INPUTS-1],
    output logic signed [31:0] data_outputs [0:OUTPUTS-1],
    output logic [OUTPUT_IDX_BITS-1:0] predicted_class
);


    //Layer 0: 784 inputs, 16 neurons
    localparam logic signed [31:0] layer0_weights [0:15][0:783] = '{
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd576437, -32'sd134934, -32'sd132625, -32'sd211687, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd42583, 32'sd417758, -32'sd455149, -32'sd785490, -32'sd79943, 32'sd1255362, 32'sd632455, 32'sd2290942, -32'sd1413618, -32'sd584377, -32'sd140943, 32'sd48516, 32'sd512141, 32'sd548504, 32'sd1474634, 32'sd1315657, 32'sd1044969, 32'sd461847, -32'sd23884, 32'sd67519, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd877736, -32'sd678181, 32'sd1258707, -32'sd1763061, 32'sd1244745, 32'sd153429, 32'sd1120537, -32'sd1974464, 32'sd1079757, 32'sd1794727, 32'sd17899, -32'sd1285147, -32'sd2882779, -32'sd2931639, -32'sd2097483, 32'sd415342, 32'sd3075134, 32'sd1759827, 32'sd1027760, 32'sd313639, 32'sd1167800, 32'sd489974, 32'sd1242402, 32'sd1188199, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1619513, 32'sd838514, -32'sd1253803, 32'sd1201391, 32'sd749510, 32'sd1081086, 32'sd812664, -32'sd175109, -32'sd538840, 32'sd847621, 32'sd1745904, 32'sd907639, 32'sd1224301, 32'sd3186722, -32'sd1892930, 32'sd961903, 32'sd763202, -32'sd900981, 32'sd159021, -32'sd2947287, 32'sd699564, -32'sd778619, 32'sd612518, -32'sd598666, 32'sd100252, 32'sd0, 32'sd0, 32'sd89037, 32'sd316483, 32'sd821300, -32'sd111111, 32'sd347529, -32'sd103190, -32'sd1095633, 32'sd1262944, -32'sd256656, -32'sd149537, 32'sd568630, 32'sd2123767, 32'sd2211442, 32'sd2648719, 32'sd4308951, 32'sd2674573, -32'sd569362, 32'sd2022966, 32'sd791136, 32'sd764593, 32'sd2329965, 32'sd2576541, -32'sd2041024, -32'sd1727640, 32'sd389439, -32'sd264502, -32'sd201380, 32'sd0, 32'sd267213, 32'sd1358724, -32'sd752563, 32'sd1452878, 32'sd511960, -32'sd992450, 32'sd970699, 32'sd956560, -32'sd2313091, 32'sd1353897, 32'sd1433358, 32'sd764700, 32'sd868081, -32'sd44658, 32'sd1048849, 32'sd1143282, 32'sd31822, 32'sd1466966, 32'sd187344, 32'sd1998966, -32'sd89824, 32'sd1227745, 32'sd1616891, 32'sd104736, 32'sd2854291, 32'sd598918, -32'sd1827489, 32'sd0, 32'sd1263953, -32'sd305768, -32'sd355697, 32'sd822392, 32'sd1601550, 32'sd2353390, -32'sd1308877, 32'sd139038, 32'sd1224923, -32'sd99370, 32'sd1112882, 32'sd2349572, 32'sd947606, 32'sd1295819, -32'sd801425, -32'sd501866, 32'sd370462, 32'sd286783, -32'sd1793577, -32'sd1572325, -32'sd43432, -32'sd318871, 32'sd635523, -32'sd713453, -32'sd2642037, -32'sd2005130, 32'sd175721, 32'sd2113293, -32'sd490783, 32'sd1233970, -32'sd348335, -32'sd301326, -32'sd243407, -32'sd1091916, -32'sd1203840, 32'sd1302216, -32'sd910597, 32'sd944096, 32'sd338265, 32'sd2672203, 32'sd2034337, 32'sd1098223, 32'sd502477, 32'sd1703983, -32'sd730020, -32'sd1066284, -32'sd230781, 32'sd71899, -32'sd531495, 32'sd942387, 32'sd161689, 32'sd671002, 32'sd544786, 32'sd714157, 32'sd1123546, 32'sd946177, -32'sd1446098, 32'sd638869, -32'sd459341, 32'sd1385236, -32'sd505317, -32'sd461771, -32'sd1382199, -32'sd236257, 32'sd1544834, -32'sd14865, 32'sd625281, 32'sd2038995, -32'sd60363, 32'sd143589, 32'sd1732870, 32'sd518881, 32'sd337050, 32'sd1199738, 32'sd3418530, 32'sd498131, 32'sd185810, 32'sd1345206, -32'sd1386992, 32'sd2355623, -32'sd3198512, -32'sd2784435, 32'sd1337640, 32'sd915069, 32'sd973154, 32'sd1479041, -32'sd243936, 32'sd1512378, 32'sd600473, -32'sd169491, 32'sd1546191, 32'sd539798, -32'sd266165, -32'sd594726, -32'sd1626386, 32'sd499394, 32'sd473019, 32'sd1091250, 32'sd2895943, 32'sd1717317, 32'sd5115137, 32'sd1918845, -32'sd52355, 32'sd2985172, 32'sd627046, 32'sd2694672, 32'sd1396556, -32'sd2420841, -32'sd1153067, -32'sd3172506, 32'sd1825109, -32'sd83502, -32'sd893196, 32'sd87449, 32'sd1761045, -32'sd284974, -32'sd118824, 32'sd276592, 32'sd19243, -32'sd968396, -32'sd3420212, -32'sd1834175, -32'sd1719151, -32'sd2089917, -32'sd480584, 32'sd250894, -32'sd778700, 32'sd2857957, 32'sd1744816, 32'sd2231533, 32'sd1363709, 32'sd1168925, 32'sd114697, 32'sd973645, 32'sd594652, -32'sd186680, -32'sd1421922, -32'sd376596, 32'sd295110, 32'sd166036, -32'sd118225, -32'sd1326, 32'sd2273663, 32'sd1445017, -32'sd2683058, -32'sd573188, -32'sd1179762, -32'sd1467663, -32'sd2221296, -32'sd3479385, -32'sd653893, 32'sd698025, 32'sd1008779, 32'sd729752, -32'sd1324095, -32'sd281313, 32'sd897304, 32'sd1086695, -32'sd429042, 32'sd438108, -32'sd7953, -32'sd920917, -32'sd1384828, -32'sd1642568, 32'sd1045966, 32'sd1578386, 32'sd1821093, 32'sd311723, -32'sd214347, -32'sd2893766, -32'sd762750, -32'sd2388308, -32'sd1458051, -32'sd1000075, -32'sd1850335, -32'sd1227108, -32'sd349994, 32'sd361060, 32'sd659262, 32'sd1772371, 32'sd2764752, 32'sd956401, 32'sd276317, 32'sd183048, -32'sd95594, 32'sd473653, -32'sd2302206, 32'sd361536, -32'sd3790884, -32'sd841665, -32'sd771407, -32'sd2892655, -32'sd1062438, 32'sd1143925, -32'sd1572051, 32'sd189914, -32'sd463164, -32'sd336336, 32'sd127972, -32'sd400824, 32'sd798888, -32'sd1087870, -32'sd696612, -32'sd969982, 32'sd1002581, -32'sd379306, 32'sd1469003, 32'sd3650253, 32'sd2552995, 32'sd2383893, -32'sd250381, 32'sd1830490, -32'sd281264, 32'sd117591, -32'sd2313352, -32'sd2567031, -32'sd956239, -32'sd1767399, -32'sd722065, -32'sd277698, 32'sd106851, -32'sd277902, -32'sd2425869, 32'sd617694, 32'sd1306023, -32'sd426246, 32'sd1770743, -32'sd2342036, -32'sd1482096, 32'sd1010482, 32'sd1788340, 32'sd1556363, 32'sd633570, 32'sd1365823, 32'sd724759, 32'sd2632339, 32'sd345873, -32'sd613570, -32'sd1171209, 32'sd65256, -32'sd1121492, -32'sd1860404, -32'sd2583436, -32'sd1329645, 32'sd1652823, -32'sd1088141, 32'sd498754, -32'sd178099, 32'sd248205, 32'sd219780, -32'sd295359, -32'sd1392370, 32'sd1165048, -32'sd154710, 32'sd761220, -32'sd1276159, -32'sd1563138, -32'sd1834464, -32'sd2826662, -32'sd1937011, -32'sd89463, 32'sd1680065, 32'sd2884492, 32'sd880226, -32'sd45486, 32'sd190363, -32'sd1174376, 32'sd543959, -32'sd1040263, -32'sd1889539, 32'sd835679, 32'sd747175, 32'sd1332546, 32'sd2271882, 32'sd1165290, -32'sd3200718, 32'sd920191, 32'sd1024809, 32'sd301660, 32'sd280761, -32'sd943226, 32'sd1811297, 32'sd818581, 32'sd251478, -32'sd1021043, -32'sd2191094, -32'sd3352995, -32'sd4805939, -32'sd2751949, 32'sd1406202, 32'sd184247, 32'sd2301009, 32'sd134255, -32'sd569585, -32'sd4225718, -32'sd1291273, -32'sd791163, 32'sd1602698, 32'sd1023639, -32'sd112297, 32'sd2332125, 32'sd1857318, 32'sd2207781, 32'sd3029700, -32'sd1843354, 32'sd1238321, -32'sd171613, 32'sd0, 32'sd1185125, 32'sd188813, -32'sd143418, 32'sd797682, -32'sd2466598, -32'sd6070751, -32'sd6437010, -32'sd7559187, -32'sd4932734, -32'sd6189825, -32'sd6298088, -32'sd5611312, -32'sd2903608, -32'sd3053259, 32'sd318795, -32'sd2898941, -32'sd1520478, 32'sd1147605, 32'sd1176573, -32'sd229981, 32'sd1029657, 32'sd439110, 32'sd1115461, 32'sd428521, -32'sd4677047, -32'sd1066537, 32'sd389012, 32'sd243409, -32'sd48773, 32'sd111777, 32'sd1338330, 32'sd170717, -32'sd931485, -32'sd2437846, -32'sd2276995, -32'sd3406678, -32'sd8577099, -32'sd7543485, -32'sd13373582, -32'sd10311574, -32'sd6124780, -32'sd1419008, -32'sd1419309, 32'sd751889, 32'sd1775179, -32'sd216575, 32'sd1864044, 32'sd825619, 32'sd1895580, 32'sd2158423, -32'sd1107650, -32'sd2219959, -32'sd4435480, -32'sd391453, 32'sd119799, 32'sd236459, -32'sd441921, 32'sd130327, 32'sd1143681, -32'sd902788, -32'sd1177939, -32'sd29790, 32'sd91289, -32'sd1283570, -32'sd1561769, -32'sd1825055, -32'sd6092668, -32'sd6059000, -32'sd3277433, -32'sd522876, -32'sd292634, -32'sd805932, 32'sd2402242, 32'sd557501, -32'sd1204413, 32'sd21794, 32'sd696852, -32'sd1940151, -32'sd21733, -32'sd855472, -32'sd2672811, 32'sd92924, -32'sd643715, 32'sd0, 32'sd363934, 32'sd285000, 32'sd46950, 32'sd895208, 32'sd1500088, 32'sd2511832, 32'sd1774142, 32'sd2696444, 32'sd2407343, 32'sd975839, -32'sd124478, -32'sd1019793, -32'sd1437819, -32'sd428553, -32'sd2111342, -32'sd2832085, -32'sd1097631, -32'sd1647153, -32'sd624490, 32'sd298169, 32'sd569813, 32'sd108775, 32'sd510298, -32'sd880619, -32'sd4498988, -32'sd637024, -32'sd228131, -32'sd591983, 32'sd1362340, 32'sd897015, 32'sd1052332, 32'sd1405271, -32'sd340988, 32'sd1153721, 32'sd3119165, 32'sd2509817, 32'sd2123072, 32'sd3538117, 32'sd2520541, 32'sd2591781, 32'sd1237188, 32'sd556227, -32'sd393105, 32'sd1569912, -32'sd838887, -32'sd397917, 32'sd996269, -32'sd347676, 32'sd26528, -32'sd570528, 32'sd1704927, -32'sd2527912, -32'sd137336, 32'sd715663, 32'sd228091, 32'sd114301, 32'sd1060895, 32'sd1824716, 32'sd9664, 32'sd740165, 32'sd1041851, 32'sd127903, 32'sd2065174, 32'sd3205240, 32'sd1601897, 32'sd3275079, 32'sd3823218, 32'sd1575022, 32'sd2052258, 32'sd839359, 32'sd669865, -32'sd551236, -32'sd506311, -32'sd131500, -32'sd1101061, 32'sd276231, -32'sd329951, 32'sd1096111, -32'sd730240, -32'sd965213, -32'sd1081143, 32'sd750019, -32'sd61293, 32'sd0, 32'sd2026874, 32'sd1294275, -32'sd196620, -32'sd384732, 32'sd406554, 32'sd274044, 32'sd3590138, 32'sd446083, 32'sd1194331, 32'sd3210004, 32'sd3550329, 32'sd485407, 32'sd597475, 32'sd144163, 32'sd1261160, -32'sd497534, 32'sd914705, -32'sd605260, -32'sd225118, -32'sd322326, -32'sd1739569, -32'sd1318044, 32'sd356489, -32'sd289241, -32'sd1729817, -32'sd28503, 32'sd0, 32'sd0, 32'sd0, 32'sd22375, -32'sd177804, 32'sd1513535, -32'sd663683, 32'sd1185131, 32'sd1743428, 32'sd733624, 32'sd964003, 32'sd2870425, -32'sd40204, -32'sd1790474, 32'sd855601, 32'sd344669, 32'sd1711783, -32'sd766275, 32'sd727308, -32'sd1212356, -32'sd1059611, -32'sd1049519, -32'sd155216, -32'sd1381745, 32'sd501976, 32'sd1396345, -32'sd1101011, -32'sd600647, 32'sd0, 32'sd0, 32'sd0, 32'sd811375, -32'sd753793, 32'sd115777, 32'sd218906, -32'sd162175, 32'sd731432, 32'sd706894, -32'sd1569278, 32'sd1260543, 32'sd1565596, 32'sd333982, 32'sd1058776, -32'sd1425757, -32'sd643486, -32'sd34857, 32'sd501521, -32'sd359733, -32'sd692194, -32'sd950562, -32'sd475228, 32'sd477558, -32'sd588867, -32'sd471938, -32'sd44235, -32'sd144052, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1654194, 32'sd564224, 32'sd694703, -32'sd1196933, -32'sd427790, -32'sd223208, 32'sd1169424, 32'sd1598605, -32'sd179674, 32'sd1686965, 32'sd2562916, 32'sd2385375, -32'sd833104, -32'sd335033, 32'sd1093580, 32'sd1305397, 32'sd514337, 32'sd1723817, 32'sd3403777, -32'sd1360187, -32'sd222952, 32'sd795630, -32'sd65426, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd529721, -32'sd1227489, 32'sd1094041, 32'sd736958, -32'sd278006, -32'sd410573, 32'sd1391695, 32'sd884725, -32'sd1512482, 32'sd1962144, 32'sd1609668, -32'sd780963, 32'sd12350, -32'sd145897, 32'sd1356122, 32'sd206619, 32'sd1911933, 32'sd645767, -32'sd1053444, 32'sd1477142, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd306247, -32'sd271355, -32'sd572795, -32'sd709412, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd29781, -32'sd236101, -32'sd2068351, -32'sd71680, -32'sd1358665, -32'sd433339, 32'sd2035516, 32'sd1042335, 32'sd1815241, -32'sd610553, -32'sd571421, 32'sd1328640, 32'sd1204668, 32'sd2037390, 32'sd126283, -32'sd79843, -32'sd757056, -32'sd533267, 32'sd292084, -32'sd381145, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1206448, 32'sd680366, 32'sd1349831, -32'sd370439, 32'sd132605, 32'sd1543234, 32'sd1773717, 32'sd1299382, 32'sd11779, 32'sd1551377, 32'sd2751530, 32'sd1181272, -32'sd1045036, 32'sd1676251, 32'sd18599, 32'sd2060556, 32'sd1534657, 32'sd40414, 32'sd1123615, 32'sd1577645, -32'sd1110627, 32'sd264836, -32'sd1424433, 32'sd846834, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2935895, 32'sd362755, -32'sd424118, 32'sd2404560, 32'sd859459, -32'sd1401778, 32'sd2268817, 32'sd391066, -32'sd396937, -32'sd616783, 32'sd2448732, 32'sd2929472, -32'sd702362, 32'sd510062, 32'sd1727948, -32'sd459576, 32'sd713846, 32'sd1825100, 32'sd628771, -32'sd2358126, -32'sd639504, 32'sd674270, 32'sd1363523, -32'sd5109883, 32'sd11177, 32'sd0, 32'sd0, 32'sd398578, 32'sd15921, -32'sd576075, -32'sd597473, 32'sd842315, 32'sd22361, 32'sd72769, 32'sd2976990, 32'sd2137633, 32'sd4044605, 32'sd2095603, 32'sd1584435, 32'sd893448, -32'sd550583, -32'sd138529, 32'sd696269, -32'sd1890497, 32'sd1124433, 32'sd2438989, 32'sd130567, -32'sd585992, -32'sd2296530, -32'sd998448, 32'sd965623, -32'sd644501, 32'sd209235, -32'sd1190078, 32'sd0, 32'sd740249, 32'sd835318, 32'sd1586952, 32'sd548183, -32'sd1524023, -32'sd640286, 32'sd754055, -32'sd3509694, -32'sd309156, -32'sd2601277, -32'sd3134609, -32'sd4117, 32'sd1929574, 32'sd470990, 32'sd1658948, 32'sd95460, -32'sd2268624, 32'sd1917428, 32'sd1340957, -32'sd2044050, 32'sd388715, -32'sd413103, -32'sd651664, -32'sd1368498, -32'sd631819, 32'sd774533, -32'sd911400, 32'sd0, 32'sd891353, 32'sd1140880, 32'sd1658569, 32'sd620718, 32'sd286875, 32'sd2059425, -32'sd524747, -32'sd1136486, -32'sd703784, -32'sd1877146, 32'sd1962633, 32'sd114746, -32'sd483110, 32'sd1281221, -32'sd1511641, -32'sd1155331, -32'sd1869676, 32'sd115573, -32'sd767406, -32'sd1420661, -32'sd2197585, 32'sd1456510, 32'sd1899081, 32'sd1107709, 32'sd664234, 32'sd972864, -32'sd494471, 32'sd2662832, 32'sd357988, 32'sd1320198, 32'sd1783881, 32'sd2236858, -32'sd1481057, -32'sd1090267, -32'sd566618, -32'sd88268, -32'sd1936077, -32'sd928001, -32'sd273701, -32'sd1327418, -32'sd1994440, 32'sd579310, 32'sd458171, -32'sd4363728, -32'sd3545223, -32'sd3084418, -32'sd2846023, -32'sd91033, -32'sd2426400, -32'sd1014637, 32'sd157177, -32'sd265231, -32'sd946974, 32'sd130440, -32'sd3556374, 32'sd1567919, 32'sd1765935, -32'sd1032518, -32'sd437757, -32'sd1927762, -32'sd112284, -32'sd20268, -32'sd1049708, -32'sd443757, -32'sd2680389, -32'sd1394129, -32'sd1911983, -32'sd2671716, -32'sd3136928, -32'sd1004779, -32'sd1423043, -32'sd3542752, -32'sd1726890, -32'sd2513485, -32'sd3252126, 32'sd2594073, -32'sd609391, 32'sd202273, -32'sd323277, 32'sd716354, 32'sd1703292, 32'sd438149, 32'sd371187, 32'sd123252, -32'sd1124441, 32'sd2229093, -32'sd912458, 32'sd1278431, 32'sd1295930, -32'sd2895586, -32'sd747412, -32'sd2305661, -32'sd3472327, -32'sd1591659, -32'sd2912821, -32'sd611104, -32'sd1501221, 32'sd491738, -32'sd2418096, -32'sd1562637, -32'sd1551244, 32'sd910023, -32'sd2456197, -32'sd1368135, -32'sd893688, -32'sd1072670, -32'sd4027986, -32'sd693631, 32'sd830826, 32'sd1361559, -32'sd535272, -32'sd378979, -32'sd301034, -32'sd2479773, 32'sd989174, 32'sd1934672, 32'sd2962832, -32'sd1601041, 32'sd1045039, 32'sd1827341, -32'sd1439687, -32'sd3758756, -32'sd1760178, -32'sd547352, -32'sd1788755, 32'sd1001349, 32'sd2234235, 32'sd5161518, 32'sd350974, 32'sd91915, 32'sd1588089, 32'sd2478126, 32'sd569259, -32'sd1857403, -32'sd1080687, -32'sd204949, 32'sd1581035, 32'sd982380, -32'sd2448499, 32'sd277593, -32'sd1826594, 32'sd1688535, 32'sd304545, 32'sd1612726, 32'sd149330, -32'sd209191, 32'sd278267, -32'sd2046001, -32'sd3503499, -32'sd4119394, -32'sd1650374, -32'sd5611630, -32'sd3009120, 32'sd3016369, 32'sd849411, 32'sd2153296, -32'sd454990, -32'sd559194, 32'sd2029390, 32'sd1452949, -32'sd485893, -32'sd2125075, 32'sd67241, -32'sd1442125, 32'sd526605, -32'sd281898, 32'sd1178119, 32'sd412739, 32'sd19202, 32'sd368042, -32'sd3590624, -32'sd1142416, -32'sd2910950, -32'sd4036341, -32'sd2281337, -32'sd3014238, -32'sd1187500, -32'sd2819430, -32'sd2448709, 32'sd534981, 32'sd1298403, 32'sd3738382, 32'sd1006722, 32'sd3612415, 32'sd342805, -32'sd290353, -32'sd736611, -32'sd2080224, 32'sd1173061, -32'sd2208429, -32'sd3162014, -32'sd595030, -32'sd9407, 32'sd459964, -32'sd231106, 32'sd1390721, -32'sd987445, -32'sd116841, -32'sd1115814, -32'sd4871494, -32'sd5004222, -32'sd4141986, -32'sd4146403, -32'sd1698877, -32'sd686325, 32'sd2576615, 32'sd84432, 32'sd2694321, 32'sd4300867, 32'sd1699835, -32'sd50212, 32'sd2777417, 32'sd720140, 32'sd472274, -32'sd244579, -32'sd934063, -32'sd588507, 32'sd259560, 32'sd259720, 32'sd1694302, -32'sd1210502, -32'sd608119, -32'sd337038, 32'sd1479640, -32'sd946471, -32'sd36519, 32'sd1308753, 32'sd82130, -32'sd2955356, 32'sd1715334, -32'sd296927, -32'sd1174782, 32'sd1484759, 32'sd1663796, 32'sd692148, 32'sd909626, 32'sd3059587, 32'sd3830581, -32'sd651994, -32'sd796069, -32'sd1798321, 32'sd2276207, 32'sd151740, -32'sd758438, 32'sd801466, 32'sd162986, 32'sd676346, 32'sd1136715, 32'sd647993, 32'sd1088737, -32'sd2237511, -32'sd1567844, 32'sd790678, 32'sd1128072, 32'sd312473, 32'sd1879940, 32'sd4134920, 32'sd3908615, 32'sd306208, -32'sd418671, -32'sd1955926, 32'sd339223, -32'sd2474914, 32'sd2370, 32'sd4740901, 32'sd2844319, 32'sd482854, 32'sd404318, -32'sd772202, 32'sd1863880, 32'sd2156712, 32'sd1025384, 32'sd492789, -32'sd1321670, 32'sd2295555, 32'sd3869205, -32'sd472702, -32'sd1917727, -32'sd1056854, 32'sd209795, 32'sd592697, -32'sd1135004, 32'sd1886348, 32'sd2386109, 32'sd2479089, 32'sd1563679, 32'sd1947641, -32'sd3385443, -32'sd2749124, -32'sd786512, -32'sd2093641, -32'sd3305, 32'sd1616673, 32'sd4569037, 32'sd1238640, 32'sd2248422, 32'sd2452940, 32'sd1586203, -32'sd2159380, 32'sd2249775, 32'sd895311, 32'sd732332, 32'sd313902, 32'sd1301069, 32'sd583544, 32'sd589106, 32'sd1279832, 32'sd0, 32'sd1838090, 32'sd379376, 32'sd1258314, 32'sd1525802, 32'sd2808105, 32'sd4149730, 32'sd5370803, -32'sd361864, -32'sd1625191, 32'sd659857, -32'sd685794, -32'sd3234275, -32'sd3402848, 32'sd494844, -32'sd896282, 32'sd672083, 32'sd1982295, 32'sd320397, -32'sd600380, 32'sd101808, -32'sd148110, 32'sd351542, 32'sd877062, -32'sd1538968, 32'sd420364, 32'sd399359, 32'sd100206, -32'sd1324192, -32'sd731888, -32'sd1556002, 32'sd2717794, 32'sd1636788, 32'sd2425390, 32'sd2387221, 32'sd1843317, 32'sd1960322, -32'sd331910, 32'sd2409827, 32'sd983240, 32'sd1573901, 32'sd1198114, 32'sd554198, -32'sd415096, 32'sd471352, 32'sd1856988, -32'sd383696, 32'sd1190029, 32'sd64180, 32'sd832503, -32'sd461155, -32'sd519136, -32'sd455922, 32'sd1755464, -32'sd141916, 32'sd1750098, 32'sd794394, 32'sd1327319, 32'sd842995, -32'sd492174, -32'sd610618, 32'sd571786, 32'sd424669, 32'sd229222, 32'sd458305, -32'sd1134174, 32'sd1510255, 32'sd960673, 32'sd864596, 32'sd2602743, 32'sd2629568, 32'sd1395451, -32'sd1996528, 32'sd678696, 32'sd2902844, -32'sd217074, -32'sd406810, 32'sd435513, 32'sd2367484, -32'sd411188, -32'sd3342197, 32'sd796110, 32'sd3171507, 32'sd1215699, 32'sd0, -32'sd44985, 32'sd1047223, -32'sd1360649, -32'sd2656422, 32'sd2765231, 32'sd874151, -32'sd939138, 32'sd257033, 32'sd2030693, 32'sd3285941, 32'sd560950, -32'sd542088, 32'sd1548242, 32'sd2895730, 32'sd396425, -32'sd476788, -32'sd2497291, 32'sd1107083, -32'sd185069, 32'sd466755, 32'sd1044518, 32'sd353500, 32'sd287886, -32'sd352135, -32'sd614824, 32'sd732794, -32'sd32139, 32'sd582983, -32'sd286670, 32'sd221752, -32'sd1809019, -32'sd5582394, -32'sd1243632, -32'sd1052862, 32'sd386875, -32'sd13071, 32'sd1155553, 32'sd2074579, -32'sd1355391, 32'sd679703, -32'sd138610, 32'sd287143, -32'sd2093193, -32'sd2687300, -32'sd261837, 32'sd21848, -32'sd693471, -32'sd2115915, 32'sd107260, 32'sd319222, 32'sd475325, -32'sd1596826, 32'sd2372702, -32'sd588061, -32'sd175426, 32'sd1283929, 32'sd1752306, -32'sd152702, -32'sd372948, -32'sd4026253, -32'sd1195643, 32'sd830063, 32'sd807024, 32'sd323520, 32'sd2056594, -32'sd285111, -32'sd287697, -32'sd1222307, 32'sd1449968, -32'sd1785114, -32'sd693072, 32'sd604670, -32'sd1193854, 32'sd1760917, -32'sd2694898, -32'sd2246832, -32'sd1681759, -32'sd2527453, -32'sd764605, -32'sd516848, 32'sd587733, 32'sd683074, 32'sd1775760, 32'sd0, 32'sd2431313, 32'sd873801, 32'sd1016972, 32'sd1151603, 32'sd965561, 32'sd160404, -32'sd1425939, -32'sd1800075, 32'sd1399286, 32'sd722796, -32'sd1393137, 32'sd486095, -32'sd1624819, -32'sd4780521, -32'sd4151435, -32'sd4592336, -32'sd1173941, -32'sd1774645, -32'sd1995712, -32'sd3577103, -32'sd92656, 32'sd2145716, 32'sd345591, -32'sd1511999, -32'sd1928726, 32'sd1510731, 32'sd0, 32'sd0, 32'sd0, -32'sd613877, 32'sd8494, -32'sd472130, 32'sd759088, -32'sd160376, -32'sd886362, -32'sd2066064, -32'sd799811, -32'sd1816680, -32'sd3864174, -32'sd3661197, -32'sd7425063, -32'sd6276666, -32'sd2811749, -32'sd3299551, -32'sd1697914, -32'sd6895758, -32'sd4924156, -32'sd1669576, 32'sd2000633, 32'sd945083, -32'sd1887191, -32'sd1762112, -32'sd662080, -32'sd1056083, 32'sd0, 32'sd0, 32'sd0, 32'sd1053687, 32'sd268239, -32'sd864203, -32'sd1776673, -32'sd11486, -32'sd4071404, -32'sd193198, -32'sd931099, -32'sd4615269, -32'sd3302724, -32'sd602634, -32'sd3571952, -32'sd4096032, -32'sd5139980, -32'sd2231392, 32'sd717691, 32'sd1290889, -32'sd607437, -32'sd844721, -32'sd52169, -32'sd4101767, -32'sd854630, -32'sd3175425, 32'sd904077, 32'sd2502324, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd604447, -32'sd12547, -32'sd852435, -32'sd2172536, -32'sd505024, -32'sd422466, -32'sd1245836, -32'sd1925639, 32'sd395435, -32'sd2689487, -32'sd3170464, 32'sd925725, 32'sd2123987, 32'sd458752, -32'sd2720657, -32'sd427050, 32'sd494956, 32'sd1165003, 32'sd1026128, 32'sd480121, -32'sd11623, 32'sd1156649, 32'sd501029, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd86578, -32'sd266276, 32'sd117750, 32'sd274998, -32'sd98079, -32'sd210178, -32'sd1171166, -32'sd53283, 32'sd224346, 32'sd1112811, 32'sd424324, 32'sd894532, 32'sd219444, -32'sd156179, -32'sd795963, 32'sd208825, -32'sd109491, 32'sd699808, -32'sd812087, 32'sd456056, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd456708, -32'sd1090784, -32'sd3964742, -32'sd3975066, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd341565, 32'sd347496, -32'sd649723, -32'sd743358, -32'sd2905886, -32'sd5323499, -32'sd2385796, -32'sd1665544, -32'sd2486119, -32'sd1524555, -32'sd1356730, -32'sd3367533, -32'sd428121, -32'sd516040, -32'sd680827, -32'sd1375453, -32'sd168624, 32'sd39127, -32'sd4462101, -32'sd3654244, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5231230, -32'sd4817741, -32'sd489805, -32'sd2631338, -32'sd78657, 32'sd1062549, -32'sd492077, -32'sd3062571, -32'sd765918, 32'sd720347, -32'sd2914371, -32'sd3876626, -32'sd956474, -32'sd2511268, 32'sd162057, 32'sd631049, -32'sd83395, 32'sd90199, -32'sd1031601, -32'sd2312785, -32'sd890830, -32'sd3320959, -32'sd4015689, -32'sd3615543, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3820344, -32'sd4932556, -32'sd1977473, -32'sd2578658, 32'sd1112671, -32'sd2814550, -32'sd5037010, -32'sd1821576, -32'sd4551422, -32'sd4643084, -32'sd6127608, -32'sd5728725, -32'sd1965553, 32'sd784294, 32'sd825013, 32'sd1737710, 32'sd1941340, 32'sd2456108, 32'sd599491, -32'sd1802633, -32'sd1266427, -32'sd727362, -32'sd358896, 32'sd1060840, -32'sd5359080, 32'sd0, 32'sd0, -32'sd3577374, 32'sd1169793, 32'sd1519599, 32'sd6256, 32'sd387255, -32'sd2289397, -32'sd1783205, -32'sd374914, -32'sd2045906, -32'sd291834, -32'sd2246231, 32'sd1169850, -32'sd1023761, 32'sd140881, 32'sd706934, 32'sd4232107, 32'sd2722562, 32'sd1606783, 32'sd2412414, 32'sd4235085, 32'sd2471421, 32'sd1801244, -32'sd2002575, -32'sd150968, -32'sd2547413, 32'sd1446236, -32'sd5217490, 32'sd0, -32'sd3018529, -32'sd3320164, 32'sd475795, 32'sd2215864, 32'sd3060800, -32'sd416838, 32'sd902686, -32'sd1839820, 32'sd1587604, 32'sd1518648, 32'sd1476170, 32'sd1478834, -32'sd2942164, -32'sd3093980, -32'sd3284784, -32'sd245995, 32'sd659445, 32'sd248403, -32'sd313004, 32'sd13191, -32'sd259003, 32'sd2382150, 32'sd1192835, 32'sd3086413, 32'sd2013739, -32'sd525076, -32'sd5391921, 32'sd0, 32'sd469982, 32'sd672311, 32'sd1625699, 32'sd822013, -32'sd320454, -32'sd227325, 32'sd733644, -32'sd1847059, -32'sd526103, -32'sd645377, -32'sd92734, -32'sd481392, -32'sd2908248, -32'sd4495926, -32'sd5151208, -32'sd2601238, -32'sd1104600, -32'sd1025026, 32'sd2137054, 32'sd2517538, 32'sd2560535, -32'sd1105858, 32'sd228921, 32'sd44988, 32'sd769170, -32'sd444658, 32'sd1075640, -32'sd2957680, 32'sd900578, -32'sd392683, -32'sd446433, -32'sd343110, -32'sd1658262, 32'sd1936147, 32'sd4121791, 32'sd75720, 32'sd1461399, -32'sd328367, -32'sd703902, -32'sd1320106, -32'sd3786241, -32'sd5315945, -32'sd3740611, -32'sd1010753, 32'sd1987724, 32'sd1730348, 32'sd1779265, 32'sd3264283, 32'sd601751, 32'sd1129925, -32'sd2588423, -32'sd3126455, 32'sd1348346, -32'sd1786779, -32'sd302154, -32'sd5197708, 32'sd1164050, -32'sd311052, 32'sd1971116, 32'sd2083442, 32'sd1716045, 32'sd1646612, 32'sd2942680, 32'sd253420, 32'sd1110652, 32'sd1556016, 32'sd1822958, -32'sd820067, -32'sd2560932, -32'sd5851027, -32'sd3599636, -32'sd1393584, 32'sd631136, 32'sd3264837, 32'sd1617888, -32'sd781995, -32'sd177683, 32'sd341164, -32'sd1599488, -32'sd6931567, -32'sd1049269, -32'sd1746892, 32'sd212160, 32'sd1484360, 32'sd2768581, 32'sd1303861, 32'sd2091891, 32'sd1233314, 32'sd613479, 32'sd689879, 32'sd1023245, -32'sd756372, -32'sd369225, -32'sd1609820, -32'sd1995920, -32'sd333810, -32'sd3430378, -32'sd4534305, -32'sd719642, 32'sd124042, 32'sd1008170, 32'sd578046, -32'sd184784, 32'sd3490439, 32'sd1048232, -32'sd2560503, -32'sd1922998, -32'sd6871387, -32'sd2303008, -32'sd3757859, -32'sd3204032, 32'sd785664, 32'sd2178400, 32'sd1681430, 32'sd2035961, 32'sd1328215, -32'sd1057427, -32'sd289866, -32'sd170680, -32'sd1017181, -32'sd1325177, -32'sd1119196, -32'sd673327, -32'sd315641, -32'sd3555528, -32'sd3576434, 32'sd549376, 32'sd1924674, 32'sd5430788, 32'sd3010709, -32'sd167668, -32'sd1314416, -32'sd912834, -32'sd1705114, 32'sd2659565, -32'sd5313126, -32'sd2937359, 32'sd24256, -32'sd285218, 32'sd71813, 32'sd737405, -32'sd1144215, 32'sd2998249, 32'sd1763530, -32'sd273300, -32'sd1009277, -32'sd2078048, -32'sd3556768, -32'sd945087, 32'sd659343, 32'sd1235202, 32'sd3735769, -32'sd839839, 32'sd2148089, 32'sd3244756, 32'sd3864246, 32'sd3948448, 32'sd3584611, -32'sd484913, -32'sd3028679, -32'sd3677531, -32'sd2973151, -32'sd3528039, -32'sd6954350, 32'sd1267403, -32'sd2433836, 32'sd2386392, 32'sd971261, 32'sd3034782, 32'sd2021975, 32'sd2011296, -32'sd1083957, 32'sd97594, -32'sd1696128, 32'sd1020978, 32'sd599416, -32'sd2198857, -32'sd1261352, 32'sd1610600, 32'sd3748998, 32'sd736750, 32'sd1053441, 32'sd3006083, 32'sd6237450, 32'sd1909542, 32'sd554514, -32'sd5304725, -32'sd3723638, -32'sd3629711, -32'sd4215964, -32'sd5878571, -32'sd3267531, 32'sd35607, -32'sd305316, 32'sd3140511, -32'sd5205754, 32'sd595975, 32'sd2212754, -32'sd1207163, 32'sd880123, 32'sd497025, 32'sd1869747, -32'sd83817, 32'sd1771066, 32'sd280527, -32'sd723033, 32'sd1507820, 32'sd766796, -32'sd3180675, -32'sd3922315, 32'sd2251543, 32'sd1108095, -32'sd117936, -32'sd944692, -32'sd3059278, -32'sd223389, -32'sd1093476, -32'sd1611536, -32'sd3218097, -32'sd1531529, 32'sd1967108, 32'sd673790, -32'sd2216750, -32'sd3520421, 32'sd906517, 32'sd1343062, 32'sd65319, -32'sd363862, 32'sd1408146, -32'sd697639, -32'sd778974, -32'sd374320, 32'sd539820, 32'sd1724583, -32'sd515311, -32'sd1722970, -32'sd1141650, -32'sd575487, -32'sd700678, 32'sd2595743, 32'sd2928477, 32'sd1349290, 32'sd3303216, 32'sd2397742, 32'sd1484034, 32'sd624352, 32'sd490630, -32'sd1875686, 32'sd2302176, -32'sd3474561, -32'sd4421504, -32'sd3741756, -32'sd2869896, 32'sd755723, 32'sd910003, -32'sd50740, -32'sd821411, 32'sd523885, 32'sd232900, 32'sd16422, 32'sd3648417, 32'sd599464, -32'sd1259357, -32'sd715194, 32'sd1018912, 32'sd33861, 32'sd3227897, 32'sd1781253, 32'sd4544417, 32'sd685908, 32'sd3645110, 32'sd2370216, 32'sd3987010, 32'sd1859556, 32'sd1246468, -32'sd2601334, 32'sd927511, -32'sd1530798, -32'sd5213678, -32'sd5012792, -32'sd3532726, 32'sd32143, 32'sd2008887, -32'sd36180, -32'sd462208, 32'sd594055, 32'sd2320491, 32'sd675663, -32'sd242812, -32'sd2186800, -32'sd2911985, 32'sd430393, 32'sd720114, -32'sd1157063, 32'sd3571324, 32'sd2951293, 32'sd3972208, 32'sd4694927, 32'sd5417173, 32'sd2020278, 32'sd4711952, 32'sd4482344, -32'sd379909, 32'sd1418626, -32'sd1096476, -32'sd5416546, -32'sd5680284, 32'sd0, 32'sd543245, -32'sd9771, -32'sd1182577, 32'sd4203518, 32'sd1843766, -32'sd280614, 32'sd381999, -32'sd2008644, -32'sd2952197, -32'sd5175966, -32'sd3044069, -32'sd2633684, -32'sd1248477, 32'sd1582438, 32'sd2422386, 32'sd2391054, 32'sd4243140, 32'sd3537174, -32'sd809241, 32'sd1661891, 32'sd2774360, -32'sd1358868, -32'sd1412017, 32'sd914455, 32'sd560018, 32'sd1597209, -32'sd4754787, -32'sd1447208, -32'sd155113, 32'sd855540, -32'sd1050380, -32'sd576701, -32'sd527375, -32'sd2215752, -32'sd1735289, -32'sd650406, -32'sd92009, -32'sd2287158, -32'sd673976, -32'sd2384593, 32'sd109655, -32'sd695730, 32'sd724335, 32'sd1430980, 32'sd3189465, 32'sd960945, -32'sd1560513, 32'sd534191, 32'sd246763, -32'sd754995, -32'sd2831803, -32'sd3495213, -32'sd3588400, -32'sd790598, -32'sd1121158, 32'sd1178182, 32'sd161599, -32'sd957892, 32'sd2951046, 32'sd465967, 32'sd115628, -32'sd1878907, -32'sd572026, -32'sd466529, 32'sd1808864, -32'sd4074864, -32'sd3573019, -32'sd6600145, -32'sd3356909, -32'sd1365378, 32'sd174532, 32'sd1128097, 32'sd440115, -32'sd1083027, -32'sd846605, -32'sd1942848, -32'sd2286058, -32'sd4552590, -32'sd4589403, -32'sd1404685, -32'sd3271088, -32'sd4501727, -32'sd20598, 32'sd0, -32'sd1624836, -32'sd123891, -32'sd63384, -32'sd4393919, -32'sd4098191, -32'sd1478403, -32'sd1046633, 32'sd274593, -32'sd446134, 32'sd862364, -32'sd1765477, -32'sd2786532, -32'sd2423666, -32'sd2673388, -32'sd919240, 32'sd1142984, 32'sd668819, -32'sd545727, -32'sd1066394, -32'sd2277164, -32'sd2017952, -32'sd650771, -32'sd1077963, -32'sd1295736, -32'sd2419600, -32'sd3252507, -32'sd4296770, 32'sd623035, -32'sd1411569, -32'sd548339, -32'sd2912772, -32'sd1886090, 32'sd2072630, -32'sd6330, -32'sd1233263, 32'sd1265671, -32'sd2020995, -32'sd930445, -32'sd144473, -32'sd936369, 32'sd80431, -32'sd426886, 32'sd588421, -32'sd2023809, 32'sd1338550, 32'sd154576, 32'sd1151198, -32'sd664968, -32'sd2860845, 32'sd598486, -32'sd1954563, 32'sd1034553, 32'sd1759959, -32'sd2284196, -32'sd3924422, 32'sd973313, 32'sd335529, -32'sd1011355, 32'sd279194, 32'sd1291866, 32'sd2327495, 32'sd326319, -32'sd1498733, -32'sd903323, -32'sd265182, -32'sd649733, -32'sd569620, -32'sd2370045, -32'sd1834849, -32'sd244529, 32'sd1092279, 32'sd960386, -32'sd290799, -32'sd1664238, 32'sd2615514, 32'sd78153, -32'sd487158, 32'sd1564230, -32'sd2223512, 32'sd79548, 32'sd633876, -32'sd954351, -32'sd5170423, 32'sd0, -32'sd5364334, -32'sd1064447, 32'sd2242643, -32'sd416948, -32'sd2444266, -32'sd406097, 32'sd1507695, -32'sd1749826, 32'sd1195616, 32'sd30942, 32'sd319411, -32'sd2074023, 32'sd428022, 32'sd1060676, 32'sd1887439, -32'sd1641135, -32'sd539404, 32'sd98606, 32'sd256727, 32'sd402819, 32'sd1404777, -32'sd1171272, -32'sd1930260, 32'sd50675, -32'sd2129153, 32'sd2438147, 32'sd0, 32'sd0, 32'sd0, -32'sd4714345, 32'sd307179, 32'sd392963, -32'sd2107472, 32'sd187348, 32'sd1872568, -32'sd337744, 32'sd1267028, -32'sd909465, 32'sd1020221, -32'sd685928, -32'sd995055, -32'sd1500665, -32'sd1332139, -32'sd910722, -32'sd2707002, -32'sd1660325, -32'sd248378, 32'sd2133446, -32'sd177218, -32'sd476586, 32'sd560559, 32'sd557873, 32'sd814598, -32'sd5195922, 32'sd0, 32'sd0, 32'sd0, -32'sd4755914, -32'sd689019, -32'sd87134, 32'sd1534890, 32'sd621395, 32'sd1021330, -32'sd79456, 32'sd1240345, -32'sd949024, 32'sd1747212, 32'sd536903, -32'sd931987, -32'sd16426, -32'sd1923022, -32'sd1652244, 32'sd357253, -32'sd879712, -32'sd2799999, -32'sd620118, -32'sd638579, 32'sd934476, 32'sd239151, 32'sd65660, -32'sd4633008, -32'sd3762966, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3101647, -32'sd619949, -32'sd1948076, -32'sd775054, -32'sd31627, 32'sd1388198, 32'sd191014, 32'sd1107077, -32'sd817358, 32'sd458634, -32'sd1102253, -32'sd1095177, -32'sd1164059, -32'sd856093, 32'sd671085, -32'sd2136319, -32'sd458331, -32'sd12472, 32'sd10746, 32'sd602578, -32'sd2162433, -32'sd3387243, -32'sd5325794, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4937287, -32'sd5728673, -32'sd2466381, 32'sd912870, -32'sd1406931, 32'sd911623, -32'sd783972, 32'sd1559273, -32'sd1437407, 32'sd348620, 32'sd821115, -32'sd1893877, -32'sd956332, 32'sd1407046, 32'sd187719, 32'sd1442602, 32'sd717252, -32'sd870191, -32'sd1800982, -32'sd4926071, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd44561, 32'sd17722, -32'sd3380779, -32'sd5147527, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4351056, -32'sd5384585, -32'sd5094546, -32'sd6008236, -32'sd5103756, -32'sd2863413, -32'sd408673, -32'sd1363210, -32'sd1958815, -32'sd3616103, 32'sd901700, 32'sd982478, -32'sd334834, -32'sd1735083, -32'sd5836126, -32'sd3707126, -32'sd4149538, -32'sd4304045, -32'sd3494167, -32'sd3863081, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4552220, -32'sd2099508, 32'sd295966, -32'sd1123156, 32'sd1470437, 32'sd645681, -32'sd1163643, -32'sd822855, -32'sd2602252, -32'sd2802905, -32'sd1576453, -32'sd3069135, -32'sd3847421, -32'sd980244, 32'sd268902, -32'sd2485624, -32'sd1817480, 32'sd1093648, -32'sd409058, -32'sd1412549, 32'sd1609956, -32'sd1674351, -32'sd6048867, -32'sd5646961, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4484926, 32'sd379007, -32'sd1996679, -32'sd1547748, 32'sd1133997, -32'sd2289307, -32'sd4702218, -32'sd2517900, -32'sd940150, -32'sd4124766, -32'sd3249093, -32'sd7849034, -32'sd6506905, -32'sd6454163, -32'sd4633266, -32'sd2682556, -32'sd2105209, -32'sd1512311, -32'sd89564, -32'sd434641, 32'sd3093232, -32'sd1173144, 32'sd455342, -32'sd1615100, -32'sd4118510, 32'sd0, 32'sd0, -32'sd3774270, -32'sd699502, 32'sd199544, -32'sd3360254, -32'sd1160868, -32'sd752144, 32'sd1331613, -32'sd2806953, -32'sd2373898, -32'sd2805721, -32'sd5566169, -32'sd6079996, -32'sd3394842, -32'sd5656777, -32'sd5120118, -32'sd5753533, -32'sd5009197, -32'sd3296741, -32'sd4101425, -32'sd3428044, -32'sd1663695, -32'sd232296, -32'sd391720, 32'sd1230227, -32'sd994459, 32'sd865708, -32'sd5047762, 32'sd0, -32'sd4333936, 32'sd191601, -32'sd1095679, -32'sd1708352, -32'sd2336461, -32'sd2732368, -32'sd1643389, 32'sd1946246, -32'sd1306460, -32'sd91926, -32'sd1108667, -32'sd1410221, -32'sd1195967, -32'sd649666, -32'sd3588109, -32'sd4317323, -32'sd3019192, -32'sd5243920, -32'sd5516853, -32'sd2687776, -32'sd4319722, -32'sd2364072, -32'sd749502, 32'sd1577934, 32'sd1162599, -32'sd420985, -32'sd4890634, 32'sd0, 32'sd716794, -32'sd1790834, 32'sd777193, 32'sd3764394, -32'sd845236, -32'sd2016463, -32'sd279325, 32'sd1037559, -32'sd326737, 32'sd943158, 32'sd652446, 32'sd2117306, 32'sd689927, 32'sd2530872, 32'sd912479, 32'sd1214854, 32'sd2582239, -32'sd74928, 32'sd2082547, 32'sd1025862, 32'sd1215993, 32'sd2701304, 32'sd1451825, 32'sd2333914, 32'sd50765, 32'sd2003531, -32'sd357165, -32'sd3795256, -32'sd1688750, -32'sd1110893, 32'sd2547110, 32'sd1948474, -32'sd1339212, 32'sd360092, -32'sd1521246, -32'sd2313226, -32'sd6407, 32'sd2326625, 32'sd1443681, 32'sd3324050, 32'sd3884717, 32'sd1542060, 32'sd1119335, 32'sd3042713, 32'sd3513693, 32'sd1925066, 32'sd2451965, 32'sd2732017, 32'sd4354500, 32'sd916359, 32'sd2845398, -32'sd647816, 32'sd576248, 32'sd243535, -32'sd87770, -32'sd1195465, 32'sd2283930, -32'sd2583408, -32'sd2617231, 32'sd144440, -32'sd940884, -32'sd272682, -32'sd1419673, -32'sd619829, 32'sd1232797, -32'sd701316, 32'sd1198585, 32'sd309807, -32'sd1331220, 32'sd647615, 32'sd1454241, 32'sd1553195, 32'sd1158646, 32'sd1669624, 32'sd1325715, 32'sd497219, 32'sd2637660, -32'sd1092446, -32'sd1667602, 32'sd1890262, 32'sd3164956, 32'sd2421770, -32'sd3913557, -32'sd5371891, -32'sd4996454, -32'sd2938687, -32'sd505715, 32'sd1119964, -32'sd454469, 32'sd2894305, 32'sd1238757, -32'sd970493, 32'sd948780, 32'sd804681, 32'sd499187, 32'sd1350695, 32'sd190649, -32'sd1099765, -32'sd1320719, -32'sd654895, 32'sd2813129, 32'sd3015101, 32'sd776907, 32'sd60784, -32'sd1356357, -32'sd2098487, -32'sd2848880, -32'sd2246719, -32'sd1073712, 32'sd2033389, -32'sd5576363, -32'sd5136248, -32'sd5923312, -32'sd6358159, -32'sd948262, -32'sd795006, 32'sd1446536, 32'sd1227101, 32'sd308762, -32'sd1320222, -32'sd119966, 32'sd1489600, 32'sd791611, 32'sd1908314, -32'sd668917, -32'sd4286459, -32'sd394438, -32'sd957898, -32'sd266950, 32'sd1446687, 32'sd2650391, -32'sd613725, 32'sd984638, -32'sd1444289, -32'sd3140602, -32'sd396924, 32'sd3804938, 32'sd998762, -32'sd5561662, -32'sd5777893, -32'sd7311151, 32'sd1922106, -32'sd215068, -32'sd920225, -32'sd2258, -32'sd137467, -32'sd913512, 32'sd1880615, 32'sd326854, 32'sd951076, 32'sd2452187, 32'sd2635133, -32'sd1804650, -32'sd1037879, -32'sd653408, -32'sd416209, 32'sd2539985, 32'sd3544778, -32'sd1124179, 32'sd276414, 32'sd80887, -32'sd761160, 32'sd710366, -32'sd1697036, 32'sd1118684, -32'sd77932, -32'sd5586395, -32'sd4671448, -32'sd5385719, 32'sd1179519, -32'sd1411529, -32'sd101567, -32'sd1703337, 32'sd3211286, 32'sd87540, 32'sd2654286, 32'sd688839, 32'sd3857441, 32'sd326985, -32'sd2294591, -32'sd1889130, -32'sd2531912, -32'sd33834, 32'sd2613798, 32'sd155661, 32'sd1343177, 32'sd1216739, -32'sd967357, -32'sd144421, 32'sd419813, -32'sd251083, -32'sd2783485, -32'sd3704473, -32'sd4219510, -32'sd3300020, -32'sd3355021, -32'sd5045371, 32'sd773432, -32'sd1861834, 32'sd309066, -32'sd806409, 32'sd723087, 32'sd2661228, 32'sd2892614, 32'sd1006959, 32'sd2600047, -32'sd74333, -32'sd551182, 32'sd376638, 32'sd2005754, 32'sd858844, 32'sd2460565, 32'sd2950046, -32'sd1314850, 32'sd866176, 32'sd571766, 32'sd340362, 32'sd995612, -32'sd3217281, -32'sd2989942, -32'sd2496702, -32'sd4173754, -32'sd3870338, -32'sd4776246, -32'sd3222185, -32'sd368657, 32'sd901907, 32'sd1024973, -32'sd481988, 32'sd1760370, 32'sd2433157, 32'sd2428123, 32'sd2655671, 32'sd1779918, -32'sd325894, 32'sd154127, 32'sd149753, -32'sd523882, 32'sd1509102, 32'sd1745243, 32'sd446085, 32'sd196487, -32'sd1486041, -32'sd588634, -32'sd53677, -32'sd76691, -32'sd2773481, -32'sd4002236, -32'sd3990568, -32'sd4607240, -32'sd3573077, -32'sd3988616, -32'sd5339730, -32'sd3785877, 32'sd688751, 32'sd2407402, 32'sd141155, 32'sd478026, 32'sd2449725, 32'sd3376931, 32'sd2081522, 32'sd3135712, 32'sd1920225, 32'sd194972, -32'sd1169680, -32'sd3404742, 32'sd2697873, 32'sd1690713, 32'sd2310322, 32'sd1397144, 32'sd341440, 32'sd1157555, -32'sd344631, 32'sd966460, -32'sd10945, -32'sd1685833, -32'sd5086579, -32'sd4524678, -32'sd5302181, -32'sd4334641, -32'sd4453508, -32'sd629418, 32'sd394170, 32'sd242629, 32'sd2282912, -32'sd134742, 32'sd2608529, 32'sd2496468, -32'sd26380, 32'sd912677, 32'sd1050507, -32'sd1009980, -32'sd3182533, -32'sd3888775, 32'sd254789, 32'sd292400, 32'sd835927, 32'sd627212, -32'sd424237, -32'sd1384095, -32'sd2418080, -32'sd427210, -32'sd289653, -32'sd900741, -32'sd1582214, 32'sd83283, -32'sd781519, 32'sd0, -32'sd4232121, -32'sd999460, 32'sd734611, 32'sd259047, 32'sd2187522, 32'sd1752168, 32'sd2024296, 32'sd3455062, 32'sd944605, 32'sd2934193, -32'sd156381, -32'sd1013921, -32'sd1130504, -32'sd5271523, 32'sd395320, 32'sd386811, -32'sd42194, -32'sd298734, 32'sd135448, -32'sd664850, 32'sd821313, 32'sd1374550, -32'sd376396, -32'sd924428, 32'sd1096372, 32'sd2121331, -32'sd457193, -32'sd3911401, -32'sd5777103, -32'sd793583, 32'sd1863476, -32'sd126790, 32'sd534485, 32'sd1581910, 32'sd2029510, -32'sd252869, 32'sd1463297, 32'sd1987268, 32'sd1013499, -32'sd2351231, -32'sd2082386, -32'sd2395561, -32'sd1551183, 32'sd177455, 32'sd665199, -32'sd1729425, -32'sd567427, -32'sd213948, -32'sd634979, -32'sd1060409, -32'sd1781019, -32'sd3466168, -32'sd2679827, 32'sd4091205, -32'sd3062330, -32'sd5461405, -32'sd5668243, 32'sd535222, -32'sd1135265, -32'sd18512, 32'sd425618, -32'sd3941817, -32'sd2583058, -32'sd1431685, -32'sd2854949, -32'sd2334688, -32'sd1424453, -32'sd2445444, -32'sd3627144, -32'sd219750, -32'sd982043, 32'sd764359, -32'sd1757797, -32'sd2484331, 32'sd170578, -32'sd1271550, -32'sd2187128, -32'sd3044562, -32'sd2865333, -32'sd3194257, -32'sd271599, -32'sd2844296, -32'sd3605304, 32'sd0, -32'sd3834470, 32'sd1797297, 32'sd126476, -32'sd1763011, -32'sd2759769, -32'sd6841641, -32'sd7304139, -32'sd5062684, -32'sd3432694, -32'sd5007042, -32'sd2804203, -32'sd6101080, -32'sd3888613, -32'sd3046041, -32'sd2349652, 32'sd224673, -32'sd710500, -32'sd150163, 32'sd812120, -32'sd2401538, -32'sd557824, -32'sd2343718, -32'sd2064809, -32'sd1563767, 32'sd3488723, -32'sd4312053, -32'sd4564173, -32'sd854330, -32'sd2517717, -32'sd3584616, -32'sd2473587, -32'sd3486079, -32'sd2055079, -32'sd4253904, -32'sd6497294, -32'sd4266197, -32'sd1792680, -32'sd2211732, -32'sd2744000, -32'sd1266152, -32'sd2563645, -32'sd4675583, -32'sd3043046, -32'sd885893, -32'sd3567374, -32'sd720278, -32'sd2308604, -32'sd722310, -32'sd1058065, 32'sd32035, -32'sd758047, 32'sd758066, -32'sd355918, -32'sd3013023, 32'sd505141, 32'sd1289170, 32'sd829717, -32'sd2105102, -32'sd541069, -32'sd3685803, -32'sd1551198, 32'sd830596, -32'sd1452636, 32'sd1149366, -32'sd1475517, -32'sd1519715, -32'sd3387880, -32'sd949021, -32'sd2679955, -32'sd255761, -32'sd3724466, -32'sd1933179, -32'sd903471, -32'sd1166775, -32'sd2652276, -32'sd729896, -32'sd2106170, 32'sd927882, -32'sd163, -32'sd6276, 32'sd1500396, -32'sd2856342, 32'sd15743, 32'sd0, -32'sd4727308, -32'sd695882, -32'sd200106, -32'sd1644057, 32'sd1757827, 32'sd2698062, 32'sd149504, 32'sd334338, -32'sd1755733, 32'sd673668, 32'sd154493, -32'sd2564754, -32'sd1322775, -32'sd1048586, -32'sd3903161, -32'sd820719, -32'sd1760106, -32'sd620456, -32'sd393136, 32'sd622514, 32'sd1417237, 32'sd18010, 32'sd412588, -32'sd802022, -32'sd782411, -32'sd893523, 32'sd0, 32'sd0, 32'sd0, -32'sd2673054, -32'sd413663, 32'sd1018217, 32'sd1560380, 32'sd423754, 32'sd864657, 32'sd2465602, 32'sd127234, -32'sd494286, -32'sd1498407, -32'sd1656448, -32'sd199901, -32'sd3897668, -32'sd2607166, 32'sd366177, -32'sd461686, -32'sd10305, -32'sd1579697, 32'sd1894564, 32'sd823165, -32'sd325155, 32'sd3115263, 32'sd680788, -32'sd2609866, -32'sd3442457, 32'sd0, 32'sd0, 32'sd0, -32'sd4660712, 32'sd774369, 32'sd1452281, 32'sd348047, -32'sd2443890, 32'sd434464, -32'sd1515472, -32'sd2672907, 32'sd44047, 32'sd118970, -32'sd1283968, 32'sd415114, 32'sd436639, -32'sd122915, 32'sd1052439, 32'sd853610, -32'sd1600064, -32'sd995319, 32'sd1465883, 32'sd2480596, 32'sd1211567, 32'sd1417973, 32'sd56928, 32'sd746473, -32'sd5503877, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4399161, -32'sd2933129, -32'sd1714299, -32'sd367049, 32'sd1546393, 32'sd1878450, 32'sd605541, -32'sd1903486, 32'sd2041701, 32'sd695735, 32'sd2276814, 32'sd2976177, 32'sd1204507, 32'sd976219, 32'sd2444945, 32'sd1638310, 32'sd1036516, 32'sd1951291, 32'sd78067, -32'sd1375936, -32'sd1407292, -32'sd3569642, -32'sd4757499, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4868219, -32'sd5051025, -32'sd5171429, -32'sd5025620, -32'sd4035137, -32'sd1716117, 32'sd115463, 32'sd734756, 32'sd1399879, 32'sd2351107, -32'sd897361, -32'sd235952, 32'sd306149, 32'sd1415122, 32'sd173036, -32'sd291, -32'sd1171768, -32'sd1866054, 32'sd139930, -32'sd5445968, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2093317, -32'sd1727481, 32'sd111006, -32'sd41510, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd119545, -32'sd875086, 32'sd1221729, 32'sd1817994, -32'sd957222, -32'sd3453111, 32'sd1102847, 32'sd915877, 32'sd749291, 32'sd1091009, -32'sd284063, 32'sd2033121, 32'sd890076, -32'sd327831, 32'sd1761139, 32'sd2073733, 32'sd2826394, 32'sd2118912, 32'sd742679, 32'sd833749, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd100449, -32'sd1321548, -32'sd54366, -32'sd2505568, -32'sd1425863, 32'sd1189015, 32'sd1477363, -32'sd627051, -32'sd1458576, 32'sd247720, -32'sd1615047, -32'sd1297892, -32'sd2037501, -32'sd732776, 32'sd312188, -32'sd451739, 32'sd61234, 32'sd729199, -32'sd342694, 32'sd987585, 32'sd2020237, 32'sd1959424, 32'sd1401589, 32'sd1472882, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1177044, 32'sd2011005, 32'sd865871, 32'sd562353, 32'sd75570, 32'sd1458832, 32'sd1819258, -32'sd1321207, -32'sd1655944, -32'sd1522989, -32'sd1679826, -32'sd879732, -32'sd2524324, 32'sd314062, -32'sd2005458, 32'sd1167613, 32'sd1115826, 32'sd1472374, 32'sd1168530, 32'sd1511731, 32'sd838970, -32'sd397583, 32'sd930638, 32'sd409154, 32'sd735723, 32'sd0, 32'sd0, -32'sd139189, 32'sd1436788, -32'sd134923, -32'sd1133889, 32'sd69454, -32'sd2443470, -32'sd2711786, -32'sd4276639, -32'sd1597729, -32'sd2667517, -32'sd793664, 32'sd18795, -32'sd584822, -32'sd1005722, -32'sd1113237, 32'sd1157305, 32'sd1147842, 32'sd2044815, 32'sd2094304, -32'sd598529, 32'sd1773076, 32'sd393655, 32'sd1093024, 32'sd323084, 32'sd978300, 32'sd266404, -32'sd1042425, 32'sd0, 32'sd803240, 32'sd828501, 32'sd686163, -32'sd1678848, 32'sd1378111, 32'sd409620, -32'sd2355990, -32'sd1359089, 32'sd398212, -32'sd677398, -32'sd2083904, -32'sd2486279, -32'sd2223012, -32'sd1196105, -32'sd655658, 32'sd399916, 32'sd1406961, 32'sd1045489, 32'sd1042635, 32'sd1352004, 32'sd1919879, 32'sd2459878, 32'sd3169112, 32'sd2585491, 32'sd322016, 32'sd745097, -32'sd925993, 32'sd0, 32'sd447124, 32'sd32201, 32'sd55094, -32'sd2408033, 32'sd663901, -32'sd3472607, -32'sd285680, 32'sd1104809, -32'sd876824, -32'sd246791, 32'sd103140, -32'sd748103, -32'sd2380418, -32'sd2055115, -32'sd1244204, 32'sd279340, 32'sd847556, 32'sd1511305, 32'sd1253297, 32'sd650229, -32'sd436582, -32'sd557098, 32'sd264614, 32'sd3606230, 32'sd2374251, 32'sd829785, 32'sd1505402, 32'sd2274627, 32'sd850672, 32'sd474183, 32'sd1649921, -32'sd2923832, -32'sd900341, -32'sd646355, 32'sd293736, -32'sd1662850, -32'sd806925, -32'sd1463347, -32'sd2056562, -32'sd1522045, -32'sd2794972, 32'sd198325, 32'sd1658403, 32'sd740008, 32'sd289834, -32'sd457046, -32'sd596783, 32'sd1595297, 32'sd600854, 32'sd3179656, -32'sd471165, -32'sd391660, 32'sd160703, 32'sd2747733, -32'sd593969, 32'sd1271752, 32'sd181140, -32'sd2052775, 32'sd383381, 32'sd1190646, 32'sd1060382, -32'sd1125109, -32'sd1300540, -32'sd2484565, -32'sd2720578, -32'sd581078, -32'sd449040, 32'sd1691970, -32'sd237992, -32'sd921163, -32'sd1654485, -32'sd1584846, 32'sd1600953, 32'sd777038, 32'sd3703961, 32'sd2203749, 32'sd3427672, 32'sd3065457, 32'sd2216120, 32'sd4364529, 32'sd684702, 32'sd1995400, 32'sd838797, 32'sd311929, 32'sd788033, -32'sd2886449, 32'sd668574, -32'sd1003161, -32'sd4288446, -32'sd2560853, -32'sd1304773, -32'sd149557, 32'sd162328, 32'sd159500, 32'sd17203, -32'sd474424, 32'sd12593, -32'sd1825413, -32'sd231935, -32'sd2720022, -32'sd1482223, -32'sd3429261, -32'sd4000646, -32'sd3599744, -32'sd2434445, 32'sd511925, 32'sd1555570, 32'sd1429833, 32'sd1186260, -32'sd1073453, 32'sd134624, -32'sd311813, 32'sd1138357, -32'sd1683241, -32'sd1041591, -32'sd1120192, -32'sd2724563, -32'sd2412815, -32'sd1871817, -32'sd1132575, 32'sd613721, 32'sd1372586, 32'sd2065663, 32'sd697822, 32'sd3214798, 32'sd1961439, -32'sd756475, -32'sd1555792, -32'sd1588569, -32'sd1112999, -32'sd3163745, -32'sd9000535, -32'sd9924936, -32'sd10014435, -32'sd6156526, -32'sd2386443, -32'sd641147, 32'sd2233102, 32'sd1804353, -32'sd120735, -32'sd785520, -32'sd1224995, 32'sd1338002, -32'sd1159047, -32'sd70951, -32'sd22266, 32'sd1277128, -32'sd3401987, -32'sd3418616, -32'sd2373955, 32'sd1381547, 32'sd2023008, 32'sd1622194, 32'sd3182052, 32'sd767491, 32'sd696000, 32'sd242862, -32'sd1471277, -32'sd2473666, -32'sd8472475, -32'sd10790364, -32'sd11157768, -32'sd7230775, -32'sd4408524, 32'sd1584945, -32'sd235840, 32'sd1262732, 32'sd1471301, 32'sd121587, -32'sd642068, 32'sd2179254, -32'sd428824, -32'sd2664583, -32'sd843446, -32'sd429586, -32'sd2652765, -32'sd2778484, 32'sd204416, 32'sd418627, 32'sd132467, 32'sd3544003, 32'sd3199525, -32'sd404337, -32'sd1487858, -32'sd272050, -32'sd2397785, -32'sd2356824, -32'sd3957096, -32'sd3357192, -32'sd1759675, -32'sd2733726, -32'sd4280804, -32'sd2289756, 32'sd213327, -32'sd1478182, 32'sd846371, 32'sd1083619, -32'sd498441, 32'sd921894, -32'sd1996432, -32'sd526192, -32'sd1253794, 32'sd263989, -32'sd250180, -32'sd1635400, -32'sd166430, -32'sd154834, -32'sd1386838, 32'sd1682050, 32'sd2084850, 32'sd2031866, 32'sd708516, 32'sd922147, -32'sd1316979, 32'sd214830, 32'sd623081, 32'sd1038039, -32'sd480192, 32'sd1178696, -32'sd4421094, -32'sd2554996, -32'sd1587948, 32'sd155903, 32'sd40751, 32'sd100725, -32'sd1567105, 32'sd975260, 32'sd1115442, 32'sd282962, 32'sd152298, 32'sd997968, -32'sd2047965, 32'sd1803313, 32'sd1036710, -32'sd1214882, -32'sd1892049, 32'sd470102, 32'sd780902, -32'sd655581, 32'sd1751321, -32'sd549042, -32'sd918433, -32'sd631120, 32'sd1142779, 32'sd2505426, -32'sd1188663, -32'sd1036114, 32'sd518199, -32'sd2504107, -32'sd25412, -32'sd705993, 32'sd715352, -32'sd259026, 32'sd1163728, 32'sd1203762, -32'sd2254672, -32'sd389237, -32'sd675447, -32'sd1599367, -32'sd941548, 32'sd250496, -32'sd2183401, -32'sd2083613, 32'sd1108547, 32'sd1210336, -32'sd272968, -32'sd1614037, 32'sd2262906, -32'sd2442401, 32'sd709609, -32'sd12560, 32'sd3762430, 32'sd1931424, -32'sd595836, 32'sd158853, -32'sd744118, 32'sd343547, -32'sd598812, 32'sd260572, -32'sd733891, 32'sd1565157, -32'sd144990, -32'sd187528, -32'sd1225221, -32'sd1742804, -32'sd763712, -32'sd1420366, 32'sd255073, -32'sd3154698, -32'sd501265, -32'sd148603, -32'sd917293, 32'sd714640, 32'sd535880, 32'sd1694728, 32'sd463961, -32'sd3739870, 32'sd676818, 32'sd762981, 32'sd2875290, 32'sd1682021, -32'sd1984035, -32'sd2300017, 32'sd1196578, -32'sd1303950, -32'sd1394767, -32'sd2020088, 32'sd0, 32'sd1691187, -32'sd781177, -32'sd1428804, 32'sd1795933, 32'sd294052, -32'sd495660, 32'sd2116119, 32'sd552086, -32'sd1640161, 32'sd642440, -32'sd1073238, -32'sd1920306, -32'sd3648767, -32'sd1979013, -32'sd979256, -32'sd254215, -32'sd238796, 32'sd1557336, 32'sd1115541, 32'sd3595175, 32'sd962949, -32'sd1661899, -32'sd426143, 32'sd312004, -32'sd2048443, 32'sd1329942, -32'sd587980, -32'sd383890, -32'sd502805, 32'sd1036868, 32'sd43273, 32'sd1694224, 32'sd1927156, -32'sd80666, 32'sd558647, -32'sd769220, -32'sd894737, -32'sd494326, -32'sd2021908, -32'sd2173243, -32'sd1825319, -32'sd1066097, -32'sd1026157, -32'sd327803, 32'sd2273517, 32'sd3505493, 32'sd2875718, 32'sd2341412, 32'sd661090, -32'sd2193548, -32'sd1687455, -32'sd3420120, -32'sd2494230, 32'sd1254573, -32'sd715151, -32'sd95391, -32'sd151764, 32'sd1031858, 32'sd756743, -32'sd97780, 32'sd1062022, 32'sd1038966, -32'sd1715378, -32'sd105633, -32'sd588095, -32'sd169849, -32'sd1794808, -32'sd2026633, 32'sd414941, -32'sd154055, 32'sd1167315, 32'sd3714553, 32'sd693040, 32'sd3113470, 32'sd879627, 32'sd1684211, -32'sd362900, -32'sd1346854, -32'sd381587, -32'sd333254, -32'sd760378, 32'sd532595, -32'sd351229, 32'sd0, -32'sd764201, 32'sd654707, 32'sd998891, 32'sd1911329, -32'sd348910, 32'sd525120, -32'sd1523772, 32'sd2730901, 32'sd538666, -32'sd1241852, 32'sd237887, -32'sd1427662, 32'sd313184, 32'sd1951395, 32'sd1916882, 32'sd2359972, 32'sd588779, -32'sd31623, 32'sd1298075, -32'sd110665, 32'sd1616027, 32'sd738474, 32'sd513289, 32'sd1255186, -32'sd550275, 32'sd982928, -32'sd1349202, -32'sd502608, 32'sd90932, -32'sd951796, -32'sd474977, 32'sd58665, -32'sd1476460, 32'sd1186018, -32'sd110109, -32'sd226877, -32'sd533343, 32'sd950446, 32'sd1282913, 32'sd3401170, 32'sd826221, 32'sd2157466, 32'sd2721788, 32'sd656450, 32'sd336965, 32'sd1984161, -32'sd947029, 32'sd2019521, -32'sd1130151, -32'sd4543682, 32'sd1462378, 32'sd1584736, -32'sd964659, 32'sd301410, 32'sd454722, 32'sd1557878, 32'sd533831, 32'sd1552450, -32'sd2384801, 32'sd773963, -32'sd449216, -32'sd2988427, -32'sd993672, -32'sd474593, -32'sd677148, 32'sd637912, 32'sd1220237, 32'sd1815564, -32'sd376856, -32'sd1715078, 32'sd4786880, 32'sd2538480, 32'sd874874, 32'sd10114, 32'sd530230, -32'sd1179434, -32'sd3710973, -32'sd3065784, 32'sd992863, 32'sd194065, -32'sd1898661, 32'sd796665, 32'sd238329, 32'sd0, -32'sd522354, 32'sd269222, -32'sd1409062, 32'sd408045, 32'sd3175259, 32'sd1548220, -32'sd1090981, -32'sd186481, 32'sd1487278, 32'sd65880, 32'sd124374, 32'sd1888866, -32'sd473424, 32'sd690028, 32'sd2263669, -32'sd1813750, 32'sd595018, -32'sd383718, -32'sd2153869, -32'sd392825, -32'sd474444, -32'sd1834626, -32'sd1049181, 32'sd828407, -32'sd561380, 32'sd937936, 32'sd0, 32'sd0, 32'sd0, -32'sd403887, 32'sd710035, 32'sd958633, -32'sd67159, 32'sd813351, -32'sd805772, 32'sd2780266, 32'sd3064563, 32'sd605762, -32'sd1647312, -32'sd758457, 32'sd137382, 32'sd1470340, -32'sd204036, -32'sd922734, 32'sd520650, 32'sd1565946, -32'sd1476985, -32'sd1241495, 32'sd992400, -32'sd1084452, 32'sd49112, 32'sd924174, 32'sd603579, -32'sd82064, 32'sd0, 32'sd0, 32'sd0, 32'sd190819, 32'sd1127484, 32'sd983685, 32'sd605365, 32'sd3000771, 32'sd895814, 32'sd4437715, 32'sd2872388, 32'sd1172864, 32'sd1273102, 32'sd1201659, 32'sd2355075, 32'sd400157, -32'sd152918, -32'sd1336799, -32'sd2122870, 32'sd1677847, -32'sd920839, -32'sd1170160, 32'sd2140736, 32'sd1009600, 32'sd924300, 32'sd1147999, -32'sd1137874, -32'sd830397, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd55192, 32'sd245079, -32'sd2134263, -32'sd336192, -32'sd2222469, -32'sd1708649, 32'sd1033409, 32'sd2046832, 32'sd1066189, -32'sd248389, -32'sd1692059, -32'sd2727970, -32'sd409044, 32'sd1825086, 32'sd107523, -32'sd2939219, 32'sd793993, 32'sd2863195, 32'sd1612498, 32'sd436454, 32'sd481344, -32'sd114472, 32'sd420209, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd14971, 32'sd646207, -32'sd129685, 32'sd595409, 32'sd344462, -32'sd1563225, 32'sd1745941, 32'sd1780653, -32'sd1332520, -32'sd356101, 32'sd2611659, 32'sd3698199, 32'sd195513, 32'sd1000546, 32'sd785768, 32'sd1648645, 32'sd895397, -32'sd1978837, 32'sd31832, -32'sd301562, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2641294, -32'sd2982189, -32'sd878447, -32'sd1641406, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2778732, -32'sd1264444, -32'sd1699321, -32'sd206536, -32'sd2367413, -32'sd2412206, -32'sd2132659, -32'sd1796516, -32'sd2973198, -32'sd281761, -32'sd2667821, -32'sd2822646, -32'sd1573482, -32'sd2078314, -32'sd3273028, -32'sd1540345, -32'sd2321161, -32'sd1216914, -32'sd852978, -32'sd2589575, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2475921, -32'sd1016559, -32'sd3199755, -32'sd1932402, 32'sd1097576, 32'sd1608290, 32'sd659337, -32'sd1044923, -32'sd1689701, -32'sd1508363, -32'sd2080248, -32'sd1091438, -32'sd2552214, -32'sd5050417, -32'sd601301, -32'sd2693403, -32'sd1519049, 32'sd939728, 32'sd1620085, 32'sd967016, -32'sd2220368, -32'sd174615, -32'sd1950097, -32'sd2376457, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1866951, -32'sd420787, 32'sd1024986, 32'sd189301, -32'sd404532, -32'sd1515923, -32'sd2703829, -32'sd2588073, -32'sd268363, -32'sd2777696, -32'sd1369562, 32'sd637767, 32'sd730651, 32'sd647880, 32'sd2033047, 32'sd1296560, 32'sd1151443, 32'sd641856, 32'sd2026865, 32'sd689018, 32'sd633757, 32'sd794376, -32'sd46252, 32'sd675776, -32'sd1331871, 32'sd0, 32'sd0, -32'sd2283154, 32'sd575021, -32'sd84400, -32'sd1854986, -32'sd2568887, -32'sd2684990, 32'sd197476, -32'sd327987, -32'sd525446, -32'sd3108137, 32'sd210344, -32'sd2441142, 32'sd893431, 32'sd2484167, 32'sd2164570, 32'sd546610, 32'sd840141, 32'sd1964602, 32'sd2775285, -32'sd481924, -32'sd496495, 32'sd162979, -32'sd1018783, 32'sd43855, -32'sd2044530, 32'sd793621, -32'sd1524398, 32'sd0, 32'sd728730, 32'sd437841, -32'sd694566, -32'sd1049755, -32'sd1452174, -32'sd223371, -32'sd438973, 32'sd2107749, 32'sd3650309, 32'sd442665, -32'sd95171, 32'sd417823, -32'sd194685, 32'sd381411, 32'sd24514, 32'sd1571756, 32'sd1217163, 32'sd1482077, 32'sd1613366, -32'sd2338114, 32'sd960500, -32'sd930263, 32'sd85521, -32'sd826617, 32'sd1728553, -32'sd100574, -32'sd3297393, 32'sd0, -32'sd2703665, 32'sd714979, -32'sd1367955, -32'sd471397, 32'sd1881163, 32'sd1266357, -32'sd627921, 32'sd2346099, 32'sd13810, -32'sd277663, 32'sd324746, 32'sd2859634, 32'sd1531495, -32'sd1169771, -32'sd1392946, 32'sd204360, -32'sd754058, -32'sd436282, -32'sd248189, -32'sd1646743, 32'sd2668170, 32'sd1632710, -32'sd732614, -32'sd327816, 32'sd349675, -32'sd617871, -32'sd3393344, -32'sd2401811, 32'sd666831, -32'sd992608, 32'sd639809, 32'sd3594526, 32'sd114939, 32'sd1062924, 32'sd1093840, -32'sd266052, 32'sd2908891, 32'sd414862, 32'sd1756364, 32'sd2525192, 32'sd847022, -32'sd3598, 32'sd25515, -32'sd384266, 32'sd492913, 32'sd1797096, 32'sd847412, 32'sd903805, 32'sd1895599, 32'sd1668521, 32'sd2092747, 32'sd1365475, 32'sd2217365, -32'sd1426959, -32'sd2166066, 32'sd1707168, 32'sd80811, 32'sd792107, -32'sd31468, 32'sd1361043, 32'sd868622, -32'sd1656483, 32'sd830761, 32'sd1786657, 32'sd1722546, 32'sd879678, 32'sd187643, 32'sd2297464, -32'sd220742, 32'sd2587859, 32'sd2339439, 32'sd3526582, 32'sd1958011, 32'sd2219193, 32'sd676381, 32'sd3817339, 32'sd1854471, 32'sd2990627, 32'sd1749662, -32'sd628435, 32'sd598440, 32'sd2094445, -32'sd2852206, -32'sd3081932, -32'sd1357772, -32'sd1304211, -32'sd1003530, 32'sd399995, 32'sd919636, -32'sd596103, 32'sd1192402, -32'sd638190, 32'sd1442854, 32'sd1049019, -32'sd79381, 32'sd1805335, -32'sd826394, 32'sd2633606, 32'sd1255537, 32'sd1023344, 32'sd2012931, 32'sd4492862, 32'sd4040572, 32'sd2338091, 32'sd1359768, 32'sd771296, -32'sd341863, 32'sd2874712, 32'sd2262288, -32'sd158111, 32'sd974496, -32'sd2564162, -32'sd258611, 32'sd877242, -32'sd1287161, 32'sd688244, 32'sd1617312, 32'sd321315, 32'sd175948, -32'sd1081595, -32'sd807113, 32'sd1549284, 32'sd1281151, 32'sd1092542, 32'sd3161845, 32'sd1036279, 32'sd1794249, 32'sd1202787, 32'sd2347915, 32'sd3895504, 32'sd3087991, 32'sd3848752, 32'sd3055476, 32'sd198454, -32'sd628549, 32'sd466053, 32'sd381075, 32'sd868558, -32'sd219423, -32'sd761149, 32'sd1741767, 32'sd1316611, 32'sd2377237, -32'sd358064, -32'sd1756934, -32'sd859781, -32'sd282692, -32'sd10587, -32'sd375928, -32'sd928684, -32'sd60406, 32'sd2127800, -32'sd2410151, -32'sd6346027, -32'sd4439887, -32'sd1972547, -32'sd2099248, -32'sd429452, 32'sd139768, 32'sd822611, -32'sd273472, 32'sd1319072, -32'sd820573, -32'sd2928306, -32'sd60987, 32'sd1487009, -32'sd2579028, 32'sd370184, -32'sd443681, -32'sd430068, -32'sd1087432, 32'sd363739, -32'sd1158190, -32'sd977253, 32'sd808209, -32'sd885160, 32'sd53006, 32'sd478895, -32'sd1039127, 32'sd438652, -32'sd3728261, -32'sd8057640, -32'sd3533689, 32'sd57040, -32'sd1148138, -32'sd1726100, -32'sd4287308, -32'sd2120664, -32'sd2016068, 32'sd220787, -32'sd1665710, 32'sd2062968, -32'sd1707313, -32'sd1773264, -32'sd2803760, -32'sd2113899, 32'sd94173, 32'sd334948, 32'sd903719, -32'sd35825, -32'sd1410771, -32'sd45724, 32'sd120853, 32'sd1634131, 32'sd662832, 32'sd2907518, 32'sd496053, -32'sd2981578, -32'sd5710922, -32'sd4290519, -32'sd4358050, -32'sd3418115, -32'sd3603827, -32'sd2543956, -32'sd3633375, -32'sd1924734, -32'sd829040, -32'sd2072288, -32'sd2456096, 32'sd1493374, 32'sd652627, -32'sd1563464, -32'sd2061535, -32'sd3113223, -32'sd600722, 32'sd1376572, 32'sd459685, -32'sd1247751, -32'sd900524, 32'sd184040, 32'sd2324447, -32'sd67287, -32'sd557766, -32'sd520988, -32'sd1782543, -32'sd3816345, -32'sd6582985, -32'sd1602726, -32'sd1757448, -32'sd4061068, -32'sd3642345, -32'sd1976103, -32'sd3203839, -32'sd2712149, -32'sd1037970, 32'sd525300, 32'sd712490, -32'sd536400, -32'sd265117, 32'sd959611, -32'sd1374997, -32'sd2799359, -32'sd1669091, 32'sd836548, -32'sd1032034, -32'sd1553049, -32'sd402625, -32'sd882823, 32'sd915682, -32'sd1988100, -32'sd1529623, -32'sd953245, -32'sd2683759, -32'sd2455958, -32'sd6550917, -32'sd4297357, -32'sd1873559, -32'sd2142858, -32'sd3368892, -32'sd2352918, -32'sd3822079, -32'sd1624222, 32'sd1297008, 32'sd433846, 32'sd281982, 32'sd909447, -32'sd708019, 32'sd3132399, -32'sd484165, -32'sd2944871, 32'sd1010121, -32'sd1063898, -32'sd65904, 32'sd233923, -32'sd452055, 32'sd638090, 32'sd1096982, -32'sd54417, -32'sd688863, -32'sd3156301, -32'sd1128533, -32'sd4762188, -32'sd4242772, -32'sd1615572, -32'sd277904, -32'sd317382, -32'sd287062, -32'sd2981120, -32'sd917219, -32'sd2308160, 32'sd1528154, -32'sd1229628, 32'sd1280635, -32'sd785428, 32'sd227883, -32'sd365175, -32'sd2547622, 32'sd0, 32'sd636624, -32'sd33946, -32'sd632946, 32'sd2215743, -32'sd667268, 32'sd340343, -32'sd645298, -32'sd807191, -32'sd2514519, -32'sd1025486, -32'sd920321, -32'sd4759939, -32'sd2610363, -32'sd1818718, -32'sd896391, 32'sd825431, -32'sd1107458, 32'sd1726905, 32'sd429692, 32'sd678297, 32'sd396179, -32'sd567276, 32'sd1638788, 32'sd602374, -32'sd2683299, -32'sd2860864, -32'sd1549532, 32'sd139330, -32'sd293006, 32'sd1510788, -32'sd3602674, -32'sd1354570, -32'sd1646907, -32'sd423676, -32'sd1680487, -32'sd2598856, -32'sd2501396, -32'sd449472, -32'sd2824340, -32'sd1701415, -32'sd1573274, -32'sd1651058, -32'sd2264369, -32'sd2942514, -32'sd391816, -32'sd286487, 32'sd416337, 32'sd647854, 32'sd201681, 32'sd866408, -32'sd1492261, -32'sd979621, -32'sd1467785, -32'sd2497171, 32'sd114244, -32'sd2243387, -32'sd586387, -32'sd2390020, -32'sd1824525, 32'sd3031334, 32'sd734473, 32'sd1047262, -32'sd684477, -32'sd2167090, -32'sd1672102, -32'sd3888006, -32'sd2083407, -32'sd512148, 32'sd1152008, -32'sd174254, 32'sd499266, -32'sd346214, 32'sd495205, -32'sd363032, 32'sd31744, -32'sd29058, -32'sd965204, -32'sd2953717, 32'sd137856, -32'sd2113604, -32'sd1462242, -32'sd1310305, 32'sd250692, 32'sd0, -32'sd1830673, -32'sd939735, -32'sd1515989, -32'sd422447, 32'sd516882, -32'sd393101, 32'sd615233, 32'sd241445, -32'sd25748, 32'sd2810871, 32'sd2549987, 32'sd3629900, 32'sd2762891, 32'sd1479196, 32'sd1405260, -32'sd98944, -32'sd1637007, -32'sd1171439, -32'sd516995, 32'sd1139442, 32'sd594598, -32'sd59055, -32'sd1940064, -32'sd1174184, 32'sd459815, -32'sd451327, -32'sd695370, 32'sd712672, 32'sd1966225, 32'sd1293803, 32'sd758730, -32'sd1703900, -32'sd1916308, 32'sd1672099, -32'sd983918, -32'sd73009, 32'sd770239, 32'sd470989, 32'sd3609871, 32'sd3335881, 32'sd1875250, 32'sd233467, 32'sd1518790, 32'sd938611, 32'sd956801, -32'sd999894, 32'sd1207083, -32'sd14598, 32'sd2143149, -32'sd765726, 32'sd1550505, 32'sd1332816, 32'sd1613284, 32'sd587121, -32'sd2671770, 32'sd894747, -32'sd5199, -32'sd693868, -32'sd1396757, -32'sd1245014, 32'sd883987, 32'sd1213310, 32'sd601615, 32'sd3323429, 32'sd2926684, 32'sd3177216, 32'sd2206892, 32'sd948419, 32'sd2669298, 32'sd1530431, 32'sd1678795, 32'sd1722774, 32'sd3461224, 32'sd948837, -32'sd428082, -32'sd676115, -32'sd781331, 32'sd2586964, 32'sd282467, -32'sd2329608, 32'sd216406, 32'sd1506213, -32'sd2555038, 32'sd0, -32'sd818285, 32'sd251149, -32'sd23554, 32'sd252252, -32'sd1761494, 32'sd1436946, 32'sd331912, -32'sd1240870, 32'sd1864315, 32'sd258737, 32'sd809849, 32'sd2195946, 32'sd1307462, 32'sd2351387, 32'sd634618, 32'sd382740, 32'sd932242, 32'sd541429, -32'sd1540436, 32'sd49795, -32'sd2556096, 32'sd267458, 32'sd489456, -32'sd2828506, -32'sd1114159, -32'sd2916354, 32'sd0, 32'sd0, 32'sd0, 32'sd720067, 32'sd34027, -32'sd926819, 32'sd2144270, 32'sd700209, 32'sd263212, 32'sd1138420, -32'sd299858, -32'sd1190989, 32'sd1169572, 32'sd869705, -32'sd1965459, 32'sd2462725, 32'sd587246, -32'sd659897, 32'sd761462, 32'sd851059, -32'sd1300642, -32'sd2074138, -32'sd807059, -32'sd1076778, 32'sd1264238, 32'sd2054954, 32'sd387554, -32'sd356764, 32'sd0, 32'sd0, 32'sd0, -32'sd1454135, 32'sd940712, 32'sd1249254, -32'sd1118989, -32'sd62886, 32'sd1709399, -32'sd927504, 32'sd1189429, -32'sd1810741, 32'sd34006, 32'sd922760, 32'sd590015, -32'sd337412, 32'sd839384, 32'sd477878, 32'sd1783727, -32'sd188753, 32'sd1126095, 32'sd156105, 32'sd3343930, 32'sd606800, -32'sd597554, -32'sd384310, -32'sd2766988, -32'sd2009296, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd663738, -32'sd22598, -32'sd231363, -32'sd788353, 32'sd398104, 32'sd255750, 32'sd8997, 32'sd200825, -32'sd1102432, -32'sd92368, 32'sd810456, 32'sd713781, 32'sd66268, 32'sd1875131, 32'sd1216656, 32'sd1439188, 32'sd2500608, -32'sd68562, 32'sd72468, 32'sd784301, -32'sd2298818, -32'sd1303728, -32'sd2502802, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1705616, -32'sd402317, 32'sd2088514, 32'sd1698095, 32'sd647661, -32'sd386150, 32'sd1566116, -32'sd101938, -32'sd56166, 32'sd2906121, 32'sd171482, 32'sd200201, 32'sd620269, 32'sd644079, -32'sd595223, 32'sd1156727, 32'sd528126, 32'sd100883, -32'sd2027380, -32'sd1809730, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd40658, -32'sd1556520, 32'sd601690, -32'sd465911, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd776496, -32'sd83241, -32'sd253191, 32'sd162859, 32'sd498634, -32'sd273688, -32'sd199403, 32'sd172860, -32'sd32714, -32'sd33814, 32'sd2365627, -32'sd1246521, -32'sd950092, 32'sd1082181, 32'sd1396402, 32'sd1460867, 32'sd376486, 32'sd152134, -32'sd709354, -32'sd270264, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2176076, -32'sd903719, -32'sd1077666, 32'sd480983, -32'sd1525793, -32'sd1593547, -32'sd974287, 32'sd1986493, -32'sd174034, 32'sd2998894, -32'sd1098447, -32'sd710081, 32'sd1139376, 32'sd2186490, 32'sd2550614, 32'sd1226610, 32'sd2303864, 32'sd944700, 32'sd3545482, 32'sd632529, 32'sd1315597, 32'sd970727, -32'sd1760219, 32'sd2353465, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd943010, 32'sd676344, -32'sd171708, -32'sd657122, -32'sd124768, 32'sd372434, 32'sd418236, 32'sd4134778, 32'sd2750200, 32'sd560703, 32'sd628389, 32'sd2506191, 32'sd307753, 32'sd1316845, -32'sd167715, 32'sd2468395, 32'sd837285, 32'sd935855, 32'sd2310540, 32'sd1564096, 32'sd1968818, 32'sd966984, 32'sd2498243, -32'sd2640833, 32'sd194626, 32'sd0, 32'sd0, -32'sd613707, 32'sd41748, -32'sd846776, 32'sd454556, 32'sd821400, 32'sd249299, -32'sd343290, 32'sd37207, 32'sd114602, -32'sd10353, 32'sd734351, -32'sd325433, 32'sd120023, 32'sd490402, 32'sd666904, 32'sd1710970, 32'sd1216268, 32'sd1524133, 32'sd2282518, 32'sd1944174, 32'sd1350163, 32'sd2421968, 32'sd1771948, 32'sd19168, 32'sd674051, 32'sd611031, -32'sd617468, 32'sd0, 32'sd1015919, 32'sd1531100, -32'sd589987, -32'sd1243543, 32'sd503690, -32'sd247249, -32'sd1397530, -32'sd1121375, -32'sd835789, 32'sd1861814, 32'sd2227984, 32'sd776175, 32'sd1757200, 32'sd2296086, 32'sd1598298, 32'sd1999855, 32'sd1738650, 32'sd3176805, 32'sd554124, 32'sd1620248, 32'sd3220144, 32'sd3560008, 32'sd592178, 32'sd415924, -32'sd1643843, -32'sd245869, -32'sd47879, 32'sd0, 32'sd1028558, -32'sd736819, -32'sd59669, 32'sd376237, -32'sd654533, -32'sd991615, -32'sd963241, -32'sd1309977, 32'sd513157, 32'sd1874805, 32'sd1587262, 32'sd1800332, 32'sd139486, 32'sd3437030, -32'sd371427, 32'sd990520, 32'sd661589, -32'sd503254, 32'sd329930, 32'sd3738244, 32'sd537538, 32'sd543887, 32'sd2480259, 32'sd3689160, 32'sd1902383, 32'sd1199600, 32'sd2488130, 32'sd1178074, 32'sd607133, -32'sd181994, -32'sd181806, 32'sd64884, 32'sd902195, 32'sd490219, 32'sd2011397, 32'sd1587239, 32'sd1045066, 32'sd3344755, 32'sd2404568, 32'sd3082380, 32'sd2723621, 32'sd838877, -32'sd867756, 32'sd648653, -32'sd461769, 32'sd1965608, 32'sd1148056, 32'sd1626108, -32'sd158009, 32'sd1485867, 32'sd1459583, -32'sd46833, 32'sd2252266, 32'sd98291, -32'sd870798, 32'sd2300965, 32'sd699489, 32'sd257595, 32'sd252419, 32'sd1060070, 32'sd455734, -32'sd85739, 32'sd2476180, 32'sd2313950, 32'sd1348907, 32'sd1894511, 32'sd2507105, 32'sd426743, 32'sd534584, 32'sd2793899, 32'sd666028, -32'sd2688826, -32'sd608350, -32'sd3252879, -32'sd2609657, -32'sd3465660, -32'sd4163003, -32'sd4203938, -32'sd1308649, -32'sd3175138, -32'sd2340980, 32'sd504306, 32'sd367224, -32'sd261088, 32'sd732922, 32'sd1013998, -32'sd900148, -32'sd418943, 32'sd333373, 32'sd569005, 32'sd1247822, 32'sd3128299, 32'sd2995138, 32'sd1973008, 32'sd2424877, -32'sd530799, -32'sd2564484, -32'sd3713779, -32'sd4411253, -32'sd5638991, -32'sd8407115, -32'sd8822992, -32'sd8821159, -32'sd6973840, -32'sd5369449, -32'sd4637857, -32'sd1845068, 32'sd65841, -32'sd3070006, -32'sd175594, 32'sd1138404, 32'sd1159706, -32'sd894484, 32'sd494177, 32'sd201491, 32'sd429085, 32'sd1678100, 32'sd1651284, 32'sd2406908, 32'sd2475419, 32'sd963958, 32'sd1247109, -32'sd1669982, -32'sd1405151, -32'sd4235157, -32'sd7260633, -32'sd4463628, -32'sd3556320, -32'sd2526858, -32'sd6555241, -32'sd7397846, -32'sd6066990, -32'sd5405042, -32'sd5930391, -32'sd1474922, -32'sd2227161, -32'sd2044070, -32'sd127302, 32'sd355597, 32'sd281183, -32'sd576353, -32'sd312432, 32'sd332957, 32'sd484253, -32'sd1038975, 32'sd455810, -32'sd156435, -32'sd878808, 32'sd784274, -32'sd738154, -32'sd1081557, -32'sd1068928, -32'sd4595884, -32'sd3708538, -32'sd2497866, 32'sd3481387, 32'sd2545909, 32'sd1416313, -32'sd1707476, -32'sd3275810, -32'sd3257653, -32'sd2223105, 32'sd850461, -32'sd3118665, -32'sd663732, -32'sd31004, -32'sd11015, 32'sd550822, -32'sd484901, -32'sd593848, 32'sd3686004, -32'sd1126479, 32'sd748897, 32'sd1236837, -32'sd759926, 32'sd3176190, 32'sd468295, -32'sd34381, -32'sd210734, -32'sd1341092, -32'sd2938110, -32'sd2239217, -32'sd339513, 32'sd1132367, 32'sd1979868, 32'sd706914, 32'sd106321, 32'sd740080, 32'sd1188086, -32'sd940860, -32'sd179392, -32'sd3749373, -32'sd2912086, -32'sd1308319, 32'sd2332409, 32'sd357770, -32'sd507861, -32'sd53245, 32'sd181693, -32'sd719612, 32'sd1634628, -32'sd2731680, -32'sd1114565, -32'sd109879, -32'sd1742180, 32'sd191917, 32'sd298282, -32'sd2724639, -32'sd11260, 32'sd190466, -32'sd3670140, -32'sd633058, 32'sd791627, -32'sd630667, 32'sd1536203, 32'sd1982007, 32'sd99003, 32'sd799192, 32'sd743751, 32'sd2540634, -32'sd1235742, -32'sd3271044, 32'sd210303, 32'sd1589924, -32'sd897894, 32'sd234559, 32'sd1484435, 32'sd611354, -32'sd4452393, 32'sd67424, 32'sd2041814, -32'sd226793, -32'sd2258912, 32'sd734308, -32'sd1587033, -32'sd684383, 32'sd55240, 32'sd6712, -32'sd1161181, -32'sd79395, -32'sd1076504, -32'sd870888, 32'sd625493, 32'sd1784876, 32'sd675280, -32'sd903312, 32'sd93509, 32'sd684226, -32'sd1124240, -32'sd1976139, -32'sd408120, -32'sd1013753, 32'sd859471, 32'sd46741, 32'sd875040, -32'sd2387298, -32'sd5236225, -32'sd4156480, -32'sd4341752, -32'sd208456, 32'sd1004211, 32'sd1820157, -32'sd225769, 32'sd1196277, 32'sd560222, -32'sd526586, -32'sd1345951, -32'sd469780, 32'sd245970, -32'sd256128, -32'sd668555, -32'sd2143494, 32'sd282264, 32'sd304390, 32'sd339039, 32'sd2332805, -32'sd167980, -32'sd1137391, -32'sd791437, 32'sd46286, -32'sd784799, 32'sd515665, 32'sd1516602, -32'sd1065966, -32'sd5393119, -32'sd3570851, -32'sd5895115, -32'sd3343735, -32'sd707700, 32'sd359707, 32'sd319549, -32'sd482747, 32'sd139658, 32'sd617492, 32'sd971090, -32'sd1914231, -32'sd279529, 32'sd1151717, -32'sd701743, -32'sd1208594, 32'sd264712, 32'sd390328, -32'sd605442, -32'sd295140, 32'sd490908, 32'sd44192, 32'sd765679, 32'sd0, 32'sd381694, -32'sd205361, 32'sd1387124, -32'sd1991425, -32'sd4454775, -32'sd1705391, -32'sd2160561, -32'sd1603449, -32'sd1630077, -32'sd55233, -32'sd301723, 32'sd1978356, 32'sd194, 32'sd896022, -32'sd96766, -32'sd374455, 32'sd788503, -32'sd300751, -32'sd1849146, -32'sd1177612, 32'sd92758, 32'sd1095304, 32'sd2436664, 32'sd860000, -32'sd404417, -32'sd2038872, 32'sd842117, 32'sd420757, -32'sd743400, -32'sd443525, 32'sd61092, 32'sd734550, -32'sd888005, -32'sd5393068, -32'sd1529581, -32'sd915313, -32'sd3362267, -32'sd1967126, -32'sd2738001, -32'sd3915220, -32'sd952154, -32'sd697936, -32'sd782509, 32'sd150946, 32'sd1083326, -32'sd244049, -32'sd2056800, -32'sd790948, 32'sd1195336, 32'sd347717, 32'sd358450, 32'sd1279210, 32'sd448009, 32'sd69683, 32'sd1940816, 32'sd201859, 32'sd846786, 32'sd81683, -32'sd928153, 32'sd175194, -32'sd33990, 32'sd179050, -32'sd3984810, 32'sd948015, -32'sd2026009, -32'sd1416459, -32'sd3244254, -32'sd2073698, -32'sd1710439, -32'sd1492289, -32'sd247135, 32'sd1680386, 32'sd1522313, 32'sd555731, -32'sd259407, 32'sd515623, 32'sd5016, 32'sd1763881, 32'sd165576, 32'sd496079, 32'sd1577187, 32'sd987196, -32'sd33196, 32'sd0, 32'sd367697, 32'sd2033935, -32'sd321728, 32'sd938574, 32'sd1772766, 32'sd1016008, -32'sd1775294, 32'sd756689, 32'sd3161431, 32'sd446123, 32'sd2139934, 32'sd1515320, 32'sd2878110, 32'sd217024, 32'sd337120, 32'sd1886726, -32'sd961317, 32'sd1249329, 32'sd759994, -32'sd1796000, -32'sd109008, 32'sd2143090, -32'sd487776, -32'sd1553936, 32'sd931288, 32'sd491252, 32'sd402086, 32'sd2452228, 32'sd668517, 32'sd2350584, 32'sd10954, 32'sd1369352, 32'sd3022365, 32'sd789465, 32'sd290553, 32'sd3672057, 32'sd3339891, 32'sd2867237, 32'sd3610228, 32'sd3874862, 32'sd1751212, 32'sd2468541, 32'sd1541755, 32'sd3019488, 32'sd2556069, 32'sd1873122, 32'sd2892352, 32'sd1722257, 32'sd3285976, 32'sd493477, 32'sd159756, 32'sd338387, 32'sd1988797, 32'sd938255, -32'sd242611, 32'sd882583, 32'sd1046467, 32'sd223753, 32'sd1174848, 32'sd1908161, 32'sd543842, -32'sd1048933, 32'sd2993237, 32'sd4490601, 32'sd4139440, 32'sd3741372, 32'sd1970093, 32'sd777924, -32'sd1443456, 32'sd4418490, 32'sd458337, 32'sd616755, 32'sd1168110, 32'sd2757158, 32'sd1274971, 32'sd2575351, -32'sd400543, -32'sd1575881, 32'sd1050873, 32'sd527478, 32'sd113161, -32'sd113072, 32'sd1228565, 32'sd0, -32'sd102952, 32'sd2065484, 32'sd354820, 32'sd2423376, 32'sd282528, 32'sd446890, -32'sd918894, 32'sd1759546, 32'sd1468155, 32'sd1895288, 32'sd1193132, 32'sd701285, 32'sd836233, 32'sd1531116, 32'sd1864524, -32'sd65563, 32'sd827267, 32'sd515460, 32'sd1075537, 32'sd2239169, 32'sd1241200, 32'sd509354, -32'sd219110, 32'sd1232204, 32'sd566270, -32'sd243500, 32'sd0, 32'sd0, 32'sd0, -32'sd498703, -32'sd411135, -32'sd2536626, 32'sd1160048, 32'sd1921606, -32'sd961339, 32'sd1662663, 32'sd386825, -32'sd1996858, 32'sd174112, 32'sd3183146, 32'sd319845, -32'sd1132941, 32'sd613704, 32'sd2103813, -32'sd495128, 32'sd1600016, -32'sd155287, 32'sd547601, 32'sd724871, 32'sd1418178, 32'sd632616, 32'sd1123345, -32'sd94258, -32'sd621586, 32'sd0, 32'sd0, 32'sd0, 32'sd475208, 32'sd957655, -32'sd1899201, -32'sd3322901, -32'sd852889, -32'sd49614, -32'sd2001200, 32'sd205291, -32'sd137191, -32'sd472585, 32'sd806684, 32'sd1070223, 32'sd642694, -32'sd516681, -32'sd377901, -32'sd101133, 32'sd1634755, 32'sd933649, -32'sd1028596, 32'sd1813489, 32'sd2057659, 32'sd1099045, 32'sd1293622, -32'sd318865, 32'sd1438640, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2560247, -32'sd319359, 32'sd2021977, 32'sd577335, 32'sd547105, 32'sd1635326, 32'sd1263965, 32'sd2055102, 32'sd139119, 32'sd1425035, -32'sd184258, -32'sd411797, 32'sd2053095, -32'sd1001558, 32'sd134107, 32'sd1459104, -32'sd5184588, -32'sd425241, 32'sd47424, -32'sd89234, 32'sd1044969, -32'sd563050, 32'sd1114036, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd346840, 32'sd630492, -32'sd645949, 32'sd779994, -32'sd227126, 32'sd638585, 32'sd883930, 32'sd1008508, 32'sd1441982, 32'sd720304, 32'sd311437, -32'sd551766, 32'sd160899, 32'sd674447, -32'sd1164954, 32'sd1442433, -32'sd521395, -32'sd604638, -32'sd1895340, 32'sd906787, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3576969, -32'sd4835674, -32'sd4617118, -32'sd4949272, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3431204, -32'sd4510826, -32'sd4890322, -32'sd3834015, -32'sd5626622, -32'sd2343147, 32'sd1767932, 32'sd909276, -32'sd793683, 32'sd197926, 32'sd415838, -32'sd2980322, -32'sd820612, -32'sd425888, 32'sd792897, -32'sd1193181, -32'sd4211606, -32'sd5196051, -32'sd4635927, -32'sd5487936, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3512355, 32'sd790225, -32'sd5343550, -32'sd5731051, -32'sd4221732, -32'sd7121648, -32'sd3611402, 32'sd1636905, -32'sd133415, 32'sd1502871, 32'sd1943221, -32'sd2195638, -32'sd636230, -32'sd724988, -32'sd859718, 32'sd1534481, -32'sd1939623, 32'sd816282, 32'sd928516, -32'sd1435459, 32'sd2426429, 32'sd1788988, -32'sd941091, -32'sd3610965, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3723075, 32'sd1656424, 32'sd207119, -32'sd1437263, -32'sd5019093, -32'sd4627323, 32'sd4062092, -32'sd2012905, 32'sd802160, 32'sd1265661, -32'sd1000480, 32'sd837098, 32'sd3724402, 32'sd1086896, 32'sd728179, -32'sd744230, 32'sd1799288, 32'sd1226645, 32'sd2356960, 32'sd354530, 32'sd1640645, 32'sd23989, -32'sd2439655, -32'sd556553, -32'sd5645324, 32'sd0, 32'sd0, -32'sd4650396, -32'sd281462, 32'sd818283, 32'sd1088084, -32'sd2977697, -32'sd2889169, -32'sd5066601, 32'sd75406, -32'sd1291616, 32'sd763644, 32'sd308338, 32'sd1041063, 32'sd760301, 32'sd2530938, 32'sd810897, 32'sd2030611, 32'sd1015605, 32'sd2178786, 32'sd3172564, 32'sd2086721, 32'sd2405516, 32'sd1093166, -32'sd2108355, 32'sd1930869, 32'sd53320, 32'sd58672, -32'sd4724482, 32'sd0, 32'sd101312, 32'sd803356, -32'sd1457491, 32'sd195349, -32'sd2422908, -32'sd3310079, -32'sd1149590, 32'sd836463, 32'sd1083248, 32'sd2433651, -32'sd301211, 32'sd1405580, -32'sd1107621, 32'sd2476564, -32'sd1088521, 32'sd1533627, 32'sd1599236, -32'sd1411065, -32'sd1331930, 32'sd785566, 32'sd702431, -32'sd210668, 32'sd336592, 32'sd844863, 32'sd802473, 32'sd168954, -32'sd5818277, 32'sd0, -32'sd4173117, -32'sd4553055, -32'sd163675, 32'sd4867142, 32'sd228188, -32'sd607426, 32'sd414403, 32'sd1380082, -32'sd983158, -32'sd3324065, -32'sd1098748, 32'sd949151, -32'sd2104646, -32'sd222098, -32'sd557591, -32'sd3765506, -32'sd1321119, -32'sd5724106, -32'sd2866984, -32'sd104203, 32'sd270092, 32'sd392823, 32'sd4692460, 32'sd2628403, 32'sd98319, -32'sd243198, -32'sd770824, -32'sd3777154, -32'sd6342725, -32'sd3271005, -32'sd4456633, 32'sd2113917, -32'sd518031, -32'sd835689, -32'sd478744, -32'sd524403, -32'sd411435, -32'sd28818, 32'sd404654, -32'sd266374, 32'sd977626, -32'sd1205918, -32'sd1227796, -32'sd4411385, -32'sd3542520, -32'sd5123294, -32'sd2576196, -32'sd2936267, 32'sd758720, 32'sd1695519, 32'sd2973431, 32'sd3001231, -32'sd314311, 32'sd1287900, 32'sd804476, -32'sd5661283, -32'sd2184896, -32'sd5682648, -32'sd4195874, 32'sd400279, 32'sd588121, -32'sd51638, 32'sd1172850, 32'sd602747, 32'sd3043583, -32'sd567008, -32'sd483110, 32'sd1529766, 32'sd1101136, -32'sd2639055, -32'sd59257, -32'sd4143578, -32'sd4163370, -32'sd3830318, -32'sd3475642, -32'sd1985198, -32'sd773539, -32'sd1891598, 32'sd1044498, 32'sd282306, 32'sd123262, 32'sd2547271, 32'sd383441, -32'sd4417260, -32'sd6388193, -32'sd5462822, -32'sd6879696, -32'sd2184929, -32'sd2203506, -32'sd946596, 32'sd1094768, 32'sd2640108, 32'sd618558, 32'sd421051, -32'sd991342, -32'sd1737454, -32'sd4414731, -32'sd3541847, -32'sd1703951, -32'sd1061746, -32'sd1028478, -32'sd2571043, 32'sd380715, 32'sd377749, 32'sd390949, -32'sd1520413, -32'sd642766, -32'sd3022188, 32'sd632411, 32'sd1222902, -32'sd983700, -32'sd5353566, -32'sd4274554, -32'sd7238599, -32'sd6821179, 32'sd1112713, -32'sd1052917, 32'sd863249, 32'sd3295563, 32'sd2593203, 32'sd94459, 32'sd150162, -32'sd372666, -32'sd1027323, -32'sd5586504, -32'sd6090845, -32'sd1989641, -32'sd2600469, 32'sd873052, -32'sd810189, 32'sd1520872, -32'sd844116, -32'sd964801, 32'sd600801, -32'sd2644866, -32'sd407577, 32'sd1340504, -32'sd608051, 32'sd135170, -32'sd4999160, -32'sd2840355, -32'sd1119262, -32'sd5657460, -32'sd1679027, 32'sd78911, 32'sd98814, 32'sd1579845, 32'sd2866217, 32'sd4473141, 32'sd1692361, 32'sd757324, 32'sd4023419, -32'sd5208034, -32'sd3781914, -32'sd1156799, -32'sd462457, -32'sd2369515, -32'sd3269116, 32'sd463409, -32'sd609502, -32'sd798955, 32'sd1342132, -32'sd83334, -32'sd1111474, -32'sd227838, -32'sd1205250, -32'sd3627136, -32'sd1869046, -32'sd2363745, -32'sd3677777, -32'sd4530830, -32'sd753556, -32'sd764191, 32'sd1731841, 32'sd1968326, 32'sd2480185, 32'sd4630092, 32'sd2480670, 32'sd1219034, 32'sd2128630, -32'sd736790, -32'sd5211230, -32'sd1807924, 32'sd1850685, -32'sd80916, -32'sd734195, 32'sd944881, 32'sd2865564, 32'sd2806245, 32'sd397051, 32'sd885906, 32'sd3188652, -32'sd506176, 32'sd60542, -32'sd4839340, -32'sd5645463, -32'sd5050241, -32'sd1653679, -32'sd1983309, -32'sd2753083, -32'sd490122, -32'sd1240422, 32'sd3040564, 32'sd1542430, 32'sd1803410, 32'sd2275987, 32'sd2550437, 32'sd4938064, 32'sd2510951, 32'sd505175, 32'sd2661149, 32'sd2977023, 32'sd2687301, 32'sd2857589, 32'sd3069317, 32'sd2143247, 32'sd3512494, 32'sd2812178, 32'sd1884025, 32'sd1159477, -32'sd3087642, -32'sd3892753, -32'sd5571053, -32'sd4819410, -32'sd4628031, -32'sd3495608, -32'sd202402, -32'sd1899474, -32'sd1044158, -32'sd2059920, -32'sd817233, 32'sd653766, 32'sd1216936, 32'sd1873930, 32'sd4465381, 32'sd2491359, 32'sd2555920, 32'sd1878915, 32'sd1334572, 32'sd3898997, 32'sd1360497, -32'sd1656200, -32'sd763246, -32'sd375459, 32'sd276643, 32'sd2003522, -32'sd134469, -32'sd2148071, -32'sd955202, -32'sd3199785, -32'sd6008867, -32'sd5496700, -32'sd5275326, -32'sd2411444, 32'sd426377, -32'sd768104, -32'sd3168868, -32'sd176049, -32'sd912206, -32'sd341408, 32'sd661251, 32'sd528981, 32'sd2036235, 32'sd3801350, 32'sd2157110, 32'sd1408126, 32'sd1372905, 32'sd1964635, 32'sd2152302, -32'sd1731869, 32'sd38059, -32'sd596890, -32'sd2508694, 32'sd4008500, 32'sd3369046, -32'sd672052, 32'sd95455, -32'sd3791630, -32'sd4778020, -32'sd5340637, -32'sd5947776, -32'sd4899847, 32'sd720402, 32'sd723998, -32'sd2898813, -32'sd1258159, -32'sd2800264, 32'sd1825426, 32'sd186307, -32'sd671416, 32'sd192124, 32'sd2594907, 32'sd1702006, 32'sd3226376, 32'sd2499392, 32'sd1304340, 32'sd962322, -32'sd1675500, -32'sd702994, -32'sd2545769, -32'sd2664772, 32'sd450487, 32'sd2659241, -32'sd1149918, -32'sd612388, -32'sd5835487, -32'sd1018049, 32'sd0, -32'sd6055135, -32'sd2426036, -32'sd1724516, -32'sd634288, -32'sd630619, -32'sd2479804, -32'sd1517216, 32'sd478274, -32'sd1336402, -32'sd373224, 32'sd1043773, 32'sd1809706, 32'sd2420938, 32'sd1638482, 32'sd128656, 32'sd619256, -32'sd386604, -32'sd1529150, 32'sd290683, 32'sd225803, -32'sd400488, 32'sd1438447, -32'sd1674746, -32'sd533195, 32'sd644136, -32'sd2892469, -32'sd256775, -32'sd6037026, -32'sd5498329, -32'sd3571801, 32'sd541075, -32'sd2918548, 32'sd1247506, 32'sd1669543, -32'sd986771, -32'sd2355591, -32'sd713412, 32'sd448490, 32'sd1244184, 32'sd3727011, 32'sd6255146, 32'sd189364, 32'sd266223, 32'sd1350054, -32'sd1463464, -32'sd1850738, -32'sd2546959, -32'sd2518208, -32'sd2773513, -32'sd481615, -32'sd1258166, 32'sd1357473, -32'sd1227774, 32'sd906161, 32'sd83913, -32'sd5575959, -32'sd6106473, -32'sd4160002, -32'sd807823, -32'sd2368474, -32'sd2454052, -32'sd1121802, -32'sd4156583, -32'sd2190103, -32'sd1624783, 32'sd1326473, 32'sd2641433, -32'sd83177, 32'sd1156314, -32'sd926884, -32'sd353492, -32'sd799426, -32'sd31427, -32'sd2327541, -32'sd1189698, -32'sd2501686, 32'sd1165335, 32'sd615722, -32'sd725421, 32'sd374689, 32'sd999208, 32'sd1113604, -32'sd3949199, 32'sd0, -32'sd5793998, -32'sd2269363, -32'sd5252595, -32'sd6200668, -32'sd2550740, -32'sd2914155, -32'sd2119633, 32'sd71211, 32'sd1538329, -32'sd892887, 32'sd1609031, -32'sd56178, -32'sd1094227, 32'sd323818, -32'sd268677, -32'sd472191, 32'sd11452, -32'sd446068, -32'sd2178474, 32'sd95028, 32'sd304106, -32'sd1245032, -32'sd25695, 32'sd549153, 32'sd511692, 32'sd1576369, -32'sd761929, 32'sd364621, -32'sd1458272, -32'sd1066888, -32'sd3964493, -32'sd3450100, -32'sd4715893, -32'sd3153436, -32'sd1215097, 32'sd1455213, 32'sd3732685, 32'sd1360764, 32'sd1374566, 32'sd1089209, 32'sd3663295, 32'sd2016693, 32'sd1329652, -32'sd504448, 32'sd1103490, 32'sd1514434, 32'sd272266, -32'sd987875, -32'sd894274, 32'sd449112, 32'sd875333, -32'sd1211997, -32'sd254051, -32'sd777949, -32'sd4234434, -32'sd253215, 32'sd503473, -32'sd2731399, -32'sd1468358, -32'sd1546415, -32'sd3319707, -32'sd2471110, -32'sd2326435, -32'sd1396793, -32'sd429551, 32'sd548524, 32'sd92129, 32'sd1372040, 32'sd1174045, -32'sd775189, 32'sd1355369, 32'sd792339, -32'sd252206, 32'sd794641, 32'sd702854, 32'sd906884, -32'sd1079662, -32'sd2521887, 32'sd1251352, -32'sd358592, 32'sd518584, 32'sd495624, -32'sd5212679, 32'sd0, 32'sd90822, -32'sd368081, -32'sd1673296, 32'sd2706569, -32'sd2350541, -32'sd3454110, -32'sd1226113, -32'sd1125606, -32'sd1643627, -32'sd880725, -32'sd1927427, -32'sd1300586, -32'sd1051373, 32'sd1049315, 32'sd603985, 32'sd1711337, 32'sd2031148, 32'sd340800, -32'sd397070, -32'sd453465, 32'sd514607, -32'sd438910, 32'sd2759165, -32'sd1342506, -32'sd347578, -32'sd255048, 32'sd0, 32'sd0, 32'sd0, -32'sd4825491, -32'sd2232308, -32'sd1477663, 32'sd2030526, -32'sd816360, -32'sd550934, -32'sd2743962, -32'sd482919, 32'sd363244, 32'sd2187931, 32'sd149628, 32'sd1201625, 32'sd299962, -32'sd65821, 32'sd2927736, -32'sd258962, 32'sd176961, -32'sd638054, -32'sd141234, 32'sd833566, 32'sd1636702, 32'sd790761, -32'sd1216546, -32'sd909163, -32'sd4256830, 32'sd0, 32'sd0, 32'sd0, -32'sd4248990, -32'sd5223528, -32'sd2848, -32'sd191172, 32'sd107583, -32'sd1815650, -32'sd1675618, -32'sd2491838, -32'sd117516, -32'sd449374, -32'sd2937025, -32'sd442083, 32'sd956142, 32'sd393703, -32'sd1468130, -32'sd706506, 32'sd662012, 32'sd120896, 32'sd1308418, -32'sd200820, 32'sd1191889, 32'sd1102267, -32'sd1324119, -32'sd6122832, -32'sd5511152, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3891374, -32'sd167992, -32'sd2521658, 32'sd510516, 32'sd253960, 32'sd2738879, -32'sd2361521, -32'sd2360315, -32'sd827991, -32'sd2025209, -32'sd577415, -32'sd279502, -32'sd1968674, -32'sd1543482, 32'sd1882071, 32'sd871575, 32'sd216699, 32'sd891582, 32'sd433123, -32'sd1937970, -32'sd5383645, -32'sd4168849, -32'sd5040430, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3855348, -32'sd6290372, -32'sd261356, 32'sd136782, -32'sd1475308, -32'sd2831272, -32'sd944609, 32'sd690694, -32'sd940320, -32'sd2336091, -32'sd2677481, -32'sd4504528, -32'sd2410555, -32'sd3081918, -32'sd5853944, -32'sd5329853, -32'sd5702531, -32'sd5956639, -32'sd3674140, -32'sd3519987, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1008468, -32'sd3495392, -32'sd1388453, -32'sd1694174, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1341824, -32'sd2947993, -32'sd913724, -32'sd586181, -32'sd5974, 32'sd1253736, -32'sd394183, 32'sd2080444, 32'sd1635363, -32'sd1080533, 32'sd1919563, -32'sd156707, 32'sd1331747, 32'sd1271885, -32'sd534952, -32'sd1039804, 32'sd676627, -32'sd838653, -32'sd1784373, -32'sd2363477, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3151169, -32'sd3345343, 32'sd1221740, 32'sd111092, 32'sd1074484, 32'sd1385931, 32'sd1147940, 32'sd3167572, 32'sd277237, 32'sd1039715, 32'sd334528, 32'sd284360, 32'sd1646215, -32'sd434438, -32'sd72233, 32'sd2938485, 32'sd998200, -32'sd1877143, 32'sd409008, 32'sd2062882, 32'sd203313, -32'sd2583822, -32'sd3058750, -32'sd2565628, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd723017, -32'sd138276, 32'sd48684, 32'sd946485, 32'sd983518, 32'sd964049, -32'sd992441, 32'sd2544956, -32'sd512484, -32'sd1230126, -32'sd1156454, -32'sd828003, -32'sd440693, -32'sd2608623, -32'sd653440, 32'sd1526982, -32'sd666332, 32'sd357415, -32'sd2999248, 32'sd1123061, -32'sd647349, 32'sd1539497, 32'sd1387035, -32'sd1041155, -32'sd3469232, 32'sd0, 32'sd0, -32'sd2022794, 32'sd590848, -32'sd948094, 32'sd705533, -32'sd357036, -32'sd763041, -32'sd1327518, 32'sd1536775, 32'sd535650, 32'sd1614008, -32'sd366697, -32'sd587751, 32'sd593817, -32'sd445024, -32'sd419811, -32'sd305291, -32'sd989268, -32'sd2639107, 32'sd48647, 32'sd1387318, -32'sd221041, -32'sd547381, 32'sd346117, -32'sd1761103, -32'sd989773, -32'sd41606, -32'sd2111315, 32'sd0, -32'sd671926, 32'sd196430, 32'sd112547, -32'sd316398, -32'sd1790498, 32'sd2437572, -32'sd127052, -32'sd1746723, -32'sd990624, -32'sd225601, 32'sd265102, -32'sd2746985, 32'sd489465, 32'sd1291697, -32'sd2018359, 32'sd1720602, 32'sd1494285, 32'sd991493, -32'sd466714, 32'sd1042274, -32'sd1355902, -32'sd1552211, -32'sd179680, -32'sd1481468, 32'sd1362133, 32'sd1006680, 32'sd513830, 32'sd0, -32'sd1946347, -32'sd413672, 32'sd1142940, 32'sd599822, -32'sd780177, -32'sd461414, 32'sd1532416, -32'sd2290115, 32'sd896161, -32'sd1297955, 32'sd44894, -32'sd2046206, -32'sd3523115, -32'sd1454472, 32'sd182151, -32'sd859935, 32'sd2008172, 32'sd1621148, -32'sd357414, -32'sd1988806, -32'sd3129884, -32'sd504889, -32'sd2069651, -32'sd3301923, -32'sd2112881, -32'sd1977064, -32'sd5315544, -32'sd2654782, -32'sd2396396, -32'sd1803476, 32'sd235724, -32'sd1167848, 32'sd219736, 32'sd374847, -32'sd602300, -32'sd1149445, -32'sd2539873, -32'sd1903803, -32'sd801696, -32'sd2053083, -32'sd1185529, -32'sd318650, -32'sd3156257, -32'sd1231762, -32'sd1490336, -32'sd1953674, -32'sd3109652, -32'sd2561799, -32'sd2256165, 32'sd671401, -32'sd3598695, -32'sd2491178, -32'sd2747153, 32'sd423939, -32'sd3238917, 32'sd616386, 32'sd585930, 32'sd1406078, -32'sd908552, -32'sd909094, -32'sd134383, 32'sd530648, -32'sd3150530, -32'sd3078973, -32'sd1770732, -32'sd1583124, -32'sd2478973, -32'sd1840631, -32'sd78669, -32'sd97395, -32'sd1453110, -32'sd1471955, -32'sd2165466, -32'sd1939458, -32'sd2214411, -32'sd3216780, -32'sd661015, -32'sd1860947, 32'sd731102, -32'sd2446463, -32'sd2426327, 32'sd1321957, -32'sd3523482, -32'sd3561393, -32'sd3620425, -32'sd2031045, 32'sd354944, 32'sd746872, -32'sd945211, -32'sd1787630, -32'sd1182327, -32'sd1219164, -32'sd1370755, -32'sd1422083, -32'sd1736942, -32'sd2211084, -32'sd1594382, 32'sd874540, -32'sd3076280, -32'sd3582013, -32'sd574457, -32'sd3229705, -32'sd3012826, -32'sd30288, -32'sd270708, 32'sd1302551, -32'sd1839686, -32'sd3631847, -32'sd1796428, -32'sd387632, -32'sd555629, -32'sd1349932, 32'sd37322, -32'sd1439611, -32'sd18916, 32'sd414536, 32'sd950740, 32'sd174852, -32'sd1549149, -32'sd2811706, -32'sd1391732, -32'sd2899452, 32'sd319922, -32'sd2049665, -32'sd1050429, -32'sd3146608, -32'sd3839657, -32'sd3905404, -32'sd1754079, -32'sd591642, -32'sd2046470, -32'sd2618349, -32'sd2580854, -32'sd1999442, -32'sd929499, 32'sd695375, -32'sd2191340, 32'sd1455396, -32'sd1608190, -32'sd2317330, -32'sd4018436, 32'sd1068438, -32'sd920301, -32'sd30971, 32'sd683508, 32'sd639559, 32'sd656726, -32'sd3430877, -32'sd1736748, -32'sd2408703, -32'sd2180740, -32'sd1717694, -32'sd4811636, -32'sd4227799, -32'sd4076309, -32'sd2744128, -32'sd2362537, -32'sd1646731, 32'sd1576883, -32'sd2846269, -32'sd1092346, -32'sd766660, -32'sd1837605, -32'sd1034659, -32'sd495870, 32'sd393562, -32'sd358567, -32'sd1053402, 32'sd791269, 32'sd50888, 32'sd1329037, -32'sd646652, 32'sd852976, 32'sd1433433, -32'sd211970, -32'sd648078, 32'sd539354, -32'sd724322, -32'sd1215064, -32'sd2915531, -32'sd3570325, -32'sd2868362, -32'sd3152764, -32'sd3912056, -32'sd2844610, -32'sd2996631, -32'sd416385, -32'sd431998, 32'sd2101593, -32'sd784165, -32'sd2284339, 32'sd2101449, 32'sd585837, -32'sd360004, -32'sd2155315, -32'sd1960277, -32'sd1265411, -32'sd968993, -32'sd397141, -32'sd1800926, 32'sd1237435, 32'sd3780446, 32'sd2814834, 32'sd3397808, 32'sd1583843, 32'sd1077562, 32'sd483928, -32'sd2055330, -32'sd690310, -32'sd1385021, -32'sd2744084, 32'sd247596, 32'sd427923, -32'sd625565, -32'sd519244, -32'sd916789, 32'sd1739708, 32'sd1508458, 32'sd647856, 32'sd151015, -32'sd1019793, -32'sd244177, -32'sd1695864, -32'sd2448564, -32'sd2976897, -32'sd1403629, -32'sd716266, -32'sd987200, -32'sd1264686, 32'sd975655, 32'sd5665344, 32'sd3207761, 32'sd1654280, 32'sd1918542, 32'sd1645114, -32'sd2593566, -32'sd1880165, -32'sd109050, -32'sd999790, 32'sd635507, -32'sd591120, 32'sd155625, -32'sd431256, 32'sd214662, 32'sd105067, 32'sd1928602, 32'sd1158684, 32'sd1626903, 32'sd2515430, 32'sd976859, -32'sd2755962, -32'sd2635051, -32'sd1703712, 32'sd461720, 32'sd2554651, -32'sd31568, -32'sd685310, 32'sd1823542, 32'sd3819214, 32'sd4623972, 32'sd2375050, 32'sd4108520, 32'sd2140060, -32'sd464376, 32'sd709199, 32'sd868875, -32'sd178163, 32'sd1663362, 32'sd1876833, -32'sd126107, 32'sd2185538, 32'sd245821, -32'sd82211, 32'sd755926, -32'sd1453193, 32'sd1694096, 32'sd2363059, -32'sd534951, -32'sd714162, -32'sd959325, 32'sd411001, -32'sd525127, -32'sd688725, -32'sd1924991, 32'sd414551, 32'sd2076753, 32'sd875853, 32'sd1277321, 32'sd1454834, 32'sd4205611, 32'sd5385197, 32'sd3881803, 32'sd3107860, 32'sd796491, 32'sd311618, 32'sd3899117, 32'sd2636606, -32'sd239856, -32'sd374220, 32'sd950565, 32'sd850446, -32'sd168686, -32'sd137235, -32'sd1121942, 32'sd717201, 32'sd2093666, 32'sd113513, 32'sd0, 32'sd17033, 32'sd1227470, 32'sd763056, -32'sd505110, 32'sd485768, 32'sd712754, -32'sd1538349, 32'sd994785, 32'sd1655880, 32'sd3363733, 32'sd2935978, 32'sd2576051, 32'sd1690934, 32'sd960848, 32'sd3284941, 32'sd3562231, -32'sd64430, 32'sd1530639, -32'sd303136, 32'sd2627955, 32'sd2717117, 32'sd1729267, -32'sd222309, -32'sd1307819, 32'sd197159, 32'sd191434, 32'sd110808, -32'sd1654701, -32'sd775175, -32'sd265122, 32'sd204377, 32'sd1632367, 32'sd1703487, -32'sd155996, 32'sd2764639, 32'sd1574382, 32'sd2171973, 32'sd837951, 32'sd805981, 32'sd3404670, 32'sd2252992, 32'sd761893, 32'sd1297425, 32'sd2425264, 32'sd1107023, 32'sd2586876, 32'sd4339671, 32'sd783736, 32'sd3383719, -32'sd551257, -32'sd203160, -32'sd1340336, 32'sd1636301, -32'sd1849383, -32'sd1888679, -32'sd393127, -32'sd3380757, -32'sd41407, -32'sd1782722, 32'sd297546, 32'sd155778, -32'sd476251, 32'sd2150179, 32'sd1690327, -32'sd742481, 32'sd1628080, 32'sd4259146, 32'sd2150462, 32'sd1382959, 32'sd1036122, 32'sd4434633, 32'sd593038, 32'sd1802039, 32'sd1626334, -32'sd1206952, 32'sd1400135, 32'sd792198, 32'sd2135528, 32'sd390207, -32'sd1721813, -32'sd263354, 32'sd2432772, -32'sd3264978, 32'sd0, -32'sd3067802, 32'sd2418542, -32'sd369896, 32'sd60734, 32'sd652739, -32'sd59140, 32'sd1066035, -32'sd2169600, -32'sd2008178, -32'sd1486556, 32'sd1062987, 32'sd815926, 32'sd471406, 32'sd3486892, 32'sd2231747, 32'sd1706849, 32'sd2679562, 32'sd2333249, 32'sd1039033, -32'sd259309, 32'sd2696010, 32'sd11075, 32'sd1126246, -32'sd1466569, 32'sd886465, 32'sd495108, -32'sd3227614, -32'sd2752295, -32'sd2313273, 32'sd355381, -32'sd1833038, -32'sd783726, 32'sd1611073, 32'sd1207406, -32'sd16599, -32'sd92870, -32'sd501898, -32'sd530884, 32'sd1688691, 32'sd35025, 32'sd2602514, 32'sd1710067, 32'sd1072872, 32'sd1822388, 32'sd845612, 32'sd940986, 32'sd2966984, 32'sd650785, 32'sd485108, 32'sd975945, 32'sd2979680, -32'sd806766, 32'sd3071481, 32'sd603694, 32'sd235452, -32'sd2759008, -32'sd1546377, 32'sd891645, -32'sd103088, 32'sd3643564, 32'sd1868385, 32'sd260594, 32'sd602860, 32'sd1335922, -32'sd585293, 32'sd318843, 32'sd2871705, 32'sd2448161, 32'sd119192, -32'sd3657069, 32'sd229994, -32'sd519182, -32'sd2050077, -32'sd523170, 32'sd568455, 32'sd495391, 32'sd1338119, 32'sd433538, -32'sd797156, -32'sd733860, -32'sd389581, 32'sd500868, -32'sd50416, 32'sd0, -32'sd491120, 32'sd743145, 32'sd780026, 32'sd1046814, 32'sd888834, -32'sd673804, -32'sd1439521, 32'sd1775207, 32'sd952003, -32'sd177763, -32'sd1677219, -32'sd1919716, -32'sd3139764, -32'sd1834646, -32'sd1362802, -32'sd917174, -32'sd1960222, 32'sd1429352, -32'sd1258824, -32'sd4789, 32'sd1077197, 32'sd958073, 32'sd946891, -32'sd26236, 32'sd113969, -32'sd3091844, 32'sd0, 32'sd0, 32'sd0, -32'sd2637644, -32'sd1828788, -32'sd74729, 32'sd1457433, -32'sd4875837, -32'sd3778025, -32'sd2164091, 32'sd273627, -32'sd4379993, -32'sd5705666, -32'sd4965790, -32'sd1685729, -32'sd4894741, -32'sd3397794, -32'sd2022116, -32'sd1178385, -32'sd762055, -32'sd70237, -32'sd132841, -32'sd101813, 32'sd586718, 32'sd714901, -32'sd869535, 32'sd862924, -32'sd929491, 32'sd0, 32'sd0, 32'sd0, -32'sd934136, -32'sd1800181, -32'sd3619006, -32'sd1603081, -32'sd128785, -32'sd2339535, 32'sd964490, -32'sd5108854, -32'sd2805208, -32'sd1076049, 32'sd427232, -32'sd1906143, -32'sd1647038, -32'sd908727, 32'sd1284817, -32'sd2575335, 32'sd1490547, 32'sd738384, 32'sd1877254, -32'sd883385, -32'sd1493595, -32'sd872084, -32'sd557276, -32'sd2780275, -32'sd2616245, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd3157554, -32'sd826155, -32'sd2449079, 32'sd342036, 32'sd742041, 32'sd1506506, -32'sd1254897, -32'sd225511, 32'sd1824258, 32'sd2067355, 32'sd1675748, -32'sd952104, 32'sd610613, -32'sd1487953, 32'sd899657, -32'sd1201128, -32'sd813849, -32'sd435581, 32'sd178119, 32'sd292209, -32'sd1887012, -32'sd2915813, -32'sd1350723, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1962684, -32'sd3230298, -32'sd2667233, -32'sd1014444, -32'sd378786, -32'sd2254052, -32'sd1908388, -32'sd832257, 32'sd637913, 32'sd42092, 32'sd2255985, 32'sd1641499, -32'sd2068573, -32'sd274776, -32'sd183186, 32'sd1404612, 32'sd178989, -32'sd2018878, -32'sd2865685, -32'sd2607106, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1775267, 32'sd1542547, -32'sd1790775, 32'sd42696, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1980014, -32'sd852993, -32'sd274042, -32'sd233134, 32'sd207949, 32'sd747153, -32'sd577373, -32'sd206621, 32'sd913461, 32'sd2441182, -32'sd518342, 32'sd1084014, 32'sd553782, 32'sd1132199, 32'sd587438, 32'sd4015799, 32'sd2114690, 32'sd2098230, 32'sd237534, 32'sd547365, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2737547, 32'sd176838, 32'sd1046565, -32'sd264541, 32'sd374811, 32'sd179684, 32'sd1681088, 32'sd636085, 32'sd373403, 32'sd3082773, 32'sd1116458, -32'sd392271, 32'sd1306765, 32'sd2874664, -32'sd659312, 32'sd2867950, -32'sd892421, 32'sd3773353, -32'sd358112, -32'sd366835, 32'sd277814, 32'sd794427, 32'sd2881974, 32'sd803973, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1096574, 32'sd821182, 32'sd169513, 32'sd946597, 32'sd48010, 32'sd840379, 32'sd2781214, 32'sd1308203, 32'sd2199151, 32'sd915329, 32'sd221836, 32'sd806345, 32'sd165513, -32'sd276976, -32'sd1683024, 32'sd797221, -32'sd2520242, 32'sd1802340, 32'sd788999, 32'sd692398, 32'sd50392, -32'sd348178, -32'sd558541, -32'sd534942, 32'sd1307363, 32'sd0, 32'sd0, 32'sd67697, 32'sd1203893, -32'sd540468, 32'sd766086, 32'sd294154, 32'sd395378, 32'sd482702, 32'sd1032385, 32'sd897928, 32'sd2396519, -32'sd931578, 32'sd287327, -32'sd514266, -32'sd353303, -32'sd821166, -32'sd999851, -32'sd922128, -32'sd1245913, -32'sd1081720, -32'sd1166845, 32'sd233937, -32'sd1115571, -32'sd2535366, -32'sd2597792, -32'sd827694, -32'sd1459554, 32'sd1033667, 32'sd0, 32'sd2125935, 32'sd1470661, 32'sd1043674, 32'sd600029, -32'sd2434771, 32'sd642884, 32'sd225371, 32'sd2715, 32'sd264303, -32'sd1515263, 32'sd1315752, -32'sd556489, 32'sd1157510, 32'sd1721307, 32'sd2496887, -32'sd360154, -32'sd316267, 32'sd65745, 32'sd150663, -32'sd3233338, -32'sd794450, -32'sd2253174, -32'sd2209317, 32'sd55439, 32'sd728319, -32'sd351497, 32'sd1195889, 32'sd0, 32'sd1442037, 32'sd444712, -32'sd853978, -32'sd123117, -32'sd463950, -32'sd685071, -32'sd1492093, 32'sd162639, -32'sd436745, -32'sd100553, 32'sd2960211, -32'sd530079, -32'sd92378, -32'sd72935, 32'sd1506357, -32'sd1532400, -32'sd914920, 32'sd662621, -32'sd3165580, -32'sd1588405, 32'sd35595, -32'sd1344349, -32'sd2259632, -32'sd40959, -32'sd1714579, 32'sd1467524, -32'sd121447, 32'sd2096125, 32'sd619810, -32'sd560952, -32'sd1187637, 32'sd1565936, 32'sd2258996, 32'sd739948, 32'sd1819455, -32'sd1532109, -32'sd1026752, 32'sd1300648, 32'sd585304, 32'sd344192, 32'sd252374, -32'sd1619115, 32'sd1198544, -32'sd3128715, -32'sd1489760, -32'sd2300837, -32'sd3482704, -32'sd2459968, -32'sd3222304, -32'sd2529945, -32'sd2638491, -32'sd431248, -32'sd1441115, -32'sd397186, -32'sd81542, 32'sd1547646, 32'sd2929705, 32'sd1623696, -32'sd243194, 32'sd317019, -32'sd569813, -32'sd605637, 32'sd224904, 32'sd364350, -32'sd4193516, 32'sd1631200, -32'sd287161, -32'sd247653, 32'sd1888887, -32'sd210847, -32'sd33886, -32'sd469004, -32'sd4038340, -32'sd3560778, -32'sd4678919, -32'sd3298968, -32'sd1178235, -32'sd2602832, -32'sd2835089, -32'sd1380127, -32'sd2644287, 32'sd170955, -32'sd2663775, -32'sd909565, -32'sd1448858, -32'sd1474247, -32'sd425905, 32'sd557683, 32'sd1502040, -32'sd389817, 32'sd1469828, -32'sd799428, -32'sd2424330, -32'sd1820199, -32'sd859469, 32'sd873537, 32'sd4239323, 32'sd3579516, -32'sd1446161, -32'sd2392781, -32'sd4122072, -32'sd3121009, -32'sd5054799, -32'sd654204, -32'sd929240, -32'sd1576250, -32'sd980658, 32'sd90004, -32'sd2582125, -32'sd2443373, 32'sd1359859, 32'sd882087, -32'sd949027, -32'sd1127893, -32'sd2753451, -32'sd2746643, -32'sd989708, -32'sd416377, -32'sd650671, -32'sd21525, 32'sd949160, 32'sd2438650, 32'sd2088328, 32'sd3138376, 32'sd6374408, 32'sd756356, -32'sd5240028, -32'sd3955977, -32'sd1071271, -32'sd1677273, -32'sd2919543, -32'sd1032490, -32'sd1030699, 32'sd1338767, 32'sd495035, 32'sd84864, 32'sd637824, 32'sd218785, -32'sd193911, 32'sd787120, 32'sd2849888, 32'sd1377397, 32'sd3170408, -32'sd442268, -32'sd36672, -32'sd1597271, -32'sd1369973, 32'sd2348351, 32'sd957734, 32'sd1754086, 32'sd2565777, 32'sd3238746, 32'sd721671, -32'sd2190916, -32'sd4141531, -32'sd1266003, 32'sd893231, -32'sd1883377, -32'sd1982199, -32'sd196271, 32'sd349597, -32'sd551054, 32'sd80435, -32'sd1013092, -32'sd341511, -32'sd1253316, -32'sd1908319, -32'sd853611, 32'sd532419, 32'sd154913, -32'sd104464, -32'sd1435466, 32'sd1016864, 32'sd1129542, 32'sd1679440, 32'sd71045, 32'sd3986311, 32'sd2179861, 32'sd2549523, 32'sd635408, -32'sd2229662, -32'sd526224, -32'sd123381, -32'sd462835, -32'sd1078262, 32'sd1502381, 32'sd199999, -32'sd847902, -32'sd690731, 32'sd1081941, 32'sd1022850, 32'sd542242, -32'sd1110120, -32'sd2233734, 32'sd875192, 32'sd642522, 32'sd1470192, -32'sd118535, 32'sd761603, -32'sd438391, 32'sd844714, 32'sd3579746, 32'sd3268873, 32'sd1336493, 32'sd2005381, 32'sd2911690, -32'sd1281754, -32'sd1003493, -32'sd2869200, -32'sd1960254, -32'sd1359545, -32'sd776723, -32'sd778538, -32'sd1884513, -32'sd87930, -32'sd818648, 32'sd1038347, -32'sd22935, 32'sd3840286, -32'sd511350, 32'sd579913, -32'sd1805013, -32'sd417447, -32'sd433385, 32'sd211840, -32'sd1780304, -32'sd1037995, -32'sd1803155, 32'sd1555220, 32'sd614196, 32'sd1831552, 32'sd2463986, 32'sd1113319, 32'sd671534, -32'sd1732920, -32'sd130314, -32'sd560593, -32'sd900822, 32'sd308690, -32'sd1182661, -32'sd2831209, 32'sd700475, -32'sd960529, 32'sd1052399, 32'sd462104, 32'sd1303187, 32'sd1965250, 32'sd1299364, 32'sd208530, -32'sd1308172, -32'sd120701, 32'sd215700, -32'sd207082, -32'sd128471, -32'sd558016, 32'sd28692, 32'sd974945, 32'sd561788, 32'sd2608847, 32'sd1880977, -32'sd1772506, 32'sd152046, -32'sd1098159, -32'sd290696, -32'sd2281089, 32'sd512435, -32'sd1331100, -32'sd903366, -32'sd2187131, -32'sd9114, -32'sd647935, 32'sd3128425, 32'sd1288483, 32'sd1602243, 32'sd1725942, -32'sd301462, -32'sd624307, -32'sd3287949, -32'sd1456418, -32'sd44352, 32'sd1510127, 32'sd379579, 32'sd843342, 32'sd265409, -32'sd155357, 32'sd255612, 32'sd1445879, 32'sd3453479, 32'sd1528835, 32'sd562819, 32'sd652768, -32'sd2673939, -32'sd3236379, 32'sd11185, -32'sd1555038, -32'sd1724030, -32'sd3755315, -32'sd820743, -32'sd1913170, 32'sd139981, -32'sd1600829, -32'sd117986, -32'sd368313, 32'sd1815877, 32'sd103287, -32'sd583706, 32'sd143507, 32'sd0, 32'sd468132, -32'sd704594, 32'sd743955, -32'sd294156, 32'sd867435, -32'sd1587604, 32'sd2080165, 32'sd2297691, 32'sd1847848, 32'sd1281017, 32'sd521165, -32'sd861164, -32'sd2351778, -32'sd948946, -32'sd4813524, 32'sd560351, 32'sd139819, 32'sd792449, -32'sd145374, -32'sd577403, 32'sd440840, 32'sd454991, -32'sd19492, -32'sd1638441, -32'sd1228020, -32'sd1682352, 32'sd742174, 32'sd40164, -32'sd1253414, -32'sd477755, 32'sd94483, 32'sd1161968, 32'sd432857, -32'sd1655139, 32'sd1314136, 32'sd1535278, 32'sd3636445, 32'sd2962775, 32'sd768743, 32'sd1145664, -32'sd2375760, -32'sd2510364, -32'sd306611, 32'sd74309, 32'sd2289018, -32'sd1588537, -32'sd1002770, -32'sd498121, 32'sd136034, 32'sd1344406, -32'sd1106606, -32'sd2068840, 32'sd255450, -32'sd1286992, -32'sd564945, 32'sd1005437, 32'sd860191, -32'sd693122, -32'sd1780921, 32'sd2166804, -32'sd508943, -32'sd1895532, -32'sd2394144, -32'sd1274040, 32'sd1030196, 32'sd2566587, 32'sd4012205, 32'sd3738181, -32'sd1318975, 32'sd2578948, -32'sd845615, -32'sd575384, -32'sd412162, 32'sd220333, 32'sd933768, 32'sd1313171, -32'sd207134, 32'sd1018559, 32'sd1057409, -32'sd1794670, -32'sd2537779, -32'sd1582875, -32'sd262610, 32'sd0, 32'sd1332875, -32'sd1344179, -32'sd1893004, -32'sd662518, -32'sd644976, -32'sd4084088, -32'sd1411382, -32'sd996295, 32'sd273962, -32'sd630719, 32'sd493848, 32'sd957832, 32'sd1469219, 32'sd3973577, 32'sd4024125, 32'sd1700451, -32'sd100809, 32'sd1142048, -32'sd1649713, 32'sd381781, -32'sd36131, 32'sd282671, -32'sd354756, 32'sd1617881, 32'sd442109, -32'sd991648, 32'sd730447, -32'sd1081299, -32'sd63414, 32'sd1765275, -32'sd1303237, -32'sd781280, -32'sd2641190, -32'sd1082361, -32'sd240476, 32'sd755718, 32'sd526912, 32'sd747771, 32'sd89569, -32'sd514311, 32'sd771141, 32'sd2870127, 32'sd3756624, 32'sd2657018, -32'sd1067685, 32'sd1498114, -32'sd382165, -32'sd343089, 32'sd540778, 32'sd1391823, -32'sd257839, -32'sd3609089, -32'sd1874029, 32'sd2535112, -32'sd234251, 32'sd1122320, 32'sd2104366, 32'sd1142903, 32'sd26244, 32'sd1646964, -32'sd1760143, -32'sd190388, -32'sd1316275, 32'sd1514793, 32'sd428470, -32'sd838714, -32'sd889746, 32'sd1115846, 32'sd648743, 32'sd68986, 32'sd1987771, 32'sd2272047, 32'sd916018, -32'sd224973, -32'sd1151682, 32'sd719086, 32'sd1120458, 32'sd843407, -32'sd94541, -32'sd2254239, -32'sd912745, 32'sd1171675, 32'sd1405373, 32'sd0, 32'sd1637048, 32'sd1602059, -32'sd815222, 32'sd1471156, -32'sd1612526, -32'sd2737030, -32'sd1180646, -32'sd3393276, 32'sd843686, -32'sd89902, -32'sd486787, -32'sd140035, -32'sd404867, 32'sd1491623, 32'sd1713775, -32'sd112019, 32'sd2972217, 32'sd650985, 32'sd618611, -32'sd640882, -32'sd2223979, -32'sd200896, -32'sd1360645, -32'sd1493903, 32'sd1224435, -32'sd454685, 32'sd0, 32'sd0, 32'sd0, 32'sd2082412, -32'sd1239489, 32'sd1092888, 32'sd303650, -32'sd1097188, 32'sd926283, 32'sd44775, 32'sd226680, 32'sd875310, -32'sd1669854, 32'sd1866502, 32'sd164309, -32'sd35837, 32'sd928910, 32'sd2293128, 32'sd2135331, 32'sd1157536, -32'sd390777, -32'sd1833158, -32'sd771793, 32'sd438178, 32'sd396323, 32'sd1878943, -32'sd1652855, -32'sd1148663, 32'sd0, 32'sd0, 32'sd0, -32'sd573215, 32'sd1083522, -32'sd670341, -32'sd1096563, -32'sd1197781, 32'sd3204150, 32'sd76915, -32'sd2252787, -32'sd3759907, -32'sd4676709, 32'sd736929, 32'sd1603153, 32'sd135202, -32'sd799678, 32'sd607637, -32'sd981943, 32'sd137229, 32'sd3188971, -32'sd2262758, 32'sd103836, 32'sd3535103, -32'sd1849254, -32'sd2150824, 32'sd775146, 32'sd965864, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1906372, -32'sd244617, -32'sd302753, 32'sd1051186, -32'sd127494, 32'sd1090427, -32'sd1306126, -32'sd563504, 32'sd89564, 32'sd1427887, 32'sd151534, 32'sd210347, 32'sd2291482, 32'sd1688447, 32'sd1632964, 32'sd305025, 32'sd1068268, -32'sd1120873, -32'sd2408484, -32'sd250315, -32'sd1114869, 32'sd574548, 32'sd1055030, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd727443, -32'sd1410740, 32'sd299264, -32'sd1300345, 32'sd864919, 32'sd693843, 32'sd1791282, -32'sd923069, 32'sd2189822, 32'sd669577, -32'sd1966643, -32'sd3647252, 32'sd919858, 32'sd65792, -32'sd765792, -32'sd386281, 32'sd1009545, 32'sd260394, -32'sd949080, -32'sd204503, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd267693, 32'sd9592, -32'sd300679, -32'sd1538392, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd926650, -32'sd1591634, -32'sd1341900, -32'sd852284, 32'sd85719, -32'sd674764, -32'sd274419, 32'sd816795, 32'sd786909, 32'sd1039982, 32'sd707355, -32'sd1447086, -32'sd304691, 32'sd202586, 32'sd2516049, 32'sd1363316, 32'sd440249, -32'sd627227, -32'sd1212914, -32'sd649915, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd276223, -32'sd1101588, -32'sd198673, -32'sd1432307, -32'sd654845, -32'sd217922, 32'sd1088497, 32'sd882817, 32'sd2853801, 32'sd1585246, 32'sd1756589, 32'sd1029071, -32'sd1641808, 32'sd888245, 32'sd1693266, 32'sd669995, 32'sd1849039, 32'sd1854899, 32'sd2119490, 32'sd3469148, 32'sd1570509, 32'sd599816, 32'sd3049446, 32'sd539451, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd322177, 32'sd1010325, -32'sd792006, 32'sd1183947, -32'sd335820, -32'sd423054, 32'sd1295745, 32'sd497787, -32'sd655995, -32'sd756863, -32'sd1066751, 32'sd326553, 32'sd964597, -32'sd716075, 32'sd2600261, -32'sd435195, -32'sd602698, -32'sd981139, 32'sd60307, 32'sd132799, 32'sd239106, 32'sd3515929, -32'sd21547, -32'sd577695, 32'sd1535801, 32'sd0, 32'sd0, -32'sd539720, 32'sd640232, 32'sd301268, 32'sd367151, 32'sd505195, -32'sd1216596, -32'sd2050383, 32'sd606471, -32'sd2042307, -32'sd323558, 32'sd966692, 32'sd229316, 32'sd289031, 32'sd480414, 32'sd31394, -32'sd1069241, 32'sd526996, 32'sd1029745, 32'sd1907830, 32'sd2520548, 32'sd359675, 32'sd1515676, 32'sd1442694, 32'sd689737, -32'sd942268, -32'sd280622, -32'sd817655, 32'sd0, -32'sd221325, 32'sd854518, 32'sd1380313, -32'sd1308430, -32'sd2242941, -32'sd76639, -32'sd2056828, -32'sd1658823, -32'sd3234622, 32'sd554451, 32'sd90475, -32'sd3355474, 32'sd664846, 32'sd1637912, -32'sd753428, -32'sd3154490, 32'sd637498, 32'sd1157167, 32'sd1479560, -32'sd863068, 32'sd851427, 32'sd747669, 32'sd1573040, 32'sd279287, 32'sd1627607, 32'sd138356, -32'sd1408903, 32'sd0, -32'sd945588, -32'sd1455374, 32'sd782550, 32'sd315980, -32'sd3230992, -32'sd980034, -32'sd251717, 32'sd1152827, -32'sd4373975, 32'sd981548, 32'sd1423012, 32'sd304911, 32'sd1798018, -32'sd1737069, 32'sd3458678, -32'sd1237223, -32'sd671539, -32'sd161166, -32'sd1184237, -32'sd2590507, 32'sd80661, 32'sd1878201, 32'sd227829, -32'sd120576, 32'sd225428, -32'sd290921, 32'sd2226012, 32'sd92927, 32'sd261387, -32'sd408001, -32'sd795948, -32'sd473843, -32'sd749703, -32'sd489049, -32'sd1802395, -32'sd3716286, 32'sd302968, 32'sd514469, 32'sd1816686, 32'sd288172, 32'sd1941601, 32'sd118727, 32'sd1321945, -32'sd1246063, 32'sd201665, 32'sd2258974, 32'sd693836, -32'sd1695653, 32'sd179540, 32'sd477938, 32'sd1347466, 32'sd670286, 32'sd183802, 32'sd160692, -32'sd567284, 32'sd1338706, 32'sd58456, 32'sd1692189, -32'sd839137, -32'sd709467, -32'sd1658203, -32'sd1926871, -32'sd549797, -32'sd1000464, -32'sd670682, -32'sd423459, 32'sd1904241, 32'sd1862277, 32'sd1286350, -32'sd943710, -32'sd805762, 32'sd1501390, -32'sd273780, 32'sd1424656, 32'sd1465723, -32'sd180235, 32'sd642837, -32'sd738942, -32'sd1586174, 32'sd1388568, -32'sd41356, 32'sd237266, -32'sd1050550, -32'sd1555540, -32'sd989355, -32'sd530405, -32'sd1064825, 32'sd2714307, -32'sd1018945, -32'sd980845, 32'sd611883, -32'sd1463315, -32'sd1557062, 32'sd251202, 32'sd1056540, -32'sd2075227, 32'sd290441, 32'sd643419, -32'sd2711463, -32'sd895935, 32'sd1673182, 32'sd1249647, 32'sd1385407, 32'sd1234388, -32'sd118718, -32'sd891092, -32'sd1448037, 32'sd942605, 32'sd485131, 32'sd1381454, -32'sd3013550, 32'sd523152, -32'sd1722375, 32'sd645079, 32'sd3335161, 32'sd691926, 32'sd1738872, 32'sd227248, 32'sd154870, -32'sd1155869, -32'sd986795, -32'sd1579494, -32'sd659061, 32'sd141266, 32'sd331334, 32'sd2077109, -32'sd1725721, -32'sd2679787, 32'sd3257018, 32'sd2682262, 32'sd222204, -32'sd1981404, -32'sd1446185, 32'sd2224070, 32'sd1017171, -32'sd1124682, -32'sd1356058, 32'sd755151, -32'sd1092423, 32'sd871391, 32'sd4469983, -32'sd4777810, 32'sd1480889, -32'sd3982395, -32'sd2092999, -32'sd213428, 32'sd1160212, -32'sd1874199, -32'sd575528, -32'sd1863768, -32'sd1124400, -32'sd827819, 32'sd2262709, 32'sd856084, -32'sd2111400, -32'sd5044752, -32'sd1122300, 32'sd1220841, -32'sd338232, -32'sd92485, 32'sd145118, -32'sd11391, 32'sd270379, 32'sd793719, 32'sd342731, 32'sd1093030, 32'sd2001038, 32'sd568048, -32'sd291725, -32'sd778099, -32'sd4048489, -32'sd884544, -32'sd1871568, -32'sd256002, -32'sd793635, -32'sd2142415, 32'sd205618, -32'sd604469, -32'sd393885, 32'sd2578601, 32'sd4957472, 32'sd1499888, -32'sd2772545, -32'sd3333590, 32'sd2080719, -32'sd75668, 32'sd175297, 32'sd1158236, -32'sd824821, -32'sd789250, 32'sd1729756, 32'sd1043341, -32'sd1422642, 32'sd267538, -32'sd227051, -32'sd608813, 32'sd1311298, 32'sd1520363, -32'sd2932269, 32'sd136377, -32'sd1630346, -32'sd193818, -32'sd855534, 32'sd530136, 32'sd2727879, -32'sd506770, 32'sd2953495, 32'sd2440157, 32'sd1365236, 32'sd319529, -32'sd3116543, -32'sd2221643, -32'sd1226777, 32'sd1321532, -32'sd1675491, 32'sd259995, -32'sd453172, 32'sd717494, 32'sd1937878, -32'sd121904, -32'sd348474, 32'sd1309348, -32'sd433369, -32'sd1298374, -32'sd149316, 32'sd502893, -32'sd843548, 32'sd79757, 32'sd2422780, 32'sd126210, 32'sd2292729, -32'sd104231, 32'sd3608039, 32'sd2248234, 32'sd2982221, 32'sd4871916, 32'sd486359, -32'sd2004031, -32'sd2753966, -32'sd2894180, -32'sd1685898, -32'sd572789, -32'sd47926, -32'sd658308, 32'sd321517, -32'sd984584, 32'sd564891, 32'sd619571, -32'sd1858011, -32'sd1463057, -32'sd1553835, -32'sd1260991, 32'sd395497, -32'sd506367, 32'sd1237587, 32'sd1277484, 32'sd1752007, 32'sd858463, 32'sd2362764, 32'sd888887, 32'sd2942618, 32'sd4105466, 32'sd3728407, 32'sd3818826, -32'sd4774017, -32'sd3872639, -32'sd4530983, -32'sd1228763, -32'sd595626, 32'sd268835, 32'sd670693, 32'sd275084, 32'sd146079, -32'sd604711, 32'sd439839, 32'sd501150, 32'sd12529, -32'sd3269258, 32'sd29187, -32'sd1305637, -32'sd90249, -32'sd1879633, 32'sd1336017, 32'sd331215, 32'sd1696072, 32'sd1893674, 32'sd3632638, 32'sd3091901, 32'sd2800448, 32'sd4479506, 32'sd6916529, -32'sd565327, -32'sd6683495, -32'sd3794072, -32'sd2543564, -32'sd956780, -32'sd1060331, -32'sd1879189, 32'sd915543, 32'sd249078, 32'sd1087137, 32'sd303134, -32'sd2639013, -32'sd1115927, -32'sd567945, 32'sd704243, 32'sd935467, 32'sd0, -32'sd26324, -32'sd2629267, -32'sd159937, 32'sd3008231, 32'sd2359310, 32'sd1631021, 32'sd1685395, 32'sd2088645, 32'sd3610784, 32'sd6249588, 32'sd4082162, -32'sd4663721, -32'sd7039069, 32'sd437297, -32'sd1376507, -32'sd2067587, -32'sd298167, -32'sd20318, 32'sd1454571, 32'sd389101, 32'sd1236469, 32'sd822440, -32'sd469098, 32'sd813073, -32'sd315504, 32'sd556684, 32'sd12335, -32'sd138004, -32'sd582639, -32'sd2612700, 32'sd666029, 32'sd64423, 32'sd83135, 32'sd408697, 32'sd2259370, 32'sd2776121, 32'sd5764761, 32'sd4066943, 32'sd2190141, -32'sd5365881, -32'sd6897172, -32'sd867005, -32'sd688185, -32'sd2171854, -32'sd151270, 32'sd1798249, -32'sd1544923, -32'sd721273, -32'sd274051, 32'sd280884, 32'sd1384519, 32'sd158759, 32'sd541614, 32'sd924737, 32'sd695612, -32'sd1026409, -32'sd493844, -32'sd2093361, 32'sd901809, 32'sd726371, -32'sd909429, -32'sd838090, 32'sd229469, 32'sd2502153, 32'sd3928977, 32'sd5179565, -32'sd2045061, -32'sd4653657, -32'sd3646336, -32'sd1835867, -32'sd2907750, -32'sd2097895, 32'sd1084486, -32'sd609677, -32'sd1044429, -32'sd1052769, -32'sd276017, 32'sd385297, -32'sd868512, -32'sd734709, -32'sd987691, -32'sd19482, 32'sd568162, 32'sd0, 32'sd1317229, -32'sd1140538, -32'sd1526350, -32'sd516856, 32'sd732822, -32'sd308151, 32'sd3451932, 32'sd1902853, 32'sd3425825, 32'sd4308299, -32'sd3706075, -32'sd2001461, -32'sd2138441, -32'sd1968255, -32'sd3422805, -32'sd4815465, -32'sd3373534, -32'sd1484333, -32'sd1371897, -32'sd147444, 32'sd498513, 32'sd862661, -32'sd612952, -32'sd1340890, -32'sd1237822, -32'sd2914430, -32'sd1340652, 32'sd676399, -32'sd1730112, 32'sd1029845, 32'sd3532415, -32'sd804326, 32'sd49920, 32'sd1191397, 32'sd4804651, 32'sd1410460, 32'sd2041790, 32'sd408815, 32'sd2584632, 32'sd641506, -32'sd1531205, -32'sd934264, -32'sd1823343, -32'sd2705187, -32'sd1852056, -32'sd3526519, -32'sd1559785, 32'sd74542, 32'sd1078664, -32'sd896269, -32'sd697417, -32'sd3052341, -32'sd2678270, 32'sd717888, -32'sd85160, -32'sd280693, 32'sd312513, -32'sd192043, 32'sd999391, 32'sd774205, -32'sd349673, 32'sd1134470, 32'sd2392808, 32'sd637049, -32'sd319801, 32'sd1305039, 32'sd1466944, 32'sd3446021, 32'sd3421185, -32'sd1934840, -32'sd236190, -32'sd2090486, -32'sd2387836, -32'sd3179341, -32'sd1402787, -32'sd1209170, 32'sd795849, 32'sd860738, -32'sd2365639, -32'sd2126592, -32'sd3381350, 32'sd1260430, 32'sd1407546, 32'sd0, -32'sd1212058, 32'sd117626, -32'sd996439, -32'sd1591142, -32'sd1070331, 32'sd1114160, 32'sd2348334, 32'sd3268963, -32'sd1197868, 32'sd2084292, 32'sd2130847, 32'sd735196, 32'sd1191809, -32'sd122909, -32'sd2269840, -32'sd479214, -32'sd1361244, -32'sd2129043, 32'sd794638, -32'sd936006, -32'sd64526, -32'sd3112394, 32'sd815406, 32'sd593453, 32'sd1684805, -32'sd393858, 32'sd0, 32'sd0, 32'sd0, -32'sd908613, -32'sd1211431, 32'sd527489, 32'sd1750782, -32'sd707984, 32'sd178715, 32'sd2075605, -32'sd429731, -32'sd1968930, -32'sd1369439, 32'sd959924, 32'sd933739, -32'sd992677, -32'sd1584058, 32'sd69434, -32'sd1769509, -32'sd1230467, -32'sd692759, -32'sd696327, -32'sd2409764, -32'sd2036486, 32'sd283242, -32'sd1945219, 32'sd40773, -32'sd181103, 32'sd0, 32'sd0, 32'sd0, -32'sd267101, -32'sd943197, 32'sd148122, -32'sd1713554, -32'sd925626, -32'sd97788, 32'sd1501498, -32'sd1504667, -32'sd327421, 32'sd124167, -32'sd3584578, -32'sd836612, 32'sd399665, -32'sd467759, 32'sd93268, -32'sd2034019, -32'sd2818874, -32'sd1906380, -32'sd2135140, -32'sd524223, 32'sd660494, -32'sd966575, -32'sd1648841, 32'sd784318, -32'sd1238222, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1028948, 32'sd328390, -32'sd407689, -32'sd2563673, -32'sd2739259, -32'sd2379444, -32'sd2595289, -32'sd776368, -32'sd1155628, -32'sd2405281, -32'sd76734, -32'sd3845154, -32'sd3049625, -32'sd1072938, -32'sd2572467, 32'sd157338, -32'sd1096428, -32'sd2094796, -32'sd2926751, -32'sd1123937, -32'sd1022163, 32'sd834403, -32'sd1375419, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1460541, 32'sd391376, 32'sd201920, -32'sd117483, 32'sd180282, -32'sd484654, -32'sd735437, -32'sd1003471, 32'sd1103697, -32'sd960036, -32'sd813808, -32'sd223666, -32'sd259370, -32'sd1022096, -32'sd1073731, 32'sd474726, -32'sd1442221, -32'sd1279253, 32'sd690121, -32'sd1155252, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd7895146, -32'sd9704588, -32'sd7949293, -32'sd6989737, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd7180807, -32'sd8856438, -32'sd9148076, -32'sd7723454, -32'sd9193642, -32'sd9591848, -32'sd9140037, -32'sd10159779, -32'sd10041719, -32'sd7223934, -32'sd4717022, -32'sd9443394, -32'sd9041309, -32'sd9752799, -32'sd9029863, -32'sd9947937, -32'sd9529797, -32'sd7838457, -32'sd8822004, -32'sd9386715, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd7497057, -32'sd9400555, 32'sd1309132, -32'sd2760510, -32'sd8082768, -32'sd8559503, -32'sd10015076, -32'sd4525801, -32'sd5435427, -32'sd9670835, -32'sd7888445, -32'sd7600493, -32'sd8766672, -32'sd7798782, -32'sd7581775, -32'sd3811269, -32'sd2224962, -32'sd6913606, -32'sd3521903, -32'sd1617504, -32'sd2859942, -32'sd6680589, -32'sd7584858, -32'sd8177769, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd8957603, -32'sd2449304, -32'sd2641155, -32'sd7051125, -32'sd7781754, -32'sd6440077, -32'sd3280717, -32'sd2510076, -32'sd4136000, -32'sd4554706, -32'sd8829726, -32'sd5968515, -32'sd5463834, -32'sd1074063, 32'sd1864568, 32'sd2417654, 32'sd835255, -32'sd1569484, 32'sd573878, -32'sd622835, 32'sd569676, 32'sd2982699, -32'sd721614, -32'sd626460, -32'sd1318783, 32'sd0, 32'sd0, -32'sd7510727, -32'sd586171, 32'sd1929557, -32'sd2867700, -32'sd2556528, 32'sd834824, 32'sd2032702, 32'sd343796, 32'sd392246, -32'sd437694, -32'sd965512, 32'sd787073, 32'sd374527, 32'sd218172, -32'sd388276, 32'sd266428, 32'sd1934630, 32'sd1360670, -32'sd474062, -32'sd872035, -32'sd1009811, -32'sd179669, -32'sd265494, 32'sd1656150, -32'sd156324, -32'sd12177, -32'sd8776996, 32'sd0, -32'sd7661669, -32'sd230647, -32'sd12420, -32'sd879654, -32'sd1133131, 32'sd251238, 32'sd1479960, -32'sd1553949, -32'sd1462462, 32'sd289367, 32'sd3717277, 32'sd5918643, 32'sd3432589, 32'sd1957656, 32'sd307169, 32'sd2316220, 32'sd3473355, 32'sd2324168, -32'sd8011, 32'sd1926634, 32'sd654391, -32'sd658890, -32'sd1817860, -32'sd1209884, 32'sd1690625, 32'sd315823, 32'sd746262, 32'sd0, -32'sd8827805, -32'sd1867294, -32'sd427481, -32'sd245879, -32'sd790202, -32'sd1427792, -32'sd1097146, -32'sd627665, -32'sd462891, 32'sd254501, 32'sd3202202, 32'sd2281394, 32'sd2256068, 32'sd1960797, 32'sd5011772, 32'sd2301853, 32'sd3523010, 32'sd1911210, 32'sd2275153, 32'sd516966, -32'sd288325, -32'sd737279, -32'sd212551, -32'sd391139, 32'sd935906, -32'sd1824422, 32'sd283457, -32'sd7934077, -32'sd8363785, -32'sd1616453, -32'sd936944, 32'sd1163324, 32'sd983468, 32'sd497438, -32'sd864524, 32'sd1512451, 32'sd3589682, 32'sd1705329, 32'sd67434, -32'sd185866, 32'sd1293068, 32'sd770123, 32'sd3047690, 32'sd1478452, 32'sd1742758, 32'sd3150236, 32'sd303786, 32'sd749643, 32'sd2341236, 32'sd986411, -32'sd1039991, 32'sd2143083, 32'sd1765278, 32'sd164971, 32'sd681427, -32'sd508326, -32'sd7568839, -32'sd341183, 32'sd1551204, 32'sd1689136, 32'sd1580581, 32'sd3233236, 32'sd2444825, -32'sd218131, 32'sd1769786, 32'sd1453204, -32'sd779187, 32'sd874146, 32'sd2269507, 32'sd1519189, -32'sd420298, 32'sd2808088, 32'sd2281746, 32'sd3438321, 32'sd2850334, -32'sd117716, -32'sd585762, 32'sd105668, -32'sd1603273, 32'sd839934, 32'sd404138, 32'sd208001, 32'sd804410, -32'sd8644518, -32'sd8420694, -32'sd829483, 32'sd933050, -32'sd692374, 32'sd3346098, 32'sd1369384, 32'sd619524, 32'sd967650, -32'sd190408, 32'sd1630829, -32'sd1233490, -32'sd1132631, 32'sd3083370, 32'sd96807, -32'sd687678, -32'sd3734406, -32'sd943389, -32'sd1239243, 32'sd992855, -32'sd36838, 32'sd286623, 32'sd453163, 32'sd1953114, -32'sd1373745, 32'sd410070, 32'sd1693518, -32'sd3675409, -32'sd9493654, -32'sd6168966, -32'sd2117868, -32'sd113636, 32'sd1105143, 32'sd679321, 32'sd2761009, 32'sd1124555, 32'sd324537, 32'sd3470821, 32'sd1492386, -32'sd1129845, 32'sd950155, -32'sd1325782, 32'sd28962, -32'sd5448650, -32'sd4340986, -32'sd2004824, 32'sd2324911, 32'sd2133161, 32'sd3410199, 32'sd2738218, 32'sd4849361, 32'sd1446918, -32'sd1567570, -32'sd2310750, 32'sd703814, -32'sd9675802, -32'sd9276492, -32'sd1893490, -32'sd1557033, 32'sd740704, 32'sd2327048, 32'sd1751123, 32'sd612257, -32'sd1154644, -32'sd442950, -32'sd1263410, 32'sd1157808, -32'sd105303, 32'sd1050821, 32'sd1318651, 32'sd3394798, 32'sd543029, 32'sd854707, 32'sd1958801, 32'sd1980916, 32'sd1209306, 32'sd367338, -32'sd1377983, -32'sd858998, 32'sd1129731, 32'sd2001611, 32'sd1536222, 32'sd856668, -32'sd1701638, -32'sd2569804, -32'sd2937190, -32'sd2432313, 32'sd225012, 32'sd1277866, 32'sd455135, -32'sd1635591, 32'sd1906160, -32'sd153910, 32'sd240034, 32'sd133148, 32'sd661205, -32'sd1938172, 32'sd2143403, 32'sd2982592, 32'sd1522710, 32'sd884336, 32'sd1482057, -32'sd387200, -32'sd24514, 32'sd2501, 32'sd1176967, 32'sd139047, -32'sd1732128, -32'sd2272916, -32'sd306850, 32'sd16621, 32'sd1210908, -32'sd7735294, -32'sd6988294, -32'sd1942593, 32'sd49933, -32'sd889212, 32'sd38771, -32'sd31420, 32'sd2336739, -32'sd879753, 32'sd1016459, -32'sd502709, 32'sd1578129, -32'sd1330173, 32'sd2088635, 32'sd2574257, 32'sd564439, 32'sd989043, -32'sd1592855, 32'sd1215928, -32'sd1962801, -32'sd737447, -32'sd2956035, -32'sd2027915, -32'sd404550, -32'sd670660, 32'sd289286, 32'sd1733231, 32'sd281875, -32'sd9060344, -32'sd9075244, -32'sd1528282, -32'sd4456502, 32'sd1376773, 32'sd1323112, 32'sd841505, -32'sd2045230, -32'sd459585, -32'sd1856386, -32'sd673768, -32'sd66859, -32'sd2303117, 32'sd2649120, 32'sd3057451, 32'sd863738, -32'sd1206928, 32'sd726937, -32'sd970038, -32'sd3668967, -32'sd2655648, -32'sd3995716, -32'sd4035602, -32'sd3132425, -32'sd2990390, 32'sd503944, 32'sd951090, -32'sd7374125, -32'sd9170142, -32'sd7491634, -32'sd1710892, -32'sd1997135, -32'sd2428280, -32'sd3242700, 32'sd1248021, -32'sd107199, -32'sd1356365, 32'sd616727, -32'sd962269, 32'sd126795, 32'sd908852, 32'sd2469240, 32'sd3016030, 32'sd2351676, -32'sd1635647, 32'sd185641, -32'sd2520918, -32'sd1484532, -32'sd2307199, -32'sd3429380, -32'sd657662, -32'sd570027, 32'sd1517154, 32'sd2463504, -32'sd4907047, -32'sd1879944, -32'sd8479170, -32'sd9029991, -32'sd3885123, -32'sd2383210, -32'sd2709066, -32'sd4377568, -32'sd1226777, 32'sd2249175, 32'sd1599690, 32'sd1546144, -32'sd422409, 32'sd102810, 32'sd1413247, -32'sd364505, 32'sd580859, 32'sd358411, 32'sd690087, 32'sd499982, -32'sd2193227, -32'sd3883832, -32'sd2033034, -32'sd2482498, -32'sd613602, 32'sd1217132, 32'sd2365037, 32'sd397610, -32'sd2127444, 32'sd283524, 32'sd0, -32'sd9828797, -32'sd4408629, -32'sd2420878, 32'sd561430, -32'sd2513861, -32'sd2497141, 32'sd725639, 32'sd1372926, 32'sd1705077, -32'sd1569084, 32'sd282191, 32'sd1139027, -32'sd3418624, -32'sd564441, -32'sd2091881, -32'sd579420, -32'sd222732, -32'sd1893887, -32'sd243393, -32'sd2251737, 32'sd552746, 32'sd2942912, 32'sd75274, -32'sd347884, -32'sd2218715, -32'sd1880202, 32'sd261927, -32'sd9098391, -32'sd265942, -32'sd1491966, -32'sd5430286, -32'sd1055982, -32'sd659538, -32'sd305270, -32'sd336901, -32'sd393051, 32'sd129757, -32'sd862522, -32'sd2304671, -32'sd3965575, -32'sd1742926, -32'sd2906778, -32'sd2301600, -32'sd1971995, -32'sd413755, -32'sd476605, 32'sd322272, 32'sd1089490, 32'sd1258765, 32'sd1306235, -32'sd1840609, -32'sd269067, -32'sd2918089, -32'sd3159246, 32'sd237442, -32'sd9410571, 32'sd65653, -32'sd3784295, -32'sd902710, 32'sd2167233, 32'sd2022731, 32'sd168547, -32'sd1052346, -32'sd1083019, -32'sd1146567, -32'sd2040153, -32'sd5003936, -32'sd3834147, -32'sd2915952, -32'sd2892233, -32'sd3255747, -32'sd1567227, -32'sd1272064, 32'sd2034495, 32'sd1014457, 32'sd1046298, -32'sd326632, 32'sd800878, 32'sd1077228, -32'sd1028729, -32'sd5443030, -32'sd2923927, -32'sd9944453, 32'sd0, -32'sd455510, -32'sd3803197, 32'sd1626718, 32'sd1052497, 32'sd2639288, 32'sd2382418, 32'sd423571, -32'sd820876, -32'sd1763571, -32'sd2020148, -32'sd3212865, -32'sd1444988, 32'sd98874, -32'sd1058640, 32'sd526536, -32'sd1850076, -32'sd1244703, -32'sd298048, 32'sd2832818, 32'sd2723707, 32'sd207060, 32'sd392500, -32'sd226354, -32'sd733720, -32'sd3921972, -32'sd2082418, -32'sd9236450, 32'sd427693, -32'sd2531214, -32'sd200601, -32'sd3543335, 32'sd2044742, 32'sd2006168, 32'sd1654724, 32'sd1365592, -32'sd1186339, 32'sd721545, -32'sd26158, -32'sd393547, -32'sd810385, -32'sd2722431, -32'sd581502, 32'sd1201232, -32'sd49209, 32'sd1068865, -32'sd1458592, 32'sd2062608, 32'sd1369930, 32'sd2066010, 32'sd1346887, 32'sd670449, -32'sd2180303, -32'sd1695207, -32'sd1522761, -32'sd7694655, 32'sd803966, -32'sd1573188, -32'sd2656641, 32'sd1128705, -32'sd631814, -32'sd547117, 32'sd1370633, 32'sd1457587, 32'sd457450, -32'sd367736, -32'sd274750, 32'sd3225865, -32'sd830741, -32'sd151243, 32'sd693383, 32'sd863515, 32'sd1523357, -32'sd316349, 32'sd1274907, -32'sd913507, 32'sd516582, 32'sd578907, 32'sd1847272, -32'sd1118780, 32'sd295248, 32'sd923741, -32'sd601114, -32'sd8785679, 32'sd0, -32'sd8761415, -32'sd792131, 32'sd2321225, 32'sd2396292, 32'sd300037, 32'sd1647530, 32'sd279345, 32'sd2229221, 32'sd1436105, 32'sd1133502, 32'sd1611577, -32'sd105264, 32'sd3537280, 32'sd2494725, 32'sd365625, -32'sd1221029, 32'sd1360471, 32'sd728010, 32'sd1178514, 32'sd2764730, 32'sd1058560, -32'sd961668, 32'sd260414, -32'sd1643228, 32'sd430966, -32'sd67984, 32'sd0, 32'sd0, 32'sd0, -32'sd492123, 32'sd1051320, -32'sd697026, -32'sd1009301, 32'sd1018077, 32'sd95625, 32'sd161281, -32'sd1310053, 32'sd2323733, 32'sd2683350, 32'sd2258465, 32'sd3525555, 32'sd2437105, 32'sd1162378, 32'sd1824381, 32'sd442638, -32'sd221477, 32'sd817207, 32'sd927755, -32'sd439302, -32'sd1467557, -32'sd1013695, -32'sd157931, -32'sd1529960, -32'sd9397054, 32'sd0, 32'sd0, 32'sd0, -32'sd8463120, 32'sd557408, -32'sd20351, 32'sd64876, 32'sd2537821, 32'sd1614767, 32'sd1820850, 32'sd637035, 32'sd3204909, 32'sd2187251, 32'sd1284612, 32'sd1445720, 32'sd846819, 32'sd997989, 32'sd1153724, 32'sd1861056, -32'sd1647355, 32'sd1321707, 32'sd729086, -32'sd3069554, -32'sd148314, -32'sd3173752, -32'sd9359699, 32'sd748698, -32'sd8872872, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd7817343, 32'sd336568, -32'sd1846183, 32'sd922514, 32'sd2815612, 32'sd4810382, 32'sd1227151, 32'sd1485535, 32'sd1094675, 32'sd1530044, 32'sd156305, 32'sd556284, 32'sd1068334, 32'sd1518191, 32'sd502128, 32'sd1905981, 32'sd516526, -32'sd507599, -32'sd342576, 32'sd14349, -32'sd5588747, -32'sd7753507, -32'sd9169859, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd8035535, -32'sd9778525, -32'sd4333983, -32'sd3801518, 32'sd573619, 32'sd2547419, 32'sd1229381, -32'sd5114691, 32'sd3117849, -32'sd6084255, -32'sd5512086, -32'sd4098126, -32'sd1822840, -32'sd2370314, -32'sd4947631, -32'sd4580063, -32'sd9047515, -32'sd9695607, -32'sd9694201, -32'sd7384426, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd6204352, -32'sd6899449, -32'sd7127265, -32'sd6195762, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5630653, -32'sd6085613, -32'sd389463, 32'sd652262, -32'sd2983348, -32'sd7153819, -32'sd4921293, -32'sd713534, -32'sd711974, -32'sd779480, -32'sd4067530, -32'sd4990827, -32'sd1419632, -32'sd967388, -32'sd3084932, -32'sd7328597, -32'sd6565104, -32'sd6792905, -32'sd4954313, -32'sd5571329, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd6796838, -32'sd5601439, -32'sd6309222, 32'sd1247732, -32'sd385401, -32'sd671019, -32'sd1378782, -32'sd2418497, -32'sd2610402, -32'sd5394377, -32'sd5628765, -32'sd6955710, -32'sd7038458, -32'sd5236262, -32'sd6389895, -32'sd3248476, 32'sd790569, -32'sd6648932, -32'sd7774566, -32'sd4571651, -32'sd7341079, -32'sd7408718, -32'sd6699214, -32'sd6428809, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd7257062, -32'sd5879969, -32'sd7663621, -32'sd1399641, -32'sd1986566, -32'sd1991895, -32'sd3383314, -32'sd5110342, -32'sd6731456, -32'sd5063584, -32'sd4109496, -32'sd2322596, -32'sd5613197, -32'sd2714899, -32'sd4098181, -32'sd3519479, -32'sd2054560, -32'sd2762590, -32'sd2894534, 32'sd524737, -32'sd3722090, -32'sd3423630, -32'sd294418, -32'sd7509851, -32'sd5488370, 32'sd0, 32'sd0, -32'sd6519239, 32'sd1112200, -32'sd7275383, -32'sd534675, -32'sd1795329, -32'sd1416133, -32'sd374172, -32'sd2525925, -32'sd2764654, -32'sd2313145, -32'sd1258498, 32'sd174029, -32'sd1956810, -32'sd1378666, -32'sd1025046, -32'sd1830340, -32'sd871912, -32'sd526925, -32'sd2744390, -32'sd277589, 32'sd209384, -32'sd1901826, 32'sd619738, -32'sd1698119, 32'sd1011058, 32'sd786987, -32'sd958632, 32'sd0, -32'sd6379633, 32'sd742704, -32'sd2329572, 32'sd1288656, 32'sd1049931, 32'sd232624, -32'sd1382483, 32'sd1230608, -32'sd140793, -32'sd828718, 32'sd754109, 32'sd1611299, 32'sd1560581, -32'sd1532557, -32'sd1863055, -32'sd306185, -32'sd1269016, -32'sd1585447, -32'sd591880, -32'sd210635, -32'sd13006, -32'sd934899, 32'sd430792, 32'sd760456, -32'sd306290, 32'sd663446, 32'sd420651, 32'sd0, 32'sd24568, -32'sd758070, 32'sd895336, -32'sd722063, 32'sd618886, -32'sd1472595, 32'sd809771, -32'sd223583, 32'sd2729774, 32'sd1777184, 32'sd122226, 32'sd105500, 32'sd753381, 32'sd2508407, 32'sd2629190, 32'sd3302643, 32'sd2689925, -32'sd107021, -32'sd223279, -32'sd432297, 32'sd3875698, -32'sd1192872, 32'sd673762, -32'sd2670326, 32'sd711680, 32'sd2547287, -32'sd177246, -32'sd6081355, 32'sd991003, 32'sd839700, 32'sd2237773, 32'sd26236, -32'sd662079, 32'sd327055, 32'sd937325, 32'sd936146, 32'sd739028, -32'sd30087, 32'sd1006259, 32'sd1020436, 32'sd3116283, 32'sd1761576, 32'sd2419286, 32'sd902168, -32'sd1663358, -32'sd1522763, -32'sd3706697, -32'sd74278, -32'sd32757, 32'sd975087, 32'sd26742, -32'sd934638, -32'sd2305225, 32'sd152239, -32'sd2097500, 32'sd71236, 32'sd2575244, 32'sd732266, -32'sd104348, 32'sd409772, 32'sd674672, 32'sd1262109, 32'sd974776, 32'sd1901847, 32'sd567904, 32'sd2053209, 32'sd1155475, 32'sd1627549, 32'sd4801438, 32'sd3197222, 32'sd1557543, 32'sd88089, -32'sd3959382, 32'sd260865, -32'sd121678, -32'sd2942835, -32'sd2370400, -32'sd92048, -32'sd1391168, -32'sd2602751, -32'sd375078, -32'sd337855, -32'sd3748295, 32'sd1341729, 32'sd251458, 32'sd1178833, 32'sd1250182, 32'sd1168444, 32'sd1278047, 32'sd225859, 32'sd978216, 32'sd772130, 32'sd2398820, 32'sd3874904, 32'sd3850215, 32'sd1349663, 32'sd2763384, 32'sd2280833, 32'sd370465, -32'sd587699, 32'sd381621, -32'sd2344588, -32'sd1961430, -32'sd600340, -32'sd2482978, -32'sd1411109, 32'sd471117, -32'sd351312, -32'sd968593, 32'sd1379877, 32'sd350899, -32'sd279317, -32'sd254469, 32'sd827993, -32'sd531229, 32'sd265387, 32'sd66885, 32'sd1989445, 32'sd721730, 32'sd2037356, 32'sd2722218, 32'sd3045274, 32'sd2715922, 32'sd677833, 32'sd607598, -32'sd726195, -32'sd2584111, 32'sd2795182, -32'sd690989, 32'sd1166192, -32'sd1154892, 32'sd361303, -32'sd691325, 32'sd1146829, 32'sd366622, 32'sd400510, -32'sd284859, -32'sd274909, 32'sd108609, 32'sd1859351, -32'sd311960, -32'sd1746407, 32'sd2133418, 32'sd148314, -32'sd1737938, 32'sd1997300, 32'sd4284699, 32'sd4157682, 32'sd3006405, 32'sd2640504, 32'sd3916139, -32'sd2299490, -32'sd1278569, 32'sd815976, 32'sd1378492, 32'sd2724244, 32'sd2138928, -32'sd86495, -32'sd538871, 32'sd1016296, -32'sd424535, 32'sd3022837, -32'sd3196835, 32'sd452339, 32'sd387574, -32'sd402331, -32'sd500496, 32'sd1090599, -32'sd542391, 32'sd319529, 32'sd1158680, 32'sd2600838, 32'sd2346474, 32'sd600991, 32'sd1490299, -32'sd473951, -32'sd2448577, -32'sd6294480, -32'sd5895764, -32'sd3172868, -32'sd3285199, -32'sd1918150, 32'sd2299280, 32'sd2078625, 32'sd4221158, 32'sd1798055, 32'sd793769, 32'sd686961, 32'sd2017108, 32'sd3474326, -32'sd1064698, -32'sd274502, -32'sd205653, -32'sd455711, 32'sd477220, -32'sd225374, 32'sd254896, -32'sd72958, 32'sd871362, 32'sd629737, -32'sd247120, 32'sd688594, -32'sd1327645, -32'sd2578130, -32'sd3317593, -32'sd4293302, -32'sd3364642, -32'sd3463103, -32'sd1583344, 32'sd1175921, 32'sd1271771, 32'sd2623249, 32'sd2083584, 32'sd2885541, 32'sd589301, 32'sd1458405, 32'sd2974499, 32'sd2745712, 32'sd1615925, -32'sd771042, -32'sd833696, -32'sd3143270, -32'sd1213928, -32'sd4666871, 32'sd603628, 32'sd485154, 32'sd1179519, -32'sd2325514, -32'sd1970017, -32'sd2393923, -32'sd4714140, -32'sd3535796, -32'sd4834055, -32'sd3865107, -32'sd1057518, 32'sd108352, 32'sd770521, -32'sd279699, 32'sd1030132, 32'sd1810786, 32'sd2635872, 32'sd3856645, 32'sd327794, -32'sd143028, 32'sd1261108, 32'sd1394525, 32'sd982813, -32'sd2980105, 32'sd88924, 32'sd526503, -32'sd5551549, -32'sd6294801, -32'sd3332744, -32'sd1507735, 32'sd768096, -32'sd2202913, -32'sd3802269, -32'sd3654526, -32'sd1907689, -32'sd2881432, -32'sd494296, -32'sd695302, -32'sd938811, -32'sd53183, 32'sd1088161, 32'sd1821524, 32'sd2819949, 32'sd516547, 32'sd2599405, 32'sd1231881, 32'sd844919, 32'sd1547599, 32'sd405898, 32'sd1173396, 32'sd748750, 32'sd400302, -32'sd193112, -32'sd1899912, -32'sd7145571, -32'sd6846863, -32'sd2040607, -32'sd1276314, 32'sd892344, -32'sd406578, -32'sd1339648, -32'sd1090817, 32'sd505113, -32'sd875510, -32'sd2723863, -32'sd1603795, 32'sd221044, 32'sd1126372, 32'sd1297659, 32'sd2345230, 32'sd1022398, 32'sd1584383, -32'sd639521, -32'sd1922379, -32'sd2347917, 32'sd225689, 32'sd445812, -32'sd709041, 32'sd1563721, 32'sd492534, -32'sd192649, -32'sd919817, -32'sd3495261, 32'sd0, 32'sd953245, 32'sd1735551, -32'sd170821, -32'sd2635241, -32'sd3589245, -32'sd2555499, -32'sd3009329, -32'sd2605503, -32'sd200093, 32'sd405169, 32'sd2717214, 32'sd3579029, 32'sd2906946, 32'sd1412497, 32'sd980650, 32'sd1043840, -32'sd566260, -32'sd509586, -32'sd268678, 32'sd402499, -32'sd2452171, -32'sd739946, -32'sd387233, 32'sd550001, 32'sd2404390, 32'sd4253455, 32'sd474654, -32'sd6302248, -32'sd492457, 32'sd2616632, -32'sd3483652, -32'sd4665892, -32'sd338048, -32'sd3015043, -32'sd3386902, -32'sd4354441, -32'sd845228, 32'sd1696647, 32'sd2385645, 32'sd787941, 32'sd2746557, 32'sd135526, 32'sd1254250, -32'sd1785349, -32'sd22833, -32'sd1032767, -32'sd1331864, -32'sd27302, -32'sd4209454, -32'sd2089480, -32'sd2045380, -32'sd2637265, -32'sd1879815, 32'sd2383485, 32'sd483380, -32'sd7016417, 32'sd2266840, 32'sd896345, -32'sd1815631, 32'sd930137, -32'sd2032334, -32'sd1431686, -32'sd2150821, -32'sd3201250, -32'sd683765, 32'sd4475351, 32'sd652100, 32'sd2436039, -32'sd270062, -32'sd452350, 32'sd187231, -32'sd1021902, 32'sd479575, -32'sd1516086, -32'sd919762, -32'sd2502491, -32'sd1106852, -32'sd380350, 32'sd826156, -32'sd567675, -32'sd2806365, -32'sd1659103, -32'sd1995941, 32'sd0, -32'sd674708, -32'sd350066, -32'sd427142, -32'sd1553352, -32'sd2360270, 32'sd1098180, -32'sd486417, 32'sd1569581, 32'sd1100351, 32'sd1558960, 32'sd476290, 32'sd688801, 32'sd1258059, -32'sd167051, -32'sd74818, 32'sd190708, -32'sd2216264, -32'sd2223682, -32'sd537334, -32'sd910220, -32'sd537041, -32'sd84556, -32'sd286616, 32'sd2292003, 32'sd996780, -32'sd739556, -32'sd6163190, -32'sd7155729, -32'sd5072490, -32'sd2831921, -32'sd40529, -32'sd2700854, 32'sd91692, -32'sd2155678, -32'sd751833, 32'sd424322, -32'sd2205441, 32'sd783685, -32'sd272193, -32'sd133030, 32'sd1031706, 32'sd1314339, 32'sd1133938, 32'sd667875, 32'sd118774, -32'sd868300, -32'sd20720, -32'sd2621379, -32'sd1137084, -32'sd1655194, -32'sd1877733, -32'sd1099098, 32'sd1665, -32'sd211678, 32'sd674605, -32'sd5816066, -32'sd6369745, -32'sd2619500, -32'sd947003, 32'sd1320413, 32'sd1514227, 32'sd852054, -32'sd1816800, -32'sd627258, -32'sd1451679, -32'sd5360, -32'sd630912, 32'sd1103817, -32'sd144758, 32'sd1801461, 32'sd1141294, 32'sd567602, -32'sd1325127, -32'sd920970, -32'sd200675, -32'sd312135, 32'sd530502, -32'sd1618503, 32'sd1261370, -32'sd2044950, -32'sd608392, 32'sd1419780, 32'sd767051, 32'sd0, -32'sd6508377, 32'sd3334, -32'sd4266356, -32'sd2761879, 32'sd467445, -32'sd653877, -32'sd1676507, 32'sd1342814, 32'sd1063598, -32'sd1712159, -32'sd337095, -32'sd412460, -32'sd1450965, 32'sd2985, 32'sd2404612, -32'sd998172, 32'sd81411, -32'sd1143624, -32'sd1087856, -32'sd1140498, -32'sd1367005, 32'sd1916142, 32'sd798620, 32'sd1140728, -32'sd712590, -32'sd7395372, 32'sd0, 32'sd0, 32'sd0, 32'sd1166085, 32'sd1506872, -32'sd805643, 32'sd151616, 32'sd412276, -32'sd921124, -32'sd638350, -32'sd2183987, -32'sd2201412, -32'sd2505088, -32'sd1048973, -32'sd1591577, -32'sd1456371, -32'sd6812, -32'sd1157509, -32'sd715316, 32'sd319103, 32'sd339851, 32'sd3016070, -32'sd395618, 32'sd1638152, 32'sd160423, 32'sd928135, -32'sd511436, 32'sd1185651, 32'sd0, 32'sd0, 32'sd0, -32'sd2973019, -32'sd562797, 32'sd256361, 32'sd591257, 32'sd1283445, -32'sd1304610, 32'sd627824, -32'sd988667, -32'sd631798, 32'sd64937, -32'sd126639, 32'sd633078, 32'sd1695071, 32'sd678047, 32'sd163227, 32'sd1238303, -32'sd1878518, 32'sd1018575, 32'sd548663, -32'sd521136, -32'sd1217534, -32'sd383107, -32'sd317250, 32'sd396074, 32'sd60273, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5880773, -32'sd3013567, -32'sd1869196, -32'sd477759, 32'sd2392061, 32'sd1371314, 32'sd2820228, 32'sd1774740, 32'sd300676, 32'sd767398, 32'sd1193040, 32'sd1486922, 32'sd2446, 32'sd121704, 32'sd1268084, 32'sd1809522, 32'sd1395070, 32'sd742777, -32'sd239527, 32'sd1592502, -32'sd875844, -32'sd2088098, 32'sd1187308, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5771027, -32'sd5071387, 32'sd1246387, 32'sd1485409, -32'sd10373, 32'sd917429, 32'sd676275, 32'sd470269, -32'sd331901, -32'sd706737, 32'sd2752368, 32'sd3407270, 32'sd797119, 32'sd554994, 32'sd586658, 32'sd996291, 32'sd1087614, 32'sd1127438, 32'sd90438, -32'sd6321765, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4150389, -32'sd4650327, -32'sd3841197, -32'sd2854939, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5296159, -32'sd3601608, -32'sd3830457, -32'sd3724143, -32'sd1761586, -32'sd653635, -32'sd919485, -32'sd2364964, -32'sd4631848, -32'sd3134388, 32'sd1466349, 32'sd1202375, 32'sd991911, -32'sd1198876, -32'sd2872542, -32'sd3019432, 32'sd272128, -32'sd939056, -32'sd4721779, -32'sd3568785, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5164485, -32'sd972445, 32'sd301228, -32'sd620602, -32'sd3618381, -32'sd1167872, -32'sd2186554, -32'sd339011, 32'sd1113786, 32'sd792480, 32'sd1684216, -32'sd1848980, 32'sd224452, 32'sd169490, 32'sd1726781, -32'sd771628, -32'sd1046037, -32'sd5708479, -32'sd2258862, -32'sd1648185, -32'sd998266, -32'sd2695287, -32'sd3576719, -32'sd3760065, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2617839, 32'sd1222289, -32'sd423605, -32'sd3368393, 32'sd596716, 32'sd1791589, 32'sd2812868, 32'sd2823839, -32'sd524114, 32'sd1165116, 32'sd1245947, 32'sd1487972, 32'sd1202572, -32'sd431441, 32'sd1621283, 32'sd940508, 32'sd1084400, 32'sd366179, 32'sd812467, 32'sd848771, 32'sd29153, 32'sd645453, -32'sd2189461, -32'sd5677015, -32'sd5287854, 32'sd0, 32'sd0, -32'sd3679687, -32'sd1419337, -32'sd598976, 32'sd610570, 32'sd1855084, 32'sd957012, -32'sd324439, 32'sd769659, 32'sd805413, 32'sd2667237, 32'sd1264534, 32'sd3581083, 32'sd163505, 32'sd1833753, 32'sd132107, 32'sd359706, 32'sd267507, 32'sd1884831, 32'sd1723840, -32'sd277098, -32'sd1913811, 32'sd560038, -32'sd1430666, 32'sd204309, -32'sd2190924, -32'sd4101504, -32'sd3371910, 32'sd0, -32'sd5347773, 32'sd721028, 32'sd1381337, -32'sd842026, -32'sd136567, 32'sd821709, 32'sd453988, -32'sd671889, -32'sd1406820, 32'sd378611, -32'sd243480, 32'sd1650299, 32'sd900598, 32'sd1581625, 32'sd2857864, 32'sd2553680, 32'sd866772, 32'sd780531, -32'sd850244, 32'sd967338, -32'sd1005350, 32'sd1004645, 32'sd518341, -32'sd621140, 32'sd373906, 32'sd615140, -32'sd4970004, 32'sd0, -32'sd4685102, -32'sd2149259, 32'sd1193122, 32'sd457733, -32'sd163015, 32'sd698896, -32'sd1610064, -32'sd1116549, 32'sd294464, 32'sd1811030, 32'sd30829, 32'sd1174414, 32'sd1503042, 32'sd2063440, 32'sd1625919, 32'sd147250, -32'sd643080, 32'sd532365, 32'sd20915, 32'sd1968516, -32'sd1857575, -32'sd175818, 32'sd1204005, -32'sd2509051, -32'sd554871, 32'sd853595, -32'sd5626566, -32'sd4378867, -32'sd5743421, -32'sd1495987, 32'sd1013180, 32'sd444533, -32'sd1082640, 32'sd1087235, 32'sd746043, 32'sd1036650, 32'sd633545, 32'sd1197757, 32'sd925721, 32'sd1108814, 32'sd1745920, 32'sd3671190, 32'sd2604401, 32'sd780452, 32'sd2358901, -32'sd569281, 32'sd832688, -32'sd2270126, -32'sd455218, -32'sd507249, -32'sd1185001, 32'sd1127716, -32'sd726651, -32'sd511594, -32'sd4810483, -32'sd4177757, -32'sd2417259, 32'sd119875, 32'sd1225998, 32'sd3395880, -32'sd576076, -32'sd132923, 32'sd238373, -32'sd16408, 32'sd1108360, 32'sd2082319, 32'sd1417976, 32'sd1537246, 32'sd1247098, 32'sd1233870, 32'sd2044176, -32'sd880475, 32'sd1484493, -32'sd1662128, 32'sd4147421, 32'sd285103, -32'sd2834335, 32'sd1588638, -32'sd2119219, -32'sd2641895, -32'sd1199268, 32'sd650531, -32'sd3976672, 32'sd778138, -32'sd1182955, 32'sd225867, 32'sd577961, 32'sd924661, 32'sd779121, -32'sd1015771, 32'sd1254631, -32'sd768248, 32'sd1513921, -32'sd508918, -32'sd2054002, -32'sd1193494, -32'sd2711721, -32'sd584913, 32'sd3140567, 32'sd1177433, 32'sd1256639, -32'sd75449, 32'sd358955, -32'sd1853377, -32'sd1051637, 32'sd751359, 32'sd2703198, -32'sd4020165, -32'sd1952881, -32'sd2976731, -32'sd4298659, -32'sd612704, 32'sd98271, -32'sd573404, 32'sd1685972, -32'sd1875116, 32'sd1108667, 32'sd3618381, -32'sd413784, -32'sd231502, -32'sd4029538, -32'sd4919455, -32'sd4427183, -32'sd4760771, -32'sd5888951, -32'sd830266, -32'sd2225982, 32'sd72085, 32'sd1199364, 32'sd737458, 32'sd3017570, -32'sd1820207, -32'sd484413, -32'sd488560, 32'sd1678622, -32'sd7263770, -32'sd484147, 32'sd114354, 32'sd1689043, -32'sd417646, 32'sd412880, 32'sd1089485, 32'sd209023, 32'sd429392, 32'sd2010491, 32'sd1406261, -32'sd2328461, -32'sd5589283, -32'sd6064364, -32'sd5155823, -32'sd4890149, -32'sd4737377, -32'sd2890300, 32'sd429046, -32'sd744011, -32'sd1226741, -32'sd2469, -32'sd637535, 32'sd1450252, 32'sd2126663, -32'sd1823941, 32'sd1358567, 32'sd202220, -32'sd2910125, -32'sd1415437, 32'sd995614, 32'sd1041244, -32'sd5272080, -32'sd1685487, -32'sd1708022, 32'sd113910, 32'sd1079959, 32'sd852963, -32'sd4238134, -32'sd7370164, -32'sd5052277, -32'sd3531765, -32'sd856224, -32'sd1765568, -32'sd1579318, -32'sd1035971, 32'sd2523611, 32'sd300268, -32'sd97519, -32'sd70138, -32'sd1566018, 32'sd1440143, -32'sd3263313, -32'sd1398441, -32'sd1626398, -32'sd74289, 32'sd1238892, -32'sd1032311, 32'sd291060, -32'sd4185408, -32'sd4167427, -32'sd3663767, -32'sd1806410, -32'sd786585, -32'sd2067896, -32'sd4192656, -32'sd9388633, -32'sd6730438, -32'sd892786, 32'sd796744, -32'sd4325833, -32'sd3401158, -32'sd2732822, 32'sd3599819, 32'sd4254593, 32'sd4113, -32'sd1330714, -32'sd1623384, 32'sd77490, -32'sd2519385, -32'sd290723, -32'sd2589876, -32'sd1446702, -32'sd2452333, -32'sd2114048, 32'sd219372, 32'sd1153753, -32'sd4619392, -32'sd4279455, -32'sd5585182, -32'sd1932739, -32'sd405610, -32'sd4841067, -32'sd9516696, -32'sd6994997, -32'sd4849580, -32'sd2904300, -32'sd2018371, -32'sd758400, -32'sd556041, -32'sd1746934, 32'sd2658243, 32'sd5064886, 32'sd1417239, 32'sd294698, -32'sd2616458, -32'sd1471485, -32'sd1217288, -32'sd1024900, -32'sd1280022, -32'sd5248391, -32'sd3237187, -32'sd2612259, -32'sd205194, 32'sd337696, -32'sd4732536, -32'sd3865925, -32'sd4206013, 32'sd1043066, 32'sd1716436, -32'sd8364690, -32'sd3619489, -32'sd2349127, -32'sd1887180, -32'sd507736, -32'sd1619419, -32'sd1746345, -32'sd83928, 32'sd127082, 32'sd4536620, 32'sd4724826, 32'sd787801, -32'sd2300193, -32'sd1512777, -32'sd3175783, -32'sd4440964, -32'sd1770905, -32'sd407001, -32'sd1091316, 32'sd1187475, -32'sd1010819, 32'sd317311, -32'sd1980307, -32'sd5478146, -32'sd3939974, -32'sd4611419, 32'sd193330, 32'sd775600, -32'sd2225734, 32'sd1025858, 32'sd1638010, 32'sd1765955, 32'sd1020216, 32'sd2240005, 32'sd438270, 32'sd2905914, 32'sd3513336, 32'sd2682872, 32'sd2742888, 32'sd32788, -32'sd1453851, -32'sd2923706, -32'sd2016026, -32'sd2239896, -32'sd2840215, -32'sd975427, 32'sd1889448, -32'sd368826, 32'sd816982, 32'sd515271, -32'sd766302, 32'sd353400, 32'sd0, -32'sd4888096, -32'sd2427445, -32'sd268952, 32'sd997447, -32'sd994655, 32'sd148627, 32'sd1680687, 32'sd3019555, 32'sd2247215, 32'sd314111, 32'sd932887, 32'sd2892689, -32'sd1348625, 32'sd35723, -32'sd526593, -32'sd1318511, -32'sd2845891, -32'sd1734446, -32'sd1210304, -32'sd978305, 32'sd90333, 32'sd2619167, 32'sd1907851, 32'sd226119, 32'sd1122703, -32'sd579731, 32'sd1223992, -32'sd3178011, -32'sd5126990, -32'sd257193, 32'sd1061752, -32'sd1281846, 32'sd1699908, 32'sd2322219, -32'sd724267, -32'sd876084, 32'sd1304630, 32'sd642586, 32'sd761753, -32'sd382248, -32'sd1880357, -32'sd2950213, 32'sd113771, -32'sd59815, -32'sd868597, 32'sd1148694, 32'sd311025, 32'sd2700426, -32'sd1860577, 32'sd1708194, 32'sd772717, 32'sd931424, 32'sd2410468, -32'sd23423, 32'sd3511548, -32'sd5071194, -32'sd3398400, -32'sd861401, -32'sd791678, 32'sd1503457, 32'sd885303, -32'sd285720, 32'sd818601, -32'sd1971760, 32'sd845502, 32'sd1148066, -32'sd1993943, -32'sd1905049, 32'sd1164069, -32'sd2162499, 32'sd719872, 32'sd1630584, 32'sd1166572, 32'sd822077, 32'sd1746900, 32'sd560123, -32'sd151882, 32'sd952705, 32'sd1399343, -32'sd1645105, 32'sd3280814, 32'sd2322570, -32'sd253299, 32'sd0, -32'sd802024, 32'sd1424113, 32'sd1895612, 32'sd3187041, -32'sd24574, 32'sd2834687, 32'sd2511354, 32'sd1083549, 32'sd2007180, -32'sd1045644, -32'sd708411, 32'sd693468, -32'sd1911757, -32'sd898679, 32'sd145020, 32'sd677190, 32'sd2322967, 32'sd2643945, 32'sd2730306, 32'sd3184735, 32'sd1804895, -32'sd368702, 32'sd2923526, 32'sd616421, -32'sd1306629, 32'sd1329865, -32'sd3175932, 32'sd334499, -32'sd1103180, 32'sd3119122, 32'sd3226495, 32'sd53567, -32'sd241661, 32'sd1739761, 32'sd2471251, 32'sd1957901, 32'sd96902, -32'sd28811, 32'sd157088, 32'sd2247348, 32'sd553615, 32'sd447013, 32'sd862011, 32'sd639002, 32'sd1952127, 32'sd4593935, 32'sd3145542, 32'sd1401161, 32'sd659770, -32'sd125860, -32'sd1138467, -32'sd36180, 32'sd998420, 32'sd717307, -32'sd5041792, 32'sd888757, 32'sd118764, 32'sd1507659, 32'sd1381074, 32'sd29669, 32'sd4921520, 32'sd1065713, 32'sd1097079, 32'sd1110508, 32'sd1482516, 32'sd943104, -32'sd248836, -32'sd333279, -32'sd401475, -32'sd1114915, -32'sd900556, 32'sd750920, 32'sd1324786, 32'sd1178222, 32'sd1817529, 32'sd2251136, 32'sd2357878, -32'sd874396, -32'sd1106468, 32'sd2349464, -32'sd168140, -32'sd604824, -32'sd3414891, 32'sd0, -32'sd4178227, 32'sd788631, -32'sd803080, -32'sd269423, 32'sd3250960, 32'sd329675, 32'sd1268180, 32'sd279395, 32'sd3165517, 32'sd902275, 32'sd455810, 32'sd515764, 32'sd1023443, -32'sd864129, -32'sd679870, 32'sd754653, -32'sd314859, 32'sd1501935, 32'sd1463729, 32'sd3916782, 32'sd2955653, 32'sd9832, 32'sd1081809, 32'sd362105, 32'sd493686, -32'sd2307718, 32'sd0, 32'sd0, 32'sd0, -32'sd267589, -32'sd236829, 32'sd602, -32'sd381510, 32'sd1381628, -32'sd605623, 32'sd1234223, 32'sd630114, -32'sd2048595, 32'sd2288923, 32'sd2259101, 32'sd2431207, 32'sd1239552, -32'sd1021146, -32'sd418907, 32'sd557029, 32'sd895557, 32'sd1285897, -32'sd2327832, 32'sd180808, 32'sd994096, -32'sd552176, -32'sd1469010, 32'sd1618239, -32'sd5399143, 32'sd0, 32'sd0, 32'sd0, -32'sd4901147, 32'sd248275, 32'sd1432538, -32'sd329473, 32'sd841688, -32'sd1690656, 32'sd1209243, -32'sd103415, 32'sd2691309, 32'sd582085, -32'sd555171, -32'sd443692, 32'sd1239251, -32'sd491111, 32'sd151588, 32'sd1093439, -32'sd3227689, -32'sd1283506, -32'sd213124, -32'sd512719, -32'sd776488, -32'sd393611, -32'sd4906268, 32'sd394894, -32'sd3619206, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd4029982, -32'sd2593197, -32'sd1056606, 32'sd63544, 32'sd820688, -32'sd64674, 32'sd900890, 32'sd170767, 32'sd400986, -32'sd1706812, 32'sd2006731, 32'sd43341, 32'sd382176, -32'sd2432159, -32'sd1178613, -32'sd307893, -32'sd280791, 32'sd1082693, -32'sd891667, -32'sd70658, -32'sd5344284, -32'sd4744137, -32'sd4867496, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd5295413, -32'sd3580892, -32'sd2624697, -32'sd1095476, 32'sd586666, -32'sd295519, 32'sd2571134, -32'sd1087988, -32'sd1073075, -32'sd3303588, -32'sd4436843, -32'sd4697068, -32'sd4244356, -32'sd412367, -32'sd145857, -32'sd382550, -32'sd461904, -32'sd3621082, -32'sd4750718, -32'sd3581971, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd639565, -32'sd1033035, -32'sd173983, 32'sd320675, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd15139, -32'sd1002430, 32'sd464578, 32'sd325157, -32'sd778036, 32'sd374607, -32'sd114958, -32'sd135128, 32'sd1113511, -32'sd595172, 32'sd1624233, 32'sd1229047, -32'sd1858254, 32'sd296261, 32'sd380591, 32'sd702426, 32'sd334172, -32'sd82929, -32'sd150538, -32'sd55387, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2256454, 32'sd653756, 32'sd1164740, 32'sd424165, -32'sd2066142, -32'sd554527, -32'sd58792, -32'sd3061038, -32'sd4019818, -32'sd1154230, 32'sd944675, 32'sd4388199, 32'sd847516, 32'sd2255679, 32'sd4550087, 32'sd1284900, -32'sd21503, 32'sd3228695, 32'sd1680866, 32'sd2126738, 32'sd578409, -32'sd2226284, 32'sd2510718, -32'sd707437, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd1665702, 32'sd2035837, -32'sd568659, -32'sd1880343, 32'sd22221, -32'sd1329256, -32'sd2029354, -32'sd416186, 32'sd897371, -32'sd2581779, 32'sd1671396, 32'sd1672232, -32'sd1018690, -32'sd1252179, -32'sd434135, 32'sd1447197, -32'sd499699, 32'sd798779, 32'sd1165246, 32'sd269812, 32'sd440448, 32'sd1576587, 32'sd1487116, -32'sd706373, 32'sd802621, 32'sd0, 32'sd0, 32'sd550365, 32'sd1023251, 32'sd920657, -32'sd238431, -32'sd2440540, -32'sd318239, -32'sd2338037, 32'sd784583, -32'sd1863980, -32'sd948083, -32'sd595568, -32'sd247980, -32'sd698964, -32'sd490779, -32'sd2276793, -32'sd911765, -32'sd1472071, -32'sd1439410, 32'sd2746461, -32'sd564185, -32'sd939933, 32'sd158534, 32'sd987572, 32'sd67688, -32'sd295818, 32'sd322563, -32'sd1377170, 32'sd0, -32'sd325595, 32'sd1573282, 32'sd136005, 32'sd283820, 32'sd3156207, 32'sd3279654, -32'sd379103, -32'sd2103647, -32'sd4200548, -32'sd2421143, -32'sd1996044, -32'sd1517718, 32'sd807059, 32'sd45063, 32'sd2041912, -32'sd4005440, -32'sd2440863, -32'sd3066250, -32'sd1115832, -32'sd4269799, -32'sd2456290, -32'sd569899, 32'sd296911, -32'sd329367, -32'sd875448, 32'sd95643, -32'sd794922, 32'sd0, 32'sd337907, -32'sd1286293, -32'sd455499, -32'sd229244, -32'sd1944383, 32'sd310545, -32'sd501908, -32'sd1161577, -32'sd4333580, -32'sd1143083, 32'sd482945, 32'sd2022367, 32'sd47427, -32'sd1530852, -32'sd538785, -32'sd1914634, -32'sd219531, -32'sd822823, -32'sd541047, 32'sd3312, 32'sd765504, 32'sd276197, -32'sd2296947, -32'sd914135, -32'sd1083662, 32'sd866874, -32'sd724641, 32'sd1566472, 32'sd1034720, -32'sd383618, 32'sd626138, 32'sd687448, -32'sd1616013, 32'sd303721, 32'sd271840, -32'sd2144815, -32'sd719688, 32'sd138616, 32'sd296433, 32'sd2541956, 32'sd915352, -32'sd562827, -32'sd2970297, 32'sd1253951, 32'sd607656, -32'sd1877642, 32'sd109439, 32'sd1354978, -32'sd1342491, 32'sd552515, 32'sd2827139, 32'sd1143433, -32'sd1402987, 32'sd673741, -32'sd32958, 32'sd1123967, -32'sd2010973, -32'sd180082, -32'sd561678, -32'sd2259014, -32'sd96460, -32'sd289929, 32'sd1928050, 32'sd612575, 32'sd2940479, 32'sd1047420, 32'sd1604132, 32'sd334600, 32'sd1473046, 32'sd4066818, 32'sd2323419, -32'sd3612063, -32'sd632229, -32'sd3009866, -32'sd610044, 32'sd93418, 32'sd1246789, 32'sd3357031, 32'sd1315938, 32'sd3527875, 32'sd486710, 32'sd303017, 32'sd254685, 32'sd682881, 32'sd243295, 32'sd375943, 32'sd1575383, -32'sd4117948, -32'sd2628700, 32'sd2666404, 32'sd2116744, -32'sd926311, -32'sd2240509, 32'sd1089198, -32'sd104636, -32'sd579877, 32'sd4677426, 32'sd2676788, 32'sd2557676, -32'sd990259, 32'sd309270, -32'sd1960009, 32'sd1487971, -32'sd120765, -32'sd1532366, -32'sd1445312, 32'sd2476498, 32'sd514473, 32'sd1808241, -32'sd968987, 32'sd1106626, 32'sd305152, -32'sd1447145, 32'sd1427589, -32'sd1743393, 32'sd758807, -32'sd3089304, -32'sd741944, -32'sd2142858, 32'sd793680, -32'sd695328, 32'sd981618, 32'sd699562, -32'sd877503, 32'sd2701177, 32'sd1842480, 32'sd2411629, 32'sd634356, 32'sd497598, -32'sd1798647, -32'sd993272, -32'sd420650, -32'sd1606336, 32'sd611955, -32'sd261631, -32'sd886684, 32'sd307673, 32'sd201886, 32'sd1526294, 32'sd349519, -32'sd968175, -32'sd1150469, 32'sd1301287, 32'sd1763577, -32'sd2249549, -32'sd3129119, -32'sd1813583, 32'sd1310411, 32'sd307809, 32'sd889370, 32'sd242878, 32'sd594408, 32'sd2125779, 32'sd4101524, 32'sd4512232, 32'sd2333922, 32'sd1275521, 32'sd1311755, 32'sd781410, 32'sd1159947, 32'sd1118415, 32'sd1971978, -32'sd46402, -32'sd1743876, -32'sd4112693, 32'sd827483, 32'sd217661, -32'sd214910, -32'sd1032185, 32'sd512839, -32'sd585002, -32'sd2011835, -32'sd1182286, -32'sd2090615, -32'sd1025176, 32'sd483573, 32'sd63383, -32'sd307068, 32'sd1746816, 32'sd2777912, 32'sd4590140, 32'sd4721342, 32'sd3217847, 32'sd1711753, 32'sd223226, -32'sd825008, 32'sd1696333, 32'sd2624095, 32'sd410780, -32'sd1162217, -32'sd1852977, -32'sd2215398, -32'sd3586932, -32'sd2075815, -32'sd1278677, 32'sd633774, 32'sd537429, 32'sd1783063, -32'sd616198, 32'sd518886, 32'sd19509, 32'sd409402, -32'sd184184, -32'sd699185, -32'sd249355, 32'sd384098, 32'sd407965, 32'sd832919, 32'sd2249107, 32'sd4896390, 32'sd4376845, 32'sd2759414, 32'sd269447, -32'sd967003, -32'sd5516, 32'sd2910059, 32'sd2594991, 32'sd143830, -32'sd2528776, -32'sd1169848, -32'sd445359, -32'sd1853177, -32'sd465983, 32'sd1111682, -32'sd605859, 32'sd2224347, 32'sd573098, 32'sd1632030, 32'sd643715, -32'sd1147713, -32'sd664559, -32'sd794939, -32'sd1252647, -32'sd1586758, -32'sd1106331, 32'sd931345, 32'sd2404324, 32'sd5450521, 32'sd4792377, 32'sd1796146, 32'sd945576, 32'sd580392, -32'sd861600, -32'sd714310, -32'sd1792447, -32'sd2253481, -32'sd2649296, -32'sd3455288, -32'sd906760, 32'sd832318, 32'sd91473, -32'sd1422475, -32'sd481747, -32'sd812432, 32'sd1614911, -32'sd332762, -32'sd3868581, -32'sd3744870, -32'sd3571114, -32'sd1619375, -32'sd200376, -32'sd1399985, 32'sd2584744, 32'sd267851, 32'sd3546735, 32'sd5885194, 32'sd1034273, 32'sd821318, -32'sd712922, -32'sd45461, -32'sd2822541, -32'sd1301041, 32'sd441247, -32'sd2394116, 32'sd347119, -32'sd3437322, -32'sd544118, 32'sd579339, -32'sd456603, 32'sd101388, 32'sd1197553, 32'sd741903, -32'sd1797141, -32'sd112888, -32'sd940920, 32'sd21202, 32'sd1170303, 32'sd964026, -32'sd2080583, 32'sd283987, 32'sd3401883, 32'sd1496864, 32'sd3484175, 32'sd3922371, 32'sd1631009, 32'sd2264624, -32'sd266592, -32'sd3267919, -32'sd4429206, -32'sd1696663, -32'sd490286, -32'sd5313803, -32'sd408102, -32'sd1801715, -32'sd5464439, 32'sd22898, -32'sd718486, 32'sd0, 32'sd1478384, 32'sd79145, -32'sd552836, 32'sd1834819, -32'sd4093927, -32'sd525091, -32'sd1564392, 32'sd1146088, -32'sd909140, 32'sd1593112, -32'sd1182215, -32'sd1389279, 32'sd2130474, 32'sd4559432, 32'sd1461775, 32'sd30572, -32'sd2414019, -32'sd5021476, -32'sd3516158, -32'sd3109574, -32'sd1488979, -32'sd1891832, -32'sd1273106, -32'sd2136795, -32'sd3818510, 32'sd650311, 32'sd95811, 32'sd1037769, -32'sd896528, -32'sd5170, -32'sd167781, -32'sd2905403, -32'sd5532634, -32'sd2364306, 32'sd211614, -32'sd1452125, -32'sd2983425, -32'sd5511369, -32'sd2858360, -32'sd2833281, 32'sd772872, 32'sd1505259, -32'sd203274, -32'sd2653591, -32'sd4220436, -32'sd3386384, -32'sd2261964, -32'sd2043633, -32'sd1484226, -32'sd6082154, -32'sd3631561, -32'sd5509747, -32'sd513119, 32'sd2577784, 32'sd113571, 32'sd559135, -32'sd900116, -32'sd812611, -32'sd1723041, -32'sd526330, -32'sd5038486, -32'sd2081099, -32'sd1300549, -32'sd3872158, -32'sd768139, -32'sd3925322, -32'sd4473171, -32'sd3412285, -32'sd345372, 32'sd812174, -32'sd2392008, -32'sd4210743, -32'sd3346153, -32'sd2624323, 32'sd685095, 32'sd132205, 32'sd1430330, -32'sd4549291, -32'sd3237609, -32'sd3100723, 32'sd1667594, 32'sd1043804, 32'sd140265, 32'sd0, 32'sd1469245, -32'sd3197313, -32'sd5649255, -32'sd3749965, -32'sd3819205, 32'sd148851, -32'sd1284282, -32'sd2487211, -32'sd949685, -32'sd2424492, -32'sd1705157, -32'sd422211, -32'sd2223306, 32'sd2458860, -32'sd1606731, 32'sd192132, 32'sd475300, -32'sd2183317, 32'sd477401, -32'sd2650865, -32'sd2241496, -32'sd4369894, -32'sd902023, -32'sd251075, 32'sd2232982, 32'sd1264605, 32'sd172690, 32'sd305821, -32'sd1362151, -32'sd633981, -32'sd732641, -32'sd3451360, -32'sd823918, 32'sd2219131, 32'sd2618866, 32'sd663969, 32'sd2275595, 32'sd2178878, -32'sd1224707, 32'sd244817, -32'sd1897364, -32'sd1600345, -32'sd948797, -32'sd2491842, -32'sd3051401, -32'sd1763374, -32'sd3006430, -32'sd2381971, -32'sd1077299, -32'sd4035534, -32'sd1133287, -32'sd1411812, 32'sd293689, -32'sd1169547, 32'sd464155, 32'sd904641, 32'sd1468348, 32'sd683898, 32'sd2867070, 32'sd250421, 32'sd1574653, 32'sd2693631, 32'sd498204, -32'sd11, 32'sd1618140, 32'sd3253090, 32'sd583667, -32'sd3108, -32'sd882716, -32'sd775141, -32'sd2662135, -32'sd3414402, -32'sd615648, -32'sd181059, -32'sd444596, -32'sd795755, -32'sd1639627, -32'sd43674, 32'sd2394243, -32'sd1040055, -32'sd277999, 32'sd59418, 32'sd151937, 32'sd0, 32'sd101353, -32'sd1083222, -32'sd4041458, -32'sd1960994, 32'sd2204715, -32'sd263179, 32'sd316209, 32'sd2354134, 32'sd572204, 32'sd1427499, 32'sd55791, 32'sd221312, -32'sd1463993, -32'sd3217070, -32'sd2404571, -32'sd1276015, 32'sd1770293, -32'sd1451285, 32'sd12550, -32'sd861854, -32'sd454576, -32'sd1406385, -32'sd3440447, -32'sd1580338, -32'sd24549, 32'sd977056, 32'sd0, 32'sd0, 32'sd0, -32'sd1488037, 32'sd975903, -32'sd559963, 32'sd1036665, 32'sd503777, -32'sd1061916, -32'sd313534, -32'sd869028, 32'sd1577895, 32'sd644050, -32'sd1449002, -32'sd785829, -32'sd209686, 32'sd286371, -32'sd4230845, -32'sd2040434, -32'sd1770646, -32'sd1736706, 32'sd1000170, 32'sd1779226, -32'sd792338, 32'sd1157716, 32'sd508267, -32'sd637637, -32'sd1641428, 32'sd0, 32'sd0, 32'sd0, 32'sd1622904, 32'sd1064034, -32'sd385222, 32'sd660801, -32'sd949776, -32'sd580034, 32'sd592814, 32'sd892465, -32'sd734981, 32'sd240304, -32'sd879541, -32'sd2947450, -32'sd697219, -32'sd846184, -32'sd3425451, -32'sd4379965, -32'sd187502, 32'sd1242481, -32'sd985530, 32'sd1016765, -32'sd1009274, 32'sd3213973, -32'sd925671, 32'sd477322, 32'sd117447, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2580479, 32'sd1531156, 32'sd1638322, -32'sd137227, 32'sd1116437, -32'sd758637, 32'sd2186221, 32'sd1524469, 32'sd1778604, -32'sd2108682, -32'sd2049753, 32'sd667126, 32'sd83190, 32'sd236021, 32'sd306778, -32'sd2113363, 32'sd373840, 32'sd893592, 32'sd417742, 32'sd2167572, 32'sd2336262, 32'sd385982, 32'sd106283, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd2764514, 32'sd875252, 32'sd3062879, 32'sd1694495, -32'sd62740, 32'sd548740, 32'sd1907802, 32'sd630949, -32'sd3019368, -32'sd1367681, 32'sd1214888, 32'sd4476973, 32'sd2028075, 32'sd2250380, -32'sd2396360, 32'sd919271, 32'sd1944455, 32'sd3912170, 32'sd2148515, 32'sd285186, 32'sd0, 32'sd0, 32'sd0, 32'sd0},
        '{32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1365263, -32'sd710634, -32'sd686209, -32'sd630769, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2600806, -32'sd1662752, -32'sd1286874, 32'sd88360, 32'sd554541, 32'sd98603, 32'sd288211, -32'sd673218, -32'sd1270899, -32'sd607567, -32'sd245725, -32'sd1900402, -32'sd2461292, -32'sd1057595, -32'sd681160, 32'sd720897, 32'sd1182277, 32'sd547256, -32'sd1737504, -32'sd1106906, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd713041, -32'sd1373902, -32'sd2205607, -32'sd800255, 32'sd347013, 32'sd1328682, 32'sd1126843, -32'sd67096, -32'sd80007, -32'sd2598311, -32'sd2208978, -32'sd3590038, -32'sd3728825, 32'sd1198119, 32'sd1035646, -32'sd1193335, 32'sd2762909, 32'sd571582, 32'sd1245563, -32'sd388510, -32'sd905060, -32'sd1054029, 32'sd95372, -32'sd2569787, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2078563, -32'sd989671, -32'sd945300, 32'sd503768, -32'sd28953, -32'sd772771, -32'sd2485765, -32'sd2200322, 32'sd663902, -32'sd1844480, 32'sd1013301, -32'sd3344259, -32'sd1940045, 32'sd518130, -32'sd2652576, -32'sd967541, 32'sd1211815, -32'sd1224083, -32'sd2773578, 32'sd815460, 32'sd177350, -32'sd256856, -32'sd365535, 32'sd733679, 32'sd313131, 32'sd0, 32'sd0, -32'sd2760314, 32'sd480769, 32'sd23070, 32'sd345321, -32'sd831999, -32'sd1107983, 32'sd1304238, -32'sd666940, 32'sd247245, -32'sd3498078, -32'sd1492687, -32'sd989739, -32'sd3368830, 32'sd264347, -32'sd392271, -32'sd45326, 32'sd2082894, 32'sd730265, -32'sd2740497, -32'sd307017, -32'sd1568282, 32'sd211028, -32'sd747313, -32'sd1463559, 32'sd1527817, 32'sd449059, -32'sd1998464, 32'sd0, 32'sd225318, -32'sd558562, 32'sd69078, 32'sd223287, 32'sd1295978, -32'sd2334657, -32'sd1799781, -32'sd285496, -32'sd1070750, -32'sd3812391, 32'sd659228, -32'sd1454644, -32'sd812131, 32'sd175611, -32'sd2454790, -32'sd3900439, -32'sd3317610, -32'sd1966435, -32'sd1241972, 32'sd2517024, -32'sd328800, -32'sd218252, -32'sd38153, -32'sd179487, 32'sd150703, 32'sd408669, 32'sd990323, 32'sd0, 32'sd369968, -32'sd835494, 32'sd221553, -32'sd1164071, -32'sd1159766, -32'sd654545, 32'sd463122, -32'sd662331, -32'sd1409083, -32'sd2870836, -32'sd219666, 32'sd54957, -32'sd3725391, -32'sd549213, -32'sd1721833, -32'sd1992537, -32'sd1087563, -32'sd2797602, 32'sd279812, -32'sd29972, 32'sd1981313, 32'sd403943, 32'sd1615375, 32'sd935625, 32'sd1256118, 32'sd986356, -32'sd336325, -32'sd1391939, -32'sd1402856, -32'sd518843, 32'sd40879, 32'sd249661, -32'sd750157, -32'sd3290130, -32'sd2325538, 32'sd631599, -32'sd3626318, 32'sd539933, 32'sd2338171, 32'sd2016611, -32'sd551854, -32'sd2266991, 32'sd995717, 32'sd1147626, -32'sd88001, 32'sd2007377, -32'sd371297, 32'sd514449, 32'sd2854214, 32'sd1910878, 32'sd1024942, -32'sd1286776, -32'sd922795, -32'sd410836, 32'sd904992, -32'sd2835518, -32'sd1238304, -32'sd2878628, -32'sd1724621, 32'sd1096173, 32'sd356506, -32'sd3215349, -32'sd2552443, -32'sd2373911, -32'sd585250, 32'sd14375, 32'sd2474036, 32'sd823913, 32'sd1373533, -32'sd2648282, -32'sd2069906, 32'sd1185466, 32'sd799986, 32'sd503324, 32'sd2244333, 32'sd2855968, 32'sd2041074, 32'sd1614731, 32'sd626624, 32'sd1199549, 32'sd541696, 32'sd228771, -32'sd254981, 32'sd510769, -32'sd836973, -32'sd639933, 32'sd473049, 32'sd2079317, -32'sd1527756, -32'sd2391820, -32'sd939155, -32'sd1707744, -32'sd126672, 32'sd1104179, 32'sd4953286, 32'sd2262602, 32'sd3593541, -32'sd984343, -32'sd964580, -32'sd99071, 32'sd1936577, 32'sd287748, 32'sd3550436, 32'sd962350, 32'sd3293778, 32'sd590963, 32'sd1330330, 32'sd3410570, 32'sd2909422, 32'sd1141191, -32'sd632801, -32'sd265220, 32'sd326112, -32'sd1930497, -32'sd615464, -32'sd205941, -32'sd3498568, -32'sd2075864, -32'sd3993784, -32'sd101051, 32'sd1757353, 32'sd2978704, 32'sd3692271, 32'sd2933481, 32'sd1498067, 32'sd1146462, -32'sd228630, -32'sd2053170, -32'sd89734, 32'sd267114, -32'sd5862, -32'sd492624, 32'sd2199613, 32'sd1464064, 32'sd957202, 32'sd1939525, -32'sd189806, 32'sd895062, 32'sd2046777, 32'sd308663, 32'sd1049400, -32'sd1326313, -32'sd3265800, -32'sd755271, -32'sd736851, -32'sd3470295, -32'sd1132373, -32'sd2320605, -32'sd30217, 32'sd153160, 32'sd2192166, 32'sd1678356, 32'sd3290743, -32'sd261836, -32'sd670186, 32'sd1672262, -32'sd2499809, -32'sd1759701, 32'sd325475, -32'sd3255999, -32'sd906874, 32'sd1702901, 32'sd3075518, 32'sd3176398, 32'sd1654230, 32'sd2242733, -32'sd196075, -32'sd2056281, -32'sd1629915, -32'sd328854, -32'sd572498, 32'sd2001004, 32'sd704393, -32'sd392834, -32'sd48506, 32'sd187736, 32'sd74392, -32'sd2918815, -32'sd1746666, 32'sd2049184, 32'sd2790762, 32'sd475603, -32'sd1248063, -32'sd2204133, -32'sd114870, -32'sd2442234, -32'sd1884894, -32'sd1235237, -32'sd380228, 32'sd1497680, 32'sd2975244, 32'sd2237043, -32'sd895892, 32'sd454491, -32'sd1119305, -32'sd169587, -32'sd512776, 32'sd1418416, -32'sd327996, -32'sd2353651, 32'sd2083752, -32'sd191506, -32'sd2568633, -32'sd622062, 32'sd2534593, -32'sd1316402, 32'sd85206, 32'sd1336768, -32'sd1156828, -32'sd543089, 32'sd339464, -32'sd711945, -32'sd2091410, -32'sd4635316, -32'sd155993, -32'sd1954357, -32'sd1703532, -32'sd1558993, -32'sd1491088, -32'sd66395, -32'sd2064665, 32'sd869758, -32'sd1077253, -32'sd2164797, -32'sd1088490, 32'sd380261, -32'sd261542, -32'sd3923174, -32'sd522516, -32'sd1399113, -32'sd2252793, -32'sd1590051, 32'sd92807, 32'sd1071350, -32'sd2404010, -32'sd1433633, 32'sd279399, 32'sd2545629, 32'sd543524, -32'sd807461, 32'sd152080, -32'sd2457838, -32'sd546685, -32'sd368757, -32'sd1915577, -32'sd3183391, -32'sd2422446, 32'sd315500, 32'sd1882819, 32'sd706736, -32'sd2690301, -32'sd2176590, -32'sd240683, -32'sd559903, 32'sd1170746, 32'sd632458, -32'sd733368, -32'sd1873338, -32'sd1617822, -32'sd131670, 32'sd2780796, -32'sd551232, -32'sd913759, 32'sd591338, 32'sd448647, 32'sd824691, -32'sd358390, -32'sd3133342, -32'sd727670, -32'sd950060, -32'sd3051199, -32'sd3484078, -32'sd799432, -32'sd1940105, -32'sd4109349, -32'sd1308928, -32'sd4592947, -32'sd3237662, -32'sd2311500, -32'sd623231, -32'sd353223, 32'sd336122, 32'sd302460, -32'sd1035210, -32'sd2074982, -32'sd2449524, -32'sd1902485, -32'sd648017, 32'sd30651, -32'sd1846213, -32'sd541520, 32'sd3043679, 32'sd2998544, -32'sd647781, -32'sd290426, -32'sd2744508, -32'sd528010, -32'sd1209811, -32'sd4463500, -32'sd3550772, -32'sd2127847, -32'sd3038721, -32'sd2554230, -32'sd3210349, -32'sd375934, -32'sd1747466, -32'sd1712078, 32'sd0, -32'sd2510469, -32'sd3283482, 32'sd531983, 32'sd884429, -32'sd1331738, 32'sd2758975, -32'sd831809, -32'sd1119624, -32'sd215586, 32'sd2259730, 32'sd3695264, 32'sd2662597, 32'sd884401, -32'sd509818, 32'sd436948, -32'sd2537899, -32'sd2137615, -32'sd3299904, -32'sd2974149, -32'sd418676, -32'sd3472129, -32'sd2421386, -32'sd2995580, -32'sd4619655, 32'sd2068695, 32'sd45435, -32'sd2385077, -32'sd1609030, -32'sd1648100, -32'sd1746900, 32'sd1987069, 32'sd240409, -32'sd1907396, 32'sd2153899, -32'sd94041, -32'sd1115967, 32'sd2123212, 32'sd1381716, 32'sd921440, 32'sd1596690, -32'sd2278710, -32'sd2100994, 32'sd648977, -32'sd679125, -32'sd1620959, -32'sd3658305, -32'sd4826325, -32'sd1774477, -32'sd971839, -32'sd1025106, -32'sd1841417, -32'sd52340, 32'sd972730, -32'sd622836, -32'sd1263613, 32'sd771715, -32'sd1570135, -32'sd709613, 32'sd597189, -32'sd1588938, -32'sd2351060, -32'sd1469180, -32'sd2172403, -32'sd2365337, -32'sd11331, 32'sd1775240, 32'sd1207586, 32'sd1739317, -32'sd1208263, -32'sd771451, -32'sd370171, 32'sd277265, -32'sd1765618, -32'sd1826821, 32'sd568099, 32'sd1367898, -32'sd77184, 32'sd203608, -32'sd527072, 32'sd883565, 32'sd32969, -32'sd867928, -32'sd5096308, 32'sd0, -32'sd926345, -32'sd564867, -32'sd1275476, -32'sd1896817, -32'sd1819038, 32'sd282737, 32'sd600915, 32'sd2539875, 32'sd2639260, 32'sd3394277, 32'sd1410501, 32'sd1140260, 32'sd842147, -32'sd1372027, 32'sd256919, -32'sd762579, 32'sd905961, 32'sd215911, 32'sd2354995, 32'sd1086230, -32'sd1077264, -32'sd703476, -32'sd511419, -32'sd105249, 32'sd764792, 32'sd675144, 32'sd106470, -32'sd1841406, -32'sd2646156, -32'sd1594996, -32'sd722214, -32'sd58842, -32'sd1400273, -32'sd351534, 32'sd1162653, 32'sd200449, 32'sd2818480, -32'sd327550, 32'sd1111914, 32'sd1318930, 32'sd1608881, -32'sd337345, -32'sd68342, 32'sd971196, 32'sd3976553, 32'sd855689, -32'sd521903, 32'sd988145, 32'sd884874, 32'sd2752043, 32'sd1862682, 32'sd2407379, -32'sd514603, 32'sd758868, 32'sd1190373, -32'sd1320623, -32'sd2491069, -32'sd1278472, 32'sd1366125, -32'sd2430197, 32'sd1428221, 32'sd1051062, -32'sd206237, -32'sd154056, 32'sd1051555, 32'sd998116, 32'sd590016, 32'sd1733412, 32'sd1966657, 32'sd1274745, 32'sd1303504, 32'sd82416, 32'sd1626631, 32'sd2767451, -32'sd538987, 32'sd572119, 32'sd411122, 32'sd2387265, 32'sd2868875, 32'sd211705, 32'sd1187541, -32'sd16020, -32'sd917950, 32'sd0, -32'sd391488, 32'sd494074, 32'sd2240126, -32'sd1512315, -32'sd767954, 32'sd237413, -32'sd1915697, 32'sd1400478, 32'sd1417699, 32'sd1248017, -32'sd400260, 32'sd851623, -32'sd676945, 32'sd2320323, -32'sd981865, 32'sd1118517, -32'sd525624, 32'sd419782, 32'sd2699451, 32'sd1535816, -32'sd590927, 32'sd465486, 32'sd287604, -32'sd512222, -32'sd1158696, -32'sd2279076, 32'sd0, 32'sd0, 32'sd0, -32'sd884, -32'sd2216425, -32'sd3219528, -32'sd1054042, -32'sd720403, -32'sd1136435, -32'sd1652429, 32'sd1067009, -32'sd1349343, 32'sd706218, 32'sd684229, 32'sd1129135, -32'sd282159, 32'sd764227, 32'sd2842012, -32'sd602549, -32'sd316006, 32'sd120419, 32'sd1234228, 32'sd32403, 32'sd847758, 32'sd1089928, 32'sd636912, -32'sd1051987, -32'sd2187508, 32'sd0, 32'sd0, 32'sd0, -32'sd1493970, -32'sd1843034, -32'sd4747356, -32'sd1221493, 32'sd232324, -32'sd3602764, -32'sd3119638, -32'sd2409796, -32'sd3143922, 32'sd222375, -32'sd2447059, -32'sd894644, -32'sd2870722, -32'sd217459, -32'sd418302, 32'sd1652400, -32'sd1771727, -32'sd853927, 32'sd587106, 32'sd1433138, -32'sd261533, 32'sd640707, 32'sd1188136, 32'sd642010, -32'sd2353888, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd2165526, -32'sd2961063, -32'sd1548089, -32'sd4749896, -32'sd1832801, -32'sd1512346, -32'sd1379976, -32'sd2609236, 32'sd483919, -32'sd247518, -32'sd486095, -32'sd177064, 32'sd486115, -32'sd331926, 32'sd2432830, 32'sd1761846, 32'sd1059674, 32'sd2650438, -32'sd154823, -32'sd204116, 32'sd1666024, -32'sd1968551, -32'sd1941850, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, 32'sd0, -32'sd1424282, -32'sd2863463, 32'sd294056, 32'sd890389, -32'sd151153, -32'sd779804, -32'sd1226322, 32'sd756274, 32'sd709877, 32'sd1819420, 32'sd613499, -32'sd1293390, -32'sd123644, -32'sd767327, 32'sd1680039, -32'sd158317, 32'sd793756, -32'sd241272, 32'sd981197, -32'sd1234592, 32'sd0, 32'sd0, 32'sd0, 32'sd0}
    };

    localparam logic signed [31:0] layer0_biases [0:15] = '{
        -32'sd1734829, -32'sd1209072, 32'sd5805217, 32'sd5674008, -32'sd887668, 32'sd1119514, -32'sd1474121, 32'sd5404959, 32'sd1786766, -32'sd2501000, 32'sd1156473, 32'sd8201868, 32'sd5205138, 32'sd5003254, -32'sd3137167, 32'sd1492095
    };

    //Layer 1: 16 inputs, 16 neurons
    localparam logic signed [31:0] layer1_weights [0:15][0:15] = '{
        '{32'sd14551974, -32'sd8798943, 32'sd292946, 32'sd6845191, -32'sd1427235, -32'sd9887541, 32'sd5281540, -32'sd831282, 32'sd1291773, 32'sd518927, -32'sd6054295, 32'sd1731567, 32'sd4505952, -32'sd1913547, 32'sd2565194, -32'sd2225839},
        '{-32'sd5641444, 32'sd689052, 32'sd11046178, 32'sd6490125, -32'sd445250, -32'sd7293743, -32'sd7491332, 32'sd7308886, 32'sd5952842, -32'sd4855419, 32'sd7163779, -32'sd8040357, -32'sd4358715, 32'sd7217979, -32'sd2446276, -32'sd5612485},
        '{32'sd243355, -32'sd7368290, 32'sd7891120, 32'sd2768636, -32'sd4305233, 32'sd4518417, 32'sd5189916, -32'sd551624, -32'sd4279691, -32'sd3713160, 32'sd5723656, 32'sd2189963, -32'sd516471, -32'sd5370851, -32'sd4431395, -32'sd4945865},
        '{-32'sd1908923, 32'sd853708, -32'sd2268401, 32'sd4862830, 32'sd10522944, -32'sd8958920, 32'sd5425849, 32'sd9985784, 32'sd4493525, -32'sd6958394, 32'sd1790382, 32'sd9660145, -32'sd2955397, -32'sd6495427, -32'sd1149624, 32'sd8227320},
        '{-32'sd4133648, -32'sd3478660, 32'sd5519982, -32'sd2046394, -32'sd5632340, 32'sd1115567, -32'sd3346367, 32'sd8028410, 32'sd5913254, -32'sd3626912, 32'sd10965598, 32'sd457997, 32'sd11529328, 32'sd7794713, 32'sd2093923, 32'sd4484687},
        '{32'sd4805818, -32'sd6928656, 32'sd8735480, 32'sd5553200, -32'sd611475, 32'sd5039170, 32'sd25458, 32'sd3107141, -32'sd8246034, 32'sd3998143, -32'sd8832742, -32'sd4369489, 32'sd6386819, 32'sd6626355, 32'sd11766915, -32'sd3211776},
        '{-32'sd4776061, 32'sd2792917, -32'sd4812052, 32'sd5404054, 32'sd7374238, -32'sd5396076, -32'sd9669680, 32'sd3766422, 32'sd5841990, 32'sd6440200, -32'sd2312734, -32'sd4715548, 32'sd310332, -32'sd4154852, 32'sd6181791, -32'sd5973277},
        '{32'sd7394395, 32'sd1682734, -32'sd2642761, -32'sd520147, -32'sd7361606, 32'sd6520362, -32'sd9642472, 32'sd3657371, -32'sd6203221, -32'sd8145107, 32'sd2944626, 32'sd758497, -32'sd3405206, -32'sd4833031, 32'sd5381977, 32'sd5538567},
        '{32'sd8712578, 32'sd5372013, 32'sd4193343, -32'sd4664031, 32'sd5706593, -32'sd6883430, -32'sd7950027, 32'sd2769268, -32'sd5519674, 32'sd8346241, -32'sd990468, 32'sd5877990, -32'sd868217, 32'sd5109713, -32'sd5793989, -32'sd6448052},
        '{32'sd2497540, 32'sd5113402, 32'sd1254212, -32'sd7972482, 32'sd8992488, 32'sd3881486, 32'sd12067483, 32'sd8107015, 32'sd1395714, -32'sd906654, 32'sd1258435, -32'sd513515, -32'sd2403447, 32'sd4870839, -32'sd5652442, 32'sd10041939},
        '{32'sd9883420, 32'sd8045570, -32'sd8320550, 32'sd2242885, 32'sd3904257, 32'sd7029139, 32'sd3080426, -32'sd304871, 32'sd3991427, 32'sd2388533, 32'sd6249366, 32'sd6870025, 32'sd15266529, 32'sd5137249, -32'sd8018778, -32'sd4016919},
        '{-32'sd4440603, 32'sd7867995, 32'sd255250, 32'sd7008517, 32'sd6411843, 32'sd7316098, 32'sd1014582, -32'sd4406063, -32'sd11063200, 32'sd2232350, 32'sd338632, 32'sd1695665, -32'sd6788053, -32'sd750517, -32'sd4797024, -32'sd2017719},
        '{32'sd360316, 32'sd3462482, 32'sd1759999, -32'sd2445550, 32'sd9424739, 32'sd4481214, 32'sd4462663, -32'sd5809464, -32'sd9761651, 32'sd11479374, 32'sd6414297, -32'sd5118158, 32'sd2875739, 32'sd5433237, 32'sd9232400, 32'sd2899887},
        '{-32'sd2627208, 32'sd2756578, 32'sd2396463, 32'sd2178450, -32'sd8435827, 32'sd5549622, 32'sd5127911, -32'sd5455895, 32'sd5191184, -32'sd6775594, 32'sd2725696, -32'sd5134527, -32'sd1749399, 32'sd4701941, -32'sd6188660, 32'sd9530594},
        '{-32'sd4806341, -32'sd2263787, 32'sd3043880, -32'sd1624042, 32'sd1789423, 32'sd3541935, -32'sd572683, 32'sd6743612, 32'sd8332344, 32'sd7754530, 32'sd7977777, -32'sd5235007, -32'sd3749285, -32'sd4381081, 32'sd1077565, 32'sd2720220},
        '{32'sd1496811, -32'sd3864454, 32'sd1902677, 32'sd8385416, -32'sd5946639, 32'sd6586459, 32'sd5460532, -32'sd9681993, -32'sd3344910, 32'sd418129, -32'sd165180, -32'sd6624973, 32'sd5430495, -32'sd8447742, 32'sd4936132, 32'sd2406989}
    };

    localparam logic signed [31:0] layer1_biases [0:15] = '{
        32'sd8287540, 32'sd5023592, 32'sd1901070, 32'sd3191750, 32'sd9781365, 32'sd3985504, 32'sd586070, -32'sd5661924, -32'sd2105236, -32'sd5198851, 32'sd4231044, 32'sd2608879, 32'sd1528332, 32'sd4163394, -32'sd2965845, 32'sd5511686
    };

    //Layer 2: 16 inputs, 10 neurons
    localparam logic signed [31:0] layer2_weights [0:9][0:15] = '{
        '{-32'sd4318163, -32'sd4611655, 32'sd10123105, -32'sd9539038, 32'sd4722300, -32'sd7509887, -32'sd4667472, 32'sd3879960, -32'sd6403890, -32'sd5662311, 32'sd6635676, 32'sd7697585, 32'sd2505828, -32'sd3053363, 32'sd11425550, -32'sd2030767},
        '{-32'sd5444574, 32'sd5832410, -32'sd1225713, -32'sd11261693, -32'sd1584628, 32'sd6212451, 32'sd6516145, -32'sd9702844, -32'sd7013272, 32'sd5215876, -32'sd4836841, -32'sd1280852, 32'sd12473685, 32'sd7960592, -32'sd5414117, -32'sd6678988},
        '{-32'sd8012576, 32'sd6176376, -32'sd5777525, -32'sd8222173, 32'sd4748876, -32'sd1627500, 32'sd3821134, -32'sd6544138, -32'sd1666808, 32'sd6436123, 32'sd8328140, -32'sd6574582, -32'sd4032701, 32'sd9393907, -32'sd7605966, 32'sd7275819},
        '{32'sd9481163, 32'sd3502548, -32'sd10142244, -32'sd8640973, -32'sd2239762, 32'sd5068083, -32'sd4047206, -32'sd1710046, 32'sd11302385, 32'sd1007631, 32'sd4609549, 32'sd9237407, -32'sd749673, -32'sd602077, -32'sd2990599, -32'sd3767472},
        '{32'sd836504, 32'sd11323112, 32'sd6578982, 32'sd104612, 32'sd23025, 32'sd7293273, 32'sd9288221, 32'sd5691781, -32'sd6453288, -32'sd7297123, -32'sd11517685, -32'sd3853045, -32'sd2739861, 32'sd689629, 32'sd8081460, -32'sd5143777},
        '{32'sd4972419, 32'sd1869411, -32'sd3490418, 32'sd8731159, -32'sd17483841, -32'sd2069134, -32'sd3969863, 32'sd12208686, -32'sd2972327, 32'sd7109885, 32'sd1559036, 32'sd7052718, 32'sd1990216, 32'sd2081479, 32'sd2519251, 32'sd4101761},
        '{-32'sd12281724, -32'sd1712460, 32'sd1198866, 32'sd2336754, -32'sd1871897, -32'sd6966698, 32'sd6982215, -32'sd5341681, -32'sd160740, 32'sd7136881, 32'sd337471, -32'sd1550778, 32'sd1199484, -32'sd6927997, 32'sd8517064, -32'sd6879549},
        '{-32'sd4421998, 32'sd4317336, 32'sd2604887, -32'sd15620699, 32'sd4041028, 32'sd11063641, -32'sd1373638, -32'sd1668790, 32'sd5337578, -32'sd11139258, 32'sd2403772, 32'sd6546668, -32'sd2084969, -32'sd2083903, -32'sd883909, 32'sd8191265},
        '{-32'sd8561431, -32'sd6450089, -32'sd234462, 32'sd8904848, 32'sd9862301, -32'sd303294, -32'sd7364111, 32'sd2949855, 32'sd9221217, 32'sd1502885, 32'sd125126, -32'sd2967391, -32'sd706335, -32'sd9073348, -32'sd3703673, 32'sd2562391},
        '{32'sd12244459, 32'sd802908, -32'sd973094, 32'sd1262986, -32'sd4018186, 32'sd1656219, 32'sd9979454, 32'sd2797873, 32'sd1313497, 32'sd1429164, -32'sd617982, -32'sd3126450, -32'sd4969796, -32'sd941258, -32'sd6283163, 32'sd10703601}
    };

    localparam logic signed [31:0] layer2_biases [0:9] = '{
        32'sd4147116, -32'sd4517701, -32'sd9414776, 32'sd8640457, -32'sd6157512, 32'sd4199429, 32'sd483663, 32'sd5683063, 32'sd5311282, 32'sd3319070
    };


    //Intermediate outputs
    logic signed [31:0] layer0_out [0:15];
    logic signed [31:0] layer1_out [0:15];


    //Instantiate Layers
    //Layer 0
    layer #(
        .NEURONS(16),
        .PREV_LAYER_OUTPUTS(784)
    ) layer0 (
        .data_inputs(data_inputs),
        .weights(layer0_weights),
        .biases(layer0_biases),
        .data_outputs(layer0_out)
    );

    //Layer 1
    layer #(
        .NEURONS(16),
        .PREV_LAYER_OUTPUTS(16)
    ) layer1 (
        .data_inputs(layer0_out),
        .weights(layer1_weights),
        .biases(layer1_biases),
        .data_outputs(layer1_out)
    );

    //Layer 2
    layer #(
        .NEURONS(10),
        .PREV_LAYER_OUTPUTS(16)
    ) layer2 (
        .data_inputs(layer1_out),
        .weights(layer2_weights),
        .biases(layer2_biases),
        .data_outputs(data_outputs)
    );



    // Predicted class logic
    always_comb begin
        logic signed [31:0] max_val;
        max_val = data_outputs[0];
        predicted_class = '0;

        for (int i = 1; i < OUTPUTS; i++) begin
            if (data_outputs[i] > max_val) begin
                max_val = data_outputs[i];
                predicted_class = i[OUTPUT_IDX_BITS-1:0];
            end
        end
    end
endmodule
