module mlp_neural_net #(
    parameter int INPUTS  = 784,
    parameter int OUTPUTS = 10
) (
    input  logic signed [31:0] data_inputs  [0:INPUTS-1],
    output logic signed [31:0] data_outputs [0:OUTPUTS-1]
);

    //Layer 0: 784 inputs, 128 neurons
    localparam logic signed [31:0] layer0_weights [0:127][0:784] = '{
        '{32'sd1.718359258788821e-125, 32'sd5.352691656835491e-118, 32'sd-5.981172718220442e-126, 32'sd6.872192727514316e-122, 32'sd-1.64319177998815e-116, 32'sd7.357757788869089e-117, 32'sd-2.5306859728395336e-120, 32'sd6.3509356256817e-121, 32'sd2.4963554141764615e-126, 32'sd-5.061560824904401e-119, 32'sd1.083457284587331e-121, 32'sd5.56813996720011e-117, 32'sd-0.044733315826406314, 32'sd0.07138973985590737, 32'sd0.0782794975074838, 32'sd0.09028033667838985, 32'sd1.792212656138361e-128, 32'sd-7.122717776858756e-115, 32'sd7.288895118796694e-124, 32'sd-1.106392134437505e-118, 32'sd1.0185964871778448e-118, 32'sd-2.6477611382547744e-123, 32'sd-5.034351332250756e-119, 32'sd-7.467908727265815e-115, 32'sd2.764207270337301e-126, 32'sd-1.0403406299105053e-120, 32'sd1.374403834679118e-115, 32'sd-1.1018801344974543e-119, 32'sd1.4061623974554275e-127, 32'sd1.9284887475232276e-120, 32'sd-1.6781583397281288e-126, 32'sd-4.8221724182501905e-123, 32'sd0.019500238346360492, 32'sd0.026674336387622385, 32'sd0.12045596740893666, 32'sd0.03950927601080809, 32'sd0.07439853521001825, 32'sd0.12300041500547405, 32'sd0.11105884626390772, 32'sd0.15497991343617998, 32'sd0.04343070311165017, 32'sd0.008451869486807137, 32'sd0.016657795132763286, 32'sd0.027521540240186607, 32'sd0.08225166051362584, 32'sd0.0008608706514846763, 32'sd0.05208076293782294, 32'sd-0.032328349908395795, 32'sd-0.009567912479530474, 32'sd-0.000683928161037325, 32'sd0.03588221240025074, 32'sd0.03537256514622789, 32'sd-2.8054809990113787e-120, 32'sd-1.5712040768312306e-119, 32'sd2.6160119491561765e-121, 32'sd3.402728175840336e-117, 32'sd-1.6188546420388234e-115, 32'sd1.9236475896850427e-124, 32'sd0.06641593168862925, 32'sd0.027708487220609843, 32'sd-0.03808247285940734, 32'sd-0.04771950302679152, 32'sd0.0997096799940716, 32'sd0.012300189369226926, 32'sd0.039077477810300194, 32'sd-0.0446413515796236, 32'sd0.11769600906610031, 32'sd0.05181495371475874, 32'sd-0.05529588716210715, 32'sd-0.002472529169550334, 32'sd0.021913491451790695, 32'sd0.08024811852527886, 32'sd0.07122935337011863, 32'sd0.17272219281681866, 32'sd0.21408856366177303, 32'sd0.17847565613732896, 32'sd0.02267712394555068, 32'sd0.10907897437963913, 32'sd0.037165765178919445, 32'sd0.0456868720958468, 32'sd0.09443811789195836, 32'sd0.02985537505387772, 32'sd-2.582181988064221e-121, 32'sd8.796553700146387e-127, 32'sd-9.202144384336723e-125, 32'sd-4.759071254472596e-123, 32'sd-0.08615545911131096, 32'sd0.006212736694240674, 32'sd0.005072789937227223, 32'sd0.0364938165855177, 32'sd-0.039549040139709515, 32'sd0.013435490766974595, 32'sd-0.02802730618723184, 32'sd-0.03067014469105056, 32'sd0.06091970558426617, 32'sd0.06992112720989216, 32'sd0.016935162628421055, 32'sd-0.04611960738524131, 32'sd-0.0165242401162588, 32'sd-0.07302127218317021, 32'sd-0.03475825534438184, 32'sd0.08914899080253146, 32'sd0.03343860201753874, 32'sd-0.12523696468263762, 32'sd0.0890617344456426, 32'sd0.05434924224119682, 32'sd0.00769539932784079, 32'sd0.03325538838544562, 32'sd0.09231276464151, 32'sd7.95139168108201e-06, 32'sd0.02910721928105544, 32'sd6.426587760093643e-117, 32'sd4.222124324955341e-118, 32'sd0.006953158847783545, 32'sd0.032329718399061326, 32'sd-0.017306009760915887, 32'sd-0.05785589994012573, 32'sd0.09042980373265808, 32'sd-0.11995518398177646, 32'sd-0.11757781955284743, 32'sd-0.07700200671679286, 32'sd-0.17123226563859387, 32'sd-0.046241495987105016, 32'sd-0.05852868659739165, 32'sd-0.2110213976540472, 32'sd-0.13564057006553673, 32'sd-0.133799775216942, 32'sd0.08197458548237924, 32'sd-0.07725518699731826, 32'sd0.045410033741045526, 32'sd0.09666234768244461, 32'sd0.11239521775161113, 32'sd0.0843636419310122, 32'sd0.05247215396053713, 32'sd0.001050923667632968, 32'sd0.0838154377474873, 32'sd-0.01503355792213817, 32'sd0.06920290669490736, 32'sd0.012898520853377934, 32'sd0.07897141437262753, 32'sd5.875284069511495e-124, 32'sd0.044587069081651436, 32'sd0.008417474266953065, 32'sd-0.04903023917361535, 32'sd-0.07673745675411367, 32'sd-0.07669051170145848, 32'sd-0.024291933423423742, 32'sd-0.14460485099406153, 32'sd-0.09545545651155164, 32'sd-0.10682463076762638, 32'sd-0.047719738278823656, 32'sd-0.07250169098191687, 32'sd-0.2274508113306219, 32'sd-0.04498848653093782, 32'sd-0.06030115010844043, 32'sd0.015555492353489062, 32'sd-0.10407787603035136, 32'sd0.03630742840953154, 32'sd-0.0812705839132061, 32'sd0.06540158318187787, 32'sd0.14243802715629494, 32'sd0.008168292406141605, 32'sd0.04027704116466655, 32'sd0.0006338808914194032, 32'sd0.018173113444681414, 32'sd-0.043584363466779893, 32'sd-0.07619490395690907, 32'sd0.011301323721898172, 32'sd-1.0149134038311193e-114, 32'sd0.04140621830071325, 32'sd-0.059250764987931547, 32'sd-0.0032036535259419166, 32'sd-0.037327022793928154, 32'sd0.06777417463233981, 32'sd-0.022122283156852815, 32'sd-0.012611903452108405, 32'sd-0.17441890443331337, 32'sd-0.15982719900602785, 32'sd-0.09635943544244556, 32'sd-0.14726795694204864, 32'sd0.08417725142084292, 32'sd-0.011031606504048722, 32'sd-0.006829324587475372, 32'sd0.024259158493155637, 32'sd-0.1687982324983564, 32'sd-0.03933437996122107, 32'sd0.017202640113479314, 32'sd0.12460958554841892, 32'sd0.12334048938409586, 32'sd0.02341811170893514, 32'sd0.10085929935316199, 32'sd-0.09711052088773467, 32'sd0.06296067841909528, 32'sd0.005436348825691257, 32'sd0.03513807874604642, 32'sd-0.004062318741889441, 32'sd0.024186095878630475, 32'sd-0.0024432278866041543, 32'sd-0.0409923722516873, 32'sd0.032903250548938355, 32'sd-0.01228486069542567, 32'sd-0.042469578967466295, 32'sd-0.09242852021031414, 32'sd-0.033230605548561276, 32'sd-0.13190528065781423, 32'sd-0.09399495627623945, 32'sd-0.038453764516060356, 32'sd0.03709526222416514, 32'sd0.0057017404768128065, 32'sd0.15380391629801468, 32'sd-0.04253971491855391, 32'sd-0.14394064184984195, 32'sd0.001835446824402586, 32'sd0.027246828482557855, 32'sd0.1785676029066929, 32'sd0.10918291935905863, 32'sd0.034121219524076325, 32'sd0.057932537722494674, 32'sd0.2030824567463459, 32'sd0.08765452068780455, 32'sd0.051811920222777585, 32'sd-0.0008429086808202013, 32'sd-0.039171975492325976, 32'sd-0.0034338548250193945, 32'sd0.023747522807268478, 32'sd0.04577342121637697, 32'sd0.00911586063293625, 32'sd-0.007042234557891874, 32'sd0.06960162292027626, 32'sd0.010210274999383671, 32'sd-0.02522078395102724, 32'sd-0.035952159023693, 32'sd-0.09121915033367717, 32'sd-0.056177255236624396, 32'sd-0.14486690053643683, 32'sd-0.08159551577150895, 32'sd0.18508289627334384, 32'sd0.11531157385682049, 32'sd0.0724595902226622, 32'sd0.03671727072996815, 32'sd0.10992042266388762, 32'sd0.03830134943682187, 32'sd0.09397196861167666, 32'sd-0.0022413321107604047, 32'sd0.14599416661710632, 32'sd0.03258891281672299, 32'sd0.13003299744714003, 32'sd0.11761276296856685, 32'sd0.1778333620881442, 32'sd0.11289909846694772, 32'sd0.024106169720010666, 32'sd0.05731692823349699, 32'sd0.031123858431432522, 32'sd0.04600171696171064, 32'sd0.0861060731254349, 32'sd0.012853048663274297, 32'sd0.11253068063921771, 32'sd0.08944630352333698, 32'sd0.08151043508325896, 32'sd-0.04761595874705893, 32'sd-0.13417068739472587, 32'sd-0.1680669580666128, 32'sd-0.015927941427631032, 32'sd0.07151025509834642, 32'sd0.157345165465788, 32'sd0.08243568554345754, 32'sd0.20134819878418125, 32'sd0.09494825635752581, 32'sd-0.008607717971720422, 32'sd0.014391381683022952, 32'sd0.07701544307349248, 32'sd0.02223947606322228, 32'sd0.10765659116846206, 32'sd-2.4744871338575764e-06, 32'sd-0.011081179983202885, 32'sd0.05752733737254148, 32'sd0.11169900423293402, 32'sd0.07139052023769046, 32'sd0.0015221308578240516, 32'sd-0.07874227681526015, 32'sd-0.0625505620621783, 32'sd-0.029342996618544916, 32'sd-0.010698760386126056, 32'sd-0.017601004282806247, 32'sd0.04638639028877733, 32'sd0.14987089271606752, 32'sd0.06751029732660421, 32'sd-0.10375494108883404, 32'sd-0.08333347118825758, 32'sd0.012030181426586694, 32'sd0.011546016387755934, 32'sd0.02162377520497482, 32'sd0.06493512634300123, 32'sd0.13517717013970132, 32'sd0.12476486376722894, 32'sd0.08845903895540498, 32'sd-0.0041492073343228734, 32'sd-0.01993739211579879, 32'sd-0.020577889179262895, 32'sd-0.02522368336575963, 32'sd0.05988898626992748, 32'sd0.07096775943451498, 32'sd0.09693290157244468, 32'sd0.05535754513468415, 32'sd-0.052737031112180595, 32'sd0.037329301507425236, 32'sd0.07125356659404644, 32'sd0.03861316835619037, 32'sd0.04058185448696098, 32'sd-0.05613585114503191, 32'sd-0.09698225643942422, 32'sd-0.07059789969623324, 32'sd0.16079774875746405, 32'sd-0.04261304070086725, 32'sd0.08804886877698595, 32'sd0.10277976236203913, 32'sd0.15261570236262548, 32'sd-0.005764874734898806, 32'sd-0.058668018882285906, 32'sd0.13250158870443338, 32'sd0.0959822718309848, 32'sd0.054467080162340614, 32'sd0.0037129391120942585, 32'sd-0.06129442981291967, 32'sd-0.17114210022934578, 32'sd-0.24268950497487313, 32'sd-0.1435658336103055, 32'sd-0.05995915374828455, 32'sd0.00022645673183508967, 32'sd-0.15825371914244496, 32'sd-0.16308613268499475, 32'sd-0.07837840637326932, 32'sd-0.04558416224855497, 32'sd-0.07340522998563437, 32'sd-0.014715236992759867, 32'sd-0.019076330943666477, 32'sd0.0009268001348865947, 32'sd-0.05670355931520637, 32'sd-0.03170989692815663, 32'sd0.0891961861881832, 32'sd0.03692579537105088, 32'sd0.0013311709104404188, 32'sd0.03972816119778427, 32'sd0.0962444650030477, 32'sd0.1254824764274859, 32'sd0.08797250797803138, 32'sd-0.08133201608471836, 32'sd0.05830310563468872, 32'sd0.011593117857045719, 32'sd0.05092137409582241, 32'sd-0.09398553675631253, 32'sd-0.09170856791707188, 32'sd-0.26874108786350603, 32'sd-0.31256771291187324, 32'sd-0.1580062201976458, 32'sd-0.0832283160986729, 32'sd-0.0890905293226045, 32'sd-0.06977250213487264, 32'sd-0.09682179237122797, 32'sd-0.08734406304218954, 32'sd0.07996245850433917, 32'sd0.05304075772807813, 32'sd-0.0944209629952103, 32'sd0.011912870164227372, 32'sd0.008249546493005296, 32'sd0.01162539061845527, 32'sd-0.009954551987266283, 32'sd0.020683513900164274, 32'sd-0.07742661283441542, 32'sd0.010351993660177555, 32'sd0.10689151940694487, 32'sd0.09812389670792934, 32'sd-0.08816972217643718, 32'sd-0.021429910699209957, 32'sd0.03812890311719934, 32'sd-0.04204480467693608, 32'sd0.06574981027093264, 32'sd-0.057927466261954184, 32'sd-0.014872291277404007, 32'sd-0.024693871180371616, 32'sd-0.23445131059440602, 32'sd-0.13284738737361332, 32'sd-0.08090739588651952, 32'sd-0.12878222167931114, 32'sd-0.1660844221105122, 32'sd-0.14186254417496388, 32'sd0.08202990064613463, 32'sd0.08926956982396485, 32'sd0.027377284889650008, 32'sd-0.033385785342677624, 32'sd-0.11459959195790667, 32'sd0.08042575744713977, 32'sd-0.020923208513274647, 32'sd0.040201487165755403, 32'sd0.04599592274407219, 32'sd-0.03066701855767927, 32'sd0.0010400022487846781, 32'sd0.029512334450788064, 32'sd-0.0738853568575191, 32'sd0.02730422796899923, 32'sd-0.10826411741961431, 32'sd-0.0233441724996001, 32'sd0.05356686224984623, 32'sd-0.05813870671906158, 32'sd-0.01930332852865692, 32'sd-0.16932395257474506, 32'sd-0.149447441112215, 32'sd-0.06402992811779942, 32'sd-0.21252071216668203, 32'sd0.08745567378103893, 32'sd-0.04348585812860992, 32'sd0.012735695142692318, 32'sd0.0007680344578633836, 32'sd0.03928901827470098, 32'sd0.029285323688704474, 32'sd0.06425530439476539, 32'sd-0.035483569269287446, 32'sd-0.0426976137955557, 32'sd-0.021649327128890786, 32'sd0.06877893871940849, 32'sd-0.01837535156324155, 32'sd-0.06990442386743412, 32'sd-0.0635638055634053, 32'sd-0.0367990479739152, 32'sd0.07027205670449638, 32'sd0.06476252799026412, 32'sd-0.09497186004712423, 32'sd0.03567163726751521, 32'sd-0.037815552215226235, 32'sd-0.052820988458599, 32'sd-0.050384348123584416, 32'sd0.008504884089740568, 32'sd0.035843696662410114, 32'sd0.022195729444583243, 32'sd-0.05448556677112039, 32'sd-0.02329144460373382, 32'sd-0.06507031339549114, 32'sd0.21999187507027188, 32'sd0.12901129967983208, 32'sd-0.011501342042475118, 32'sd-0.09645336358172923, 32'sd0.10864669936457366, 32'sd0.006636906384356382, 32'sd0.046307030443972476, 32'sd0.11197127900832446, 32'sd-0.02827709116422071, 32'sd0.11875885258926869, 32'sd0.024835849165619768, 32'sd0.026930810766857324, 32'sd-0.012013431818399077, 32'sd-0.0591903214670288, 32'sd-0.07502464283578934, 32'sd-0.015566483466690182, 32'sd-0.014222331591922644, 32'sd-0.03029277018720987, 32'sd0.07696725840701765, 32'sd0.10930062644380407, 32'sd0.06551478057661042, 32'sd-0.02055490556152656, 32'sd-0.005626398351916428, 32'sd0.18872101766096516, 32'sd-0.05606556599803275, 32'sd0.09028719848219423, 32'sd-0.01304996102932319, 32'sd0.011127716202012531, 32'sd0.14827341418839665, 32'sd0.11357462150037058, 32'sd-0.004104132282585726, 32'sd-0.21695436786142897, 32'sd0.03490744353168842, 32'sd0.031166187581966067, 32'sd0.008471551333240375, 32'sd0.09154753838778343, 32'sd0.10447506950045705, 32'sd0.08656921335170358, 32'sd0.06537064981197675, 32'sd3.241390213266897e-126, 32'sd-0.016483866567762708, 32'sd0.04183065485406338, 32'sd0.03331771110172046, 32'sd-0.05971426819643531, 32'sd-0.06421221383067877, 32'sd-0.004928815247242626, 32'sd0.08360035160248003, 32'sd0.08398473200827017, 32'sd0.05888368868604785, 32'sd0.011725050561318989, 32'sd-0.03867504463207322, 32'sd-0.08004668140624831, 32'sd-0.10070292670424869, 32'sd0.014488616663797532, 32'sd0.16296211687693296, 32'sd0.049364753646027056, 32'sd0.06526103014706548, 32'sd0.006403067929518191, 32'sd-0.04452705081011293, 32'sd-0.09756005601063143, 32'sd-0.0033194199085889203, 32'sd0.0880177606418452, 32'sd0.13976563066308528, 32'sd0.05809331078123304, 32'sd0.024114042785496913, 32'sd0.030917477295020448, 32'sd-0.009582168857986326, 32'sd0.05282445910248048, 32'sd0.02470692532351081, 32'sd0.03838707556685337, 32'sd0.0737491317615476, 32'sd-0.05837101565670729, 32'sd0.05219356865160113, 32'sd0.04263921303359327, 32'sd0.1851145065522712, 32'sd0.12131318394588436, 32'sd-0.044977684456623215, 32'sd-0.10598135719967006, 32'sd-0.219303221338139, 32'sd-0.05935919409208744, 32'sd-0.1624341344546915, 32'sd0.02632051239587395, 32'sd0.09887040366532401, 32'sd0.21391313439200924, 32'sd0.06659664063489716, 32'sd0.02576857092360537, 32'sd-0.125271621560759, 32'sd-0.13604616575395925, 32'sd-0.10020570427545196, 32'sd0.02286572874653604, 32'sd0.06657755655849636, 32'sd-0.008330104036814213, 32'sd-0.09173162458454194, 32'sd-0.013997826384405238, 32'sd0.009152480654274733, 32'sd0.00365010644951575, 32'sd0.014866650667249263, 32'sd0.11091279137990961, 32'sd-0.07728173331157925, 32'sd-0.060374520157598775, 32'sd0.041197495704949696, 32'sd0.11876067804678662, 32'sd0.054034725257430964, 32'sd0.10652745468240007, 32'sd-0.06498304798948505, 32'sd-0.09901878089581824, 32'sd-0.0947305882703435, 32'sd0.018606797446216065, 32'sd-0.024587274667160115, 32'sd-0.028332332879723882, 32'sd0.12326544427395493, 32'sd0.13010240185733354, 32'sd-0.03158861144284102, 32'sd-0.043009379983152615, 32'sd-0.2354443103885305, 32'sd-0.1414346382475937, 32'sd-0.03591021267681179, 32'sd0.1692281090706862, 32'sd0.04090469952210023, 32'sd-0.03748396039281616, 32'sd-0.1014444729447252, 32'sd-0.08872421196909394, 32'sd-0.03392815820342156, 32'sd1.690716685968342e-123, 32'sd0.008847105913562145, 32'sd0.05676289868092535, 32'sd0.006506573012114852, 32'sd-0.02564092491693074, 32'sd0.09987448947525483, 32'sd0.11903849000733009, 32'sd0.0990031441282666, 32'sd0.1840584451725767, 32'sd0.05968709837926098, 32'sd0.0902819346137521, 32'sd0.0897830229335608, 32'sd0.08462075955119203, 32'sd0.07817256737980306, 32'sd-0.1031478518096292, 32'sd-0.011905524830943178, 32'sd-0.06280479913477593, 32'sd-0.06820390745835306, 32'sd-0.07858446723889548, 32'sd-0.045764511550922385, 32'sd-0.12816915742228757, 32'sd-0.052297756929253425, 32'sd0.07099893012180178, 32'sd-0.02663595984055149, 32'sd-0.00720097033305187, 32'sd-0.12868930061154712, 32'sd-0.061531040226598596, 32'sd0.029879368398413302, 32'sd-0.010925675374530189, 32'sd0.011445646399885559, 32'sd0.014658559411861857, 32'sd0.08296953234764474, 32'sd0.10158877518043993, 32'sd0.01892400793224865, 32'sd-0.021371063788497964, 32'sd0.07699846938089394, 32'sd0.0061916728847575585, 32'sd0.06839216265091887, 32'sd0.020678484409889588, 32'sd0.00476133139503208, 32'sd0.09016152573482575, 32'sd0.13421727059445482, 32'sd-0.06077595351059873, 32'sd-0.04984694721585075, 32'sd-0.04976757085152137, 32'sd0.057676312119561327, 32'sd-0.19681792099291093, 32'sd-0.0668069222643008, 32'sd-0.07736514198189193, 32'sd-0.0775973652928886, 32'sd0.009266588135038856, 32'sd-0.05346307310353452, 32'sd-0.1307397965488505, 32'sd-0.006425144126769735, 32'sd-0.045455826543742237, 32'sd0.04998968102038654, 32'sd0.03719906558475337, 32'sd0.003790073294228524, 32'sd0.008240775477716997, 32'sd0.12346810992009176, 32'sd-0.011974493651207061, 32'sd-0.07557726071790115, 32'sd0.10816339302287387, 32'sd0.005315685020134833, 32'sd-0.04050283572790517, 32'sd-0.03340656042456081, 32'sd0.14806531723267688, 32'sd-0.007458619154532146, 32'sd0.05317264420871694, 32'sd0.046986851638424317, 32'sd0.011081187341493095, 32'sd-0.04534279655254403, 32'sd0.0008917379686243861, 32'sd0.07839647831217382, 32'sd-0.0731777707833482, 32'sd0.0006724518008703196, 32'sd0.01295152133218886, 32'sd-0.05662229905185923, 32'sd0.10793629913343555, 32'sd0.046056948749794546, 32'sd-0.08301448790598068, 32'sd-0.09864819612126273, 32'sd-0.020575528394738547, 32'sd0.0436794204858755, 32'sd1.486500455606385e-125, 32'sd0.04525623316579433, 32'sd-0.0044167325803785035, 32'sd0.003695967622870799, 32'sd0.09592648772001985, 32'sd-0.06939669636275622, 32'sd0.19731431903369448, 32'sd0.16241504670087523, 32'sd0.10753616963693165, 32'sd0.022650721097135694, 32'sd0.04410575324820312, 32'sd0.055579007100040385, 32'sd0.13261768228070103, 32'sd0.08476610717514345, 32'sd0.059326853882248794, 32'sd-0.03725114882480032, 32'sd-0.06955235562690132, 32'sd-0.15275875725861507, 32'sd-0.08138018436730005, 32'sd-0.09074762716877129, 32'sd0.043401287919841096, 32'sd-0.01101218399534158, 32'sd0.09561985851060513, 32'sd-0.006812044062160761, 32'sd-0.11769587381698944, 32'sd0.04250182401576722, 32'sd-0.07577034738847437, 32'sd-4.360196852066068e-124, 32'sd3.9087675798337753e-118, 32'sd-2.0260565478313906e-117, 32'sd0.022948530216334504, 32'sd-0.0543908980825305, 32'sd-0.012464557458645604, 32'sd0.012025027559823903, 32'sd0.06060289257384895, 32'sd0.1579580394977839, 32'sd0.040113875860091505, 32'sd-0.01852768469147327, 32'sd0.003435313841812341, 32'sd0.06860710794728621, 32'sd0.014027267133333356, 32'sd-0.047622974863876066, 32'sd-0.1308086566359836, 32'sd0.015037993201434776, 32'sd0.06646855504084788, 32'sd0.057427683078665616, 32'sd-0.030164516198014205, 32'sd0.07361335665877003, 32'sd-0.015300938254468892, 32'sd-0.04352689977954262, 32'sd-0.09828755471880773, 32'sd0.06405961354038567, 32'sd-0.1330060368317141, 32'sd0.011650859124759478, 32'sd0.0031215185390541947, 32'sd8.812922070816881e-126, 32'sd-8.606790188670193e-122, 32'sd-9.303971943909326e-121, 32'sd0.016003968834440583, 32'sd0.018473581379641724, 32'sd0.001438236539607211, 32'sd-0.023756753382279082, 32'sd-0.012730376625485191, 32'sd-0.0039471909935388525, 32'sd-0.16079817187089768, 32'sd0.07466896652305527, 32'sd0.12049212721492918, 32'sd0.16365163453383708, 32'sd0.05074104349504579, 32'sd0.009988911064153715, 32'sd-0.08167775890932158, 32'sd0.03105571953416685, 32'sd0.021582137378358655, 32'sd0.12663497763587703, 32'sd0.10013265182662717, 32'sd0.16601880180369635, 32'sd0.12848090212042926, 32'sd0.09524787952052637, 32'sd0.0016388729669003844, 32'sd0.03238096112063616, 32'sd0.015264010079141218, 32'sd0.008253816849814995, 32'sd0.0026852032753487366, 32'sd6.869342007510948e-124, 32'sd5.175852121477398e-118, 32'sd2.312098653231584e-120, 32'sd-2.015731156148913e-127, 32'sd0.06815846201357159, 32'sd-0.05469880873912278, 32'sd0.0021778980429898467, 32'sd-0.12109740691596885, 32'sd0.05925234921025055, 32'sd-0.06766607944078136, 32'sd0.019344667924492714, 32'sd-0.0006364754684033419, 32'sd0.14162187128629192, 32'sd0.2132848883982843, 32'sd0.14524383824326909, 32'sd-0.04977725510573775, 32'sd0.09921180236119588, 32'sd-0.0054755438648665285, 32'sd-0.12101725915275961, 32'sd-0.06286359213820181, 32'sd-0.12233558125407179, 32'sd-0.03688259043216213, 32'sd0.03280593654978061, 32'sd-0.028131391814418323, 32'sd0.05939816818847722, 32'sd0.007162963445862385, 32'sd0.032147998571364855, 32'sd2.326305137136481e-114, 32'sd-7.848840622951873e-119, 32'sd1.278137314199453e-122, 32'sd-4.164238697286537e-126, 32'sd3.528734267141213e-122, 32'sd-2.1704408015465406e-127, 32'sd0.08703652011738165, 32'sd0.07349697834033303, 32'sd0.01709594351797168, 32'sd-0.013676718581245475, 32'sd0.011697718773427264, 32'sd0.08971775520484915, 32'sd-0.056532476667820214, 32'sd0.07299715590116364, 32'sd0.12088144944025796, 32'sd0.02837125591322104, 32'sd0.12683026467171526, 32'sd-0.015296912178412303, 32'sd-0.0735577234996024, 32'sd-0.03952319709799749, 32'sd0.043175032391424645, 32'sd-0.002845087033045942, 32'sd0.07421328162617537, 32'sd0.018306151137799986, 32'sd-0.047069172843994846, 32'sd0.018980164035975796, 32'sd1.3297393094793916e-123, 32'sd3.6323711189159675e-117, 32'sd1.6242597959907088e-120, 32'sd6.516698232394128e-124},
        '{32'sd-2.8611371006761545e-122, 32'sd3.0434313307587973e-122, 32'sd1.2299052526795653e-124, 32'sd-7.392815427439167e-122, 32'sd-2.5279326588816705e-121, 32'sd-3.840861536388677e-118, 32'sd-6.949012956085187e-128, 32'sd-1.1629638756599453e-126, 32'sd-4.05786251464148e-115, 32'sd1.984097282045606e-121, 32'sd-1.0011692354527364e-124, 32'sd-9.960836804339497e-120, 32'sd-0.04414720189230485, 32'sd0.021594112336604635, 32'sd0.059750391948036524, 32'sd0.0629904011825651, 32'sd3.0023464220734705e-120, 32'sd2.1038091410314296e-127, 32'sd-3.4646445642085794e-126, 32'sd1.553220565463195e-120, 32'sd3.2492471418581582e-118, 32'sd4.7866317302275894e-123, 32'sd3.4766732014250752e-115, 32'sd2.4889039833596725e-121, 32'sd4.622143653511934e-123, 32'sd-2.5491032324449904e-124, 32'sd-2.7149047569271117e-123, 32'sd-3.2970254160709655e-121, 32'sd-4.849586584503123e-118, 32'sd-7.081982543132779e-128, 32'sd5.4405006698928695e-127, 32'sd9.935956994602461e-123, 32'sd-0.01145556611033266, 32'sd-0.03859271146759927, 32'sd-0.04204168497142301, 32'sd-0.057264279040755046, 32'sd-0.06042780738808257, 32'sd0.013311986617333977, 32'sd0.03809503999927685, 32'sd0.0017183995737811294, 32'sd-0.009580895580339527, 32'sd-0.007126940232023461, 32'sd0.002477119970278169, 32'sd-0.02042910494234007, 32'sd-0.0685721462003698, 32'sd-0.12082281938462718, 32'sd-0.03470537392781379, 32'sd0.039163347090551075, 32'sd0.008498272049379824, 32'sd-0.042380198918576036, 32'sd-0.0612771386398766, 32'sd-0.06344787257388072, 32'sd3.4015995902579317e-125, 32'sd1.4249775757490789e-115, 32'sd-1.0033319127213198e-120, 32'sd-2.6381294361027647e-125, 32'sd1.6680926596804977e-117, 32'sd8.385632954015965e-117, 32'sd-0.008537798983148335, 32'sd-0.04726113451417423, 32'sd-0.08680408540016389, 32'sd0.04990990578005695, 32'sd-0.060479922808370334, 32'sd-0.0030946792257046606, 32'sd-0.038916929422556895, 32'sd0.07095022604821541, 32'sd0.08610810031563741, 32'sd0.08527906149543148, 32'sd0.028976476310859395, 32'sd0.019285570856768592, 32'sd0.062169700414370525, 32'sd-0.07915986313967656, 32'sd-0.07021806066648173, 32'sd-0.03673987051532244, 32'sd0.0146727774422807, 32'sd-0.18375869104580295, 32'sd-0.11292971385522262, 32'sd-0.09672175624016885, 32'sd-0.04898842191763514, 32'sd-0.010103795458344415, 32'sd-0.019180674494780964, 32'sd-0.0017982244279884968, 32'sd4.945529433481508e-118, 32'sd1.0379654834580973e-126, 32'sd5.5966812379707506e-117, 32'sd-7.548275515358404e-115, 32'sd-0.009476208551128266, 32'sd-0.08365337126446812, 32'sd-0.05036265538004424, 32'sd-0.008682607146319587, 32'sd0.021761570013646217, 32'sd-0.0004523264509002509, 32'sd0.0981424357223619, 32'sd0.08508635987693633, 32'sd0.023254856531223066, 32'sd-0.024089672892751962, 32'sd-0.01925255245532282, 32'sd0.0372522890876149, 32'sd-0.00635169298301366, 32'sd0.051919938474070594, 32'sd-0.05002291659691076, 32'sd-0.08427780328565701, 32'sd0.11202291618248617, 32'sd0.06908986696595201, 32'sd-0.020302422268483986, 32'sd-0.07739262007917064, 32'sd0.028722661727099332, 32'sd0.03716482462636446, 32'sd0.04736468543413545, 32'sd-0.005734032469297339, 32'sd0.011336333706956957, 32'sd-1.9935660978625623e-120, 32'sd1.4845261096694666e-126, 32'sd-0.03972528456531155, 32'sd-0.07386313501100131, 32'sd-0.04449589895360379, 32'sd0.04031997035706293, 32'sd-0.04899315241005042, 32'sd-0.0453796047162189, 32'sd-0.04016777380674558, 32'sd-0.05432517026103712, 32'sd0.023136575296205178, 32'sd0.010012104510763398, 32'sd0.04935965148000704, 32'sd0.011371057157255634, 32'sd-0.02861904518660331, 32'sd0.011005555653174782, 32'sd0.08709347808621297, 32'sd0.0405170947031136, 32'sd0.05804844918519934, 32'sd0.10254478232184677, 32'sd0.1027258233411389, 32'sd0.029704996204192567, 32'sd-0.0686384850690992, 32'sd0.03372995796575964, 32'sd0.03134999907145248, 32'sd-0.03448253489374462, 32'sd0.08712530525272542, 32'sd-0.026664092135400205, 32'sd-0.002455225054169595, 32'sd1.865447905381311e-118, 32'sd-0.002807263662909849, 32'sd-0.1012259291449828, 32'sd-0.0012322465653943552, 32'sd0.005296863309487209, 32'sd-0.06559208878520262, 32'sd-0.046455176447006814, 32'sd-0.16835527864455396, 32'sd0.0171672622506663, 32'sd-0.00903268320936245, 32'sd-0.045884190033516147, 32'sd-0.038117596868843306, 32'sd-0.08787865223034531, 32'sd0.009446351638521049, 32'sd-0.057138700813157424, 32'sd0.048153277862094265, 32'sd0.09920902579933819, 32'sd0.0345616034705258, 32'sd0.06545940652058028, 32'sd0.08696491806635814, 32'sd0.13748209623886007, 32'sd0.14109630440704085, 32'sd0.019617836802431864, 32'sd-0.03038582223669906, 32'sd0.002753283786602777, 32'sd0.03180803517910463, 32'sd-0.002259501608904286, 32'sd-0.01959101153896482, 32'sd2.7212066944683274e-121, 32'sd0.025001461648708076, 32'sd-0.11665175455788838, 32'sd0.028772108176475047, 32'sd0.048155165503760325, 32'sd-0.03724076282036314, 32'sd-0.01425619862525458, 32'sd-0.028081940131975264, 32'sd-0.12966774363003009, 32'sd-0.17155538853960794, 32'sd-0.10121321739541282, 32'sd-0.08030653493578241, 32'sd-0.09710404990065906, 32'sd-0.06505105781762398, 32'sd-0.05296142146065995, 32'sd0.13301231761869728, 32'sd0.25628499406249144, 32'sd0.12308730881555434, 32'sd0.18753301437816622, 32'sd0.02931453493301259, 32'sd-0.005710177189673393, 32'sd0.04971904118041704, 32'sd0.023699460431007503, 32'sd-0.016872300526598282, 32'sd-0.1778293210765721, 32'sd0.03377746323804952, 32'sd0.03343645285029184, 32'sd0.0015015043794436172, 32'sd-0.009574051218449474, 32'sd0.02998609767047575, 32'sd-0.0764973401933433, 32'sd0.025538939647648716, 32'sd-0.009895298639467524, 32'sd-0.1325944660889829, 32'sd-0.05053558952274269, 32'sd-0.19601495739209857, 32'sd-0.10859717149501161, 32'sd-0.28093195130491583, 32'sd-0.25169946771818463, 32'sd-0.049789797168373874, 32'sd0.051596421498302174, 32'sd0.0921758468655992, 32'sd0.04810526933179241, 32'sd0.15281393940573587, 32'sd0.07121678400820154, 32'sd0.14827921897055474, 32'sd-0.019368931642700392, 32'sd-0.0011763382963304086, 32'sd-0.18449762429480432, 32'sd0.05786131991250266, 32'sd0.09608701734830552, 32'sd0.06011623490533366, 32'sd-0.14293010963321773, 32'sd-0.09756026750148501, 32'sd0.04114861274558332, 32'sd-0.04087024430773197, 32'sd-0.07461587326151317, 32'sd-0.11416358001008503, 32'sd-0.030721309068502126, 32'sd-0.006470824394439982, 32'sd-0.009677054039625717, 32'sd-0.024049216380848604, 32'sd-0.07839311337695526, 32'sd-0.09994956931227876, 32'sd-0.14783279117745426, 32'sd-0.11119011758228235, 32'sd-0.02655509781203118, 32'sd-0.01839941367071341, 32'sd0.041098368355030446, 32'sd-0.01112051530819789, 32'sd0.03676732876580959, 32'sd-0.05364359811033714, 32'sd-0.011023609024809939, 32'sd-0.07641873860006687, 32'sd0.008178247977006503, 32'sd0.052390559620063094, 32'sd-0.02411450675293469, 32'sd-0.10992148772893437, 32'sd0.05171489056838176, 32'sd0.05877744942602484, 32'sd-0.08192292659030757, 32'sd0.062056038293767754, 32'sd0.06030353952767303, 32'sd0.01982538798597884, 32'sd-0.08528392062650228, 32'sd0.08404607822446593, 32'sd-0.11195061617547611, 32'sd-0.13999642967152598, 32'sd-0.08907046912577649, 32'sd-0.2094527243273724, 32'sd-0.07841701402667091, 32'sd0.05009580635852371, 32'sd-0.014475000264442305, 32'sd0.02846819656372746, 32'sd0.08609668732878951, 32'sd0.12556204441220042, 32'sd0.04206522569490701, 32'sd0.0026589410049394756, 32'sd-0.0638889767431295, 32'sd-0.07047704771772155, 32'sd-0.14567497370454607, 32'sd-0.14499297651123846, 32'sd0.08725800446839646, 32'sd0.085203037066864, 32'sd0.12300078419467023, 32'sd0.08495196298771641, 32'sd-0.03406338266101602, 32'sd0.00987461815124072, 32'sd-0.09133689980972734, 32'sd0.13524366068269741, 32'sd0.0009210158132311525, 32'sd-0.08120739389852792, 32'sd-0.0651973615066343, 32'sd0.048260157461820566, 32'sd-0.004496534657171037, 32'sd0.03288658152408704, 32'sd-0.033602893030023465, 32'sd-0.04756589890841069, 32'sd0.07421866171067483, 32'sd-0.03060449923725536, 32'sd0.018988172008920383, 32'sd0.022386446541047437, 32'sd0.05599021368227011, 32'sd0.11323089670036696, 32'sd0.002898607442310667, 32'sd-0.09564222611868126, 32'sd-0.1644230648357795, 32'sd-0.12353053728848852, 32'sd-0.1352256773538028, 32'sd-0.1231817681685584, 32'sd0.086378132983542, 32'sd0.04523559259029183, 32'sd0.065654736323416, 32'sd-0.009332922084254403, 32'sd0.09909297273806182, 32'sd0.1093824740759106, 32'sd0.046998940866352854, 32'sd-0.01701126639719822, 32'sd-0.024969120131956776, 32'sd0.045846149828635295, 32'sd-0.08189437214502475, 32'sd-0.07899426411252361, 32'sd0.004220019587031368, 32'sd-0.06263038848845728, 32'sd-0.024478619682157136, 32'sd0.07592083386953857, 32'sd0.15490920837840064, 32'sd0.1986526677865164, 32'sd-0.09243874306246859, 32'sd-0.055874123476321924, 32'sd-0.04079037010262456, 32'sd0.031996217892693496, 32'sd-0.18129173741261773, 32'sd-0.2685649180066076, 32'sd-0.14385728080327653, 32'sd-0.06376937093859528, 32'sd-0.04103892219608767, 32'sd-0.12300212684345423, 32'sd0.08623612856167424, 32'sd0.14781744068080546, 32'sd-0.007164375887010331, 32'sd0.05147616267700147, 32'sd0.049718644040910406, 32'sd0.04665644201496906, 32'sd-0.008306486881087045, 32'sd0.007616235454100684, 32'sd0.0016038784268821442, 32'sd-0.09645439578490544, 32'sd-0.08547658310243315, 32'sd-0.1215526446830263, 32'sd-0.0745452339567181, 32'sd0.07994854894059812, 32'sd0.13643801582837223, 32'sd0.12090779187611964, 32'sd0.17904227136654563, 32'sd0.021645643907529388, 32'sd-0.03756616025715129, 32'sd-0.028530742562622113, 32'sd-0.10327650684645025, 32'sd-0.20181438841285687, 32'sd-0.21946367821913604, 32'sd-0.17058546268790337, 32'sd0.10925121349201936, 32'sd-0.05542115934509718, 32'sd-0.04579596715153934, 32'sd0.02359737805717021, 32'sd-0.035824171364091065, 32'sd-0.02349241925845823, 32'sd-0.07337323169585175, 32'sd0.10872576153470281, 32'sd-0.006562902445866726, 32'sd0.12985610104200307, 32'sd0.0902535147576659, 32'sd-0.027346681083104382, 32'sd-0.11884066395871627, 32'sd0.010842601754007876, 32'sd-0.03468379398957485, 32'sd-0.11728612824369002, 32'sd0.002976201992979457, 32'sd0.17761075568218046, 32'sd0.05392098789112667, 32'sd-0.10234122945266468, 32'sd-0.005712798238360328, 32'sd-0.09128305360660939, 32'sd-0.06079193308723263, 32'sd0.02779905386547852, 32'sd-0.13233593529148938, 32'sd-0.20085131614357057, 32'sd-0.24864765426651675, 32'sd-0.07052407841081813, 32'sd0.12730057463893174, 32'sd-0.014572316501697567, 32'sd-0.05571525903694616, 32'sd-0.03810000937445467, 32'sd-0.06913200172277335, 32'sd-0.08715111785758495, 32'sd-0.03461155961181537, 32'sd-0.016826624225708738, 32'sd0.017453929070885565, 32'sd0.0077788729339047305, 32'sd-0.06090580555887438, 32'sd-0.13442279144033628, 32'sd-0.13234686500109968, 32'sd-0.08157385071909595, 32'sd-0.051320994779455543, 32'sd-0.13487779222804985, 32'sd-0.02624925972658718, 32'sd0.05797798737426517, 32'sd-0.17123879057722705, 32'sd-0.1308148742288486, 32'sd-0.15616862421074895, 32'sd-0.27242122093960236, 32'sd-0.25463739160266335, 32'sd-0.16789275634009762, 32'sd-0.17673884105818913, 32'sd-0.10618115484174633, 32'sd-0.03758281659746234, 32'sd0.022110603032011674, 32'sd0.170836059104029, 32'sd0.11100629104785607, 32'sd-0.003633525882245753, 32'sd-0.1545231399848701, 32'sd-0.05629000324478685, 32'sd-0.058240235921941975, 32'sd-0.2285111068025451, 32'sd-0.11180828784449703, 32'sd-0.08136794783409448, 32'sd-0.09776831439398703, 32'sd-0.09201170717356752, 32'sd0.015474384245990765, 32'sd0.06888833047129547, 32'sd-0.06450065091517058, 32'sd0.010002995130121489, 32'sd-0.01339769986914791, 32'sd0.017364407023288654, 32'sd-0.08033987173892479, 32'sd-0.13298309784242618, 32'sd-0.20290660732546653, 32'sd-0.18420719436950017, 32'sd-0.11182373577494095, 32'sd-0.05475947444564747, 32'sd-0.12443674078935549, 32'sd-0.04239868437645847, 32'sd-0.037226205605895984, 32'sd-0.05084076738612339, 32'sd0.1135625608991031, 32'sd0.1983955491452239, 32'sd0.0059879984971254, 32'sd-0.052420132695150425, 32'sd-0.09739101802237665, 32'sd-0.025060088831438815, 32'sd-0.06606031035490341, 32'sd-0.14338458026063586, 32'sd-0.20979323761159038, 32'sd-0.03066860491879608, 32'sd-0.06950685660362266, 32'sd-0.13320279757237383, 32'sd-0.06942264210242963, 32'sd-0.022668099745524063, 32'sd0.040703580900058704, 32'sd0.025297990870108072, 32'sd-0.06238811880632854, 32'sd-0.06886307831879354, 32'sd0.020796483820096377, 32'sd-0.07603159435678734, 32'sd-0.15720876078732018, 32'sd-0.10749087528317001, 32'sd-0.011323194198520714, 32'sd0.03403964891795797, 32'sd0.06715958393869405, 32'sd0.07536298658339687, 32'sd0.08817498321312352, 32'sd0.03337357568222741, 32'sd0.04960748745480031, 32'sd0.15600272173555893, 32'sd-0.07380593559234494, 32'sd-0.08671873397291233, 32'sd-0.12411747404020802, 32'sd-0.18698983823358017, 32'sd-0.1306639626192738, 32'sd-0.0707433875351563, 32'sd-0.03038911011321682, 32'sd-0.04691706540983746, 32'sd0.030643732722041662, 32'sd-0.013768263088252039, 32'sd-0.06146389885139095, 32'sd-0.10822296629051062, 32'sd0.009684072766104897, 32'sd-4.125072304130201e-125, 32'sd-0.05170594409246672, 32'sd-0.09752633101920145, 32'sd-0.008219060531137572, 32'sd-0.014358229035330914, 32'sd-0.022556783315606795, 32'sd-0.026139297803944264, 32'sd0.059691045092399156, 32'sd0.05721834445696912, 32'sd0.09995823741480576, 32'sd0.12219887581928027, 32'sd0.10675611054022559, 32'sd0.10956689240818107, 32'sd-0.013548037704033155, 32'sd-0.043429657327145814, 32'sd0.0894004276967792, 32'sd-0.05844205011514437, 32'sd-0.04626877893043029, 32'sd-0.14757104946874963, 32'sd-0.08186659157055808, 32'sd-0.11273216872623074, 32'sd-0.1543376078209839, 32'sd-0.03210992946076944, 32'sd-0.09342243932427512, 32'sd-0.08723034735351408, 32'sd0.04678095860663736, 32'sd-0.027213507410786795, 32'sd-0.012336525186111764, 32'sd-0.034903992738666956, 32'sd-0.0753232199196648, 32'sd-0.0486856764041034, 32'sd-0.004041126792640355, 32'sd0.04183301217199293, 32'sd0.09271676705790766, 32'sd0.11808107121603008, 32'sd0.17252309690786294, 32'sd0.03799655595445422, 32'sd0.00393548574739194, 32'sd0.03680034868119495, 32'sd-0.05779327424957739, 32'sd-0.11198331632165853, 32'sd-0.11404756573256455, 32'sd0.06234798752677011, 32'sd0.05497282447636204, 32'sd0.09980178741095032, 32'sd-0.010101655863123607, 32'sd-0.062154930367784425, 32'sd-0.15167768978297916, 32'sd-0.04496490922741608, 32'sd-0.05941434571878173, 32'sd-0.09106477253874891, 32'sd-0.15368694070587158, 32'sd-0.04841140249050863, 32'sd-0.006985398105619949, 32'sd0.052508635776184254, 32'sd0.047411350929049786, 32'sd-0.04412406952067062, 32'sd-0.07888581338554687, 32'sd-0.14687436103021226, 32'sd-0.12150575848571524, 32'sd0.04845122608351704, 32'sd0.0036112519810356293, 32'sd0.05093015617130664, 32'sd0.0586939995355658, 32'sd0.013740672986891184, 32'sd0.022781519061997456, 32'sd-0.11118729037698488, 32'sd-0.14576047363588876, 32'sd-0.06649820705909093, 32'sd-0.0800947823256921, 32'sd0.037636227484191466, 32'sd0.10051709483695534, 32'sd0.08082324820709634, 32'sd0.028298412481979472, 32'sd0.02589875996889322, 32'sd-0.06709458198494514, 32'sd0.07158172789881767, 32'sd0.053497016626328206, 32'sd-0.07149781037713154, 32'sd-0.033138114180644995, 32'sd0.07914661968898068, 32'sd-0.06844409703067263, 32'sd-0.00948792905871675, 32'sd-0.08276877953991199, 32'sd-5.804805416987397e-115, 32'sd-0.11425019569331646, 32'sd-0.10083061767759632, 32'sd-0.012400202184969402, 32'sd0.007025818879032601, 32'sd0.09865210482946593, 32'sd0.012799226907413596, 32'sd0.20132833396860428, 32'sd0.2022865030446442, 32'sd0.15599038782359112, 32'sd-0.04120894358781592, 32'sd-0.14298970881387446, 32'sd0.0020286817249125177, 32'sd-0.09116649586776618, 32'sd0.02886289102649753, 32'sd0.09979425299121153, 32'sd0.06980066596029112, 32'sd0.19970160220875685, 32'sd0.16596358556190327, 32'sd0.024219339438953706, 32'sd0.11716408507224972, 32'sd0.05315331721285336, 32'sd-0.034225555668901175, 32'sd0.004168428121211624, 32'sd-0.01961734919873627, 32'sd0.03608429124357336, 32'sd0.009674714299466688, 32'sd-0.039237442240566495, 32'sd0.0007515129982685736, 32'sd-0.07658083973768798, 32'sd-0.1025001871471365, 32'sd-0.038642053625470685, 32'sd0.08452057629819144, 32'sd0.08735457005776302, 32'sd0.04389941309047736, 32'sd0.13951037902581678, 32'sd0.15339586429868493, 32'sd-0.0017666185265695327, 32'sd-0.04300921781903868, 32'sd-0.00766861944411031, 32'sd-0.07368228889400194, 32'sd0.11030986398903068, 32'sd0.10351150036227787, 32'sd0.11996679190455035, 32'sd0.050531172977151095, 32'sd0.13225228641047004, 32'sd0.1608129870755047, 32'sd0.20941736677291276, 32'sd0.0016625694424854164, 32'sd0.04688705679683736, 32'sd0.010284215697077742, 32'sd0.018243405634367278, 32'sd-0.0075184422965009325, 32'sd0.013700810657541834, 32'sd0.0009187910029351409, 32'sd0.015693756240595075, 32'sd-0.001566908444064506, 32'sd0.0019564101933023568, 32'sd-0.017820892094398345, 32'sd0.0978878351706058, 32'sd0.11910921174020751, 32'sd0.010240267345609155, 32'sd0.12870533715847973, 32'sd0.0730950517905462, 32'sd0.008786767572648912, 32'sd-0.0010319197215138104, 32'sd-0.008674558725776335, 32'sd0.09097417949736285, 32'sd0.15141348883914638, 32'sd0.10653416191348446, 32'sd0.13133054267563052, 32'sd0.0061303933345811116, 32'sd0.03441957075627503, 32'sd0.060970338315446126, 32'sd0.07176940736557658, 32'sd0.0994109755309026, 32'sd0.004884606563818434, 32'sd0.044229879816466984, 32'sd0.05485395907100812, 32'sd0.03622936469785294, 32'sd0.01407212734220562, 32'sd0.0365415503169473, 32'sd-0.02690809935458561, 32'sd0.014393826720091592, 32'sd-9.441592369117129e-123, 32'sd-0.05407597179303549, 32'sd0.019989184132425078, 32'sd0.009873622416947905, 32'sd-0.01179258024909013, 32'sd0.057010630107329145, 32'sd-0.0007529236831076045, 32'sd-0.02988964524302604, 32'sd0.021538469711858174, 32'sd-0.02885085260088653, 32'sd0.1338796448520897, 32'sd0.17297331162966212, 32'sd0.09043505847101639, 32'sd0.08641766494221907, 32'sd0.005629926592420944, 32'sd-0.053249124264673146, 32'sd0.12377894549637068, 32'sd-0.02190469639780431, 32'sd0.0033889162185493826, 32'sd-0.019937564042401792, 32'sd-0.014135818949114629, 32'sd0.13781262991083762, 32'sd0.08129890276031733, 32'sd0.08001829726356753, 32'sd-0.016695029819580102, 32'sd-0.09362417702710753, 32'sd-0.09772991521377998, 32'sd4.876356805531312e-124, 32'sd2.975760908485609e-129, 32'sd1.0412785307572843e-125, 32'sd-0.024648590628182924, 32'sd0.015471474406873022, 32'sd0.055376854368638165, 32'sd-0.10024036903789056, 32'sd-0.05131522199234359, 32'sd-0.07036716970717137, 32'sd-0.042217590122549095, 32'sd-0.09186731579287419, 32'sd-0.016434729911529302, 32'sd0.07672012516448397, 32'sd-0.022917245661237047, 32'sd-0.03893439113731776, 32'sd-0.1486479808991776, 32'sd-0.0014139416264565758, 32'sd-0.08349094438957103, 32'sd0.02922813114149508, 32'sd0.06614755497956454, 32'sd-0.03915473109225775, 32'sd-0.023140014219134277, 32'sd0.04082122801990335, 32'sd-0.08276653333639505, 32'sd0.023750032865878914, 32'sd-0.01098591367860177, 32'sd-0.03675868752926452, 32'sd-0.004486796911537366, 32'sd-6.0218871452833e-117, 32'sd2.4169808666950206e-125, 32'sd-2.4009460764350994e-121, 32'sd-0.05994581217386131, 32'sd0.01682006492731889, 32'sd-0.12566020776307985, 32'sd-0.07133194969385478, 32'sd-0.029767542701452532, 32'sd-0.12184760594293202, 32'sd0.013931218414540265, 32'sd-0.06711949842451728, 32'sd-0.09444239190379816, 32'sd-0.04220558126114952, 32'sd-0.13870722866170762, 32'sd0.023226772289036374, 32'sd0.06032637612860888, 32'sd-0.051618471181535695, 32'sd-0.058902705330919826, 32'sd-0.08281561858568004, 32'sd-0.10209276929072926, 32'sd-0.1430598995969712, 32'sd0.0036681746420293977, 32'sd-0.03118943076326644, 32'sd-0.04161154981198935, 32'sd-0.10083567944252968, 32'sd-0.092727877469663, 32'sd0.018007504815243002, 32'sd-0.015559049496622696, 32'sd-2.837402810081404e-118, 32'sd2.8798504276300483e-120, 32'sd-2.5618982422508916e-122, 32'sd-5.830698166226577e-129, 32'sd-0.012524836467907417, 32'sd-0.024171031966443376, 32'sd-0.05995974061589276, 32'sd-0.035407772405424864, 32'sd-0.07459788158331566, 32'sd0.058330540217547716, 32'sd0.05917655494723809, 32'sd2.5812253554346735e-05, 32'sd0.01641968960212992, 32'sd-0.037631442316916015, 32'sd-0.004762692881383438, 32'sd-0.08672023828482746, 32'sd-0.12028605124607225, 32'sd-0.00864458705814975, 32'sd-0.12981414433498104, 32'sd-0.13161735744228023, 32'sd-0.10725143468405116, 32'sd-0.13269635228499632, 32'sd-0.08126018186246717, 32'sd-0.07307340142152771, 32'sd-0.10379657536269214, 32'sd-0.07165108229724435, 32'sd-0.015941474867460084, 32'sd2.0090905063457977e-117, 32'sd3.4570786125238072e-118, 32'sd2.3040672931503832e-117, 32'sd-2.5810384477492876e-121, 32'sd2.6614830540461016e-120, 32'sd7.330112227687378e-115, 32'sd0.0033034759944422384, 32'sd-0.025176578244591137, 32'sd-0.08438412494597416, 32'sd-0.03268386101345682, 32'sd-0.09702352321189224, 32'sd0.029836443177680173, 32'sd0.029342471283708326, 32'sd-0.046137752075804665, 32'sd-0.06815032180481372, 32'sd0.04080222647103935, 32'sd-0.02609580529170047, 32'sd0.03396992100384661, 32'sd0.03889872270065577, 32'sd-0.0849222371754567, 32'sd-0.03798197901589763, 32'sd-0.07821027916422749, 32'sd-0.08096540674959189, 32'sd-0.10812640651463883, 32'sd-0.013671792912303887, 32'sd-0.003268243716115142, 32'sd-1.3945500932816094e-125, 32'sd-5.530114375097967e-120, 32'sd8.868088647511567e-124, 32'sd2.8495708698821627e-125},
        '{32'sd3.6282195155808275e-114, 32'sd-1.3030342560760605e-125, 32'sd2.984278744578858e-123, 32'sd2.4353411946195372e-123, 32'sd9.437088032744328e-124, 32'sd-1.8163481147392741e-124, 32'sd-1.5219969620281675e-120, 32'sd9.965454773100257e-118, 32'sd-4.545358330099518e-118, 32'sd-5.8643585384889574e-120, 32'sd1.6807298858953663e-123, 32'sd6.955862314111214e-127, 32'sd-0.02502498429935392, 32'sd-0.038435075040335, 32'sd0.05211737828483769, 32'sd0.03547513584905297, 32'sd1.2726138897691781e-118, 32'sd-1.0527527698883845e-119, 32'sd4.096288267951394e-115, 32'sd9.889161986709614e-122, 32'sd-6.787368763072985e-126, 32'sd-7.622191924326416e-127, 32'sd3.6547808431631983e-119, 32'sd1.0063129678872209e-124, 32'sd8.061526937311883e-128, 32'sd-2.6023018474490355e-124, 32'sd-2.468236103870511e-120, 32'sd5.6364509281590336e-123, 32'sd2.9209302754640837e-118, 32'sd-2.1159864897233335e-127, 32'sd-4.6734849664843324e-124, 32'sd-1.5173243666435326e-124, 32'sd0.1156607210070177, 32'sd-0.059800254564522766, 32'sd0.06450689522105803, 32'sd0.02043788754805735, 32'sd0.07887599869056523, 32'sd0.05167028291840594, 32'sd0.008878747864080777, 32'sd0.06264739714160271, 32'sd0.0691953770707428, 32'sd0.06938824750025425, 32'sd0.026642353570935706, 32'sd0.15264003480975832, 32'sd0.07606820292159383, 32'sd0.07867444028045158, 32'sd0.09955685416923754, 32'sd0.016430325228905193, 32'sd0.03323808976869396, 32'sd0.07289609818821159, 32'sd0.015837311278107256, 32'sd0.030827301539792754, 32'sd8.548077109618619e-122, 32'sd1.9705618874288014e-126, 32'sd5.7573801016592343e-126, 32'sd-9.154539690005347e-120, 32'sd3.5203423141596745e-119, 32'sd-2.687464116156036e-124, 32'sd0.07630860371023662, 32'sd-0.001326919842896503, 32'sd0.1003341523922412, 32'sd-0.023300968534420378, 32'sd0.008562879537609936, 32'sd-0.03853512238441238, 32'sd0.08528320203025551, 32'sd0.042691783233487185, 32'sd-0.06862534090955608, 32'sd0.07499409682154594, 32'sd-0.12458713535499416, 32'sd0.05312943247332521, 32'sd-0.0698566874794207, 32'sd0.05564612227206094, 32'sd0.14324516534418769, 32'sd0.12624584733382688, 32'sd0.13982342136258785, 32'sd0.029595777134721512, 32'sd0.03791816874098813, 32'sd0.10254238241464624, 32'sd0.024774188091993454, 32'sd0.07024972012303757, 32'sd0.052712847578524694, 32'sd0.05370220286433857, 32'sd-1.4211432077191799e-118, 32'sd-5.815960091289632e-127, 32'sd2.9848711989375087e-116, 32'sd-1.2552009580919503e-127, 32'sd0.06667540984543188, 32'sd0.04607560967940635, 32'sd-0.031513023392119366, 32'sd0.06968823538645649, 32'sd0.0456583801580894, 32'sd0.09429455597232222, 32'sd0.06506485913545136, 32'sd0.032145108256980304, 32'sd-0.0027966081769413126, 32'sd-0.0856199113669314, 32'sd0.0011133524320510112, 32'sd0.023007063406634706, 32'sd0.026107255613506405, 32'sd-0.09389235652447415, 32'sd-0.01796797196094174, 32'sd0.043066855095951415, 32'sd0.060532304782069106, 32'sd-0.02810757019059411, 32'sd0.0768016261321798, 32'sd0.060663914868586716, 32'sd0.03178222328438291, 32'sd0.02677359532940206, 32'sd-0.036853760722150755, 32'sd0.03967582722978649, 32'sd0.11254705337926679, 32'sd-5.761069453456586e-119, 32'sd-3.693331740867155e-119, 32'sd0.024550026048677183, 32'sd0.01463415588249246, 32'sd-0.03633626382512909, 32'sd-0.005290164619785898, 32'sd0.16434681997761288, 32'sd0.042168578930757865, 32'sd0.07678794364209439, 32'sd-0.011938170633676089, 32'sd-0.062041577338329094, 32'sd-0.03575958129107172, 32'sd-0.08402721823760845, 32'sd0.0953064982807619, 32'sd0.12465072761738619, 32'sd0.08562311300779689, 32'sd0.043420868449026324, 32'sd-0.017479668042016214, 32'sd0.05314473769430411, 32'sd-0.04028532863859186, 32'sd0.00998160711209844, 32'sd0.04469702008113967, 32'sd0.02128322359731564, 32'sd0.040565512516458874, 32'sd-0.007163377302151817, 32'sd0.05062311872805349, 32'sd0.0400218582259168, 32'sd-0.05757833920144103, 32'sd0.011596885168821383, 32'sd-1.2154778989822904e-117, 32'sd0.05205205796744961, 32'sd0.0879289302650175, 32'sd0.07076050326215669, 32'sd0.08494586754745365, 32'sd0.054207961889528096, 32'sd0.003702821453714677, 32'sd0.03890571336799595, 32'sd0.06987278903375381, 32'sd0.01632347910341952, 32'sd-0.08969846495867695, 32'sd-0.009551321737943761, 32'sd0.03335548776049033, 32'sd0.032330269258044275, 32'sd-0.04399328964994629, 32'sd-0.05463250039193836, 32'sd0.058053517652462264, 32'sd0.06294152575119873, 32'sd0.06966779551116757, 32'sd0.13305078247212263, 32'sd0.061282002160926566, 32'sd-0.01196507805893282, 32'sd0.034953783302438486, 32'sd-0.012396722903241992, 32'sd0.012528755958415384, 32'sd0.03790547344894873, 32'sd0.05675511505225762, 32'sd0.05831181795605807, 32'sd-3.0937868125678666e-122, 32'sd-0.014470276837503342, 32'sd-0.011119388728195857, 32'sd0.05539661667715316, 32'sd-0.02145288794873877, 32'sd-0.05319402398808991, 32'sd-0.007617851456759637, 32'sd0.018364859227709064, 32'sd-0.03690892236141373, 32'sd0.005203137644380249, 32'sd-0.04712019736148725, 32'sd0.08385334222384996, 32'sd0.06362416245434933, 32'sd0.008623987193954222, 32'sd-0.1464922666328192, 32'sd-0.031163989929323933, 32'sd-0.07187384855051457, 32'sd0.1563319679742065, 32'sd0.02790854535906788, 32'sd0.03467975661404752, 32'sd0.020855254130965607, 32'sd0.0350723480714472, 32'sd0.020238974094386436, 32'sd0.011797861301800867, 32'sd-0.0735732826384627, 32'sd0.12603209963035963, 32'sd0.07822924313627427, 32'sd0.01701895070691586, 32'sd0.11364680160969551, 32'sd-0.001055052417303427, 32'sd0.009734577824560728, 32'sd-0.050089493861309814, 32'sd-0.03037489851178777, 32'sd0.03916165963956618, 32'sd0.0027205298696654544, 32'sd-0.027594190410789244, 32'sd0.036067873026724616, 32'sd0.027341116717657894, 32'sd0.0705119602957009, 32'sd0.07835344504306174, 32'sd0.09718938053544976, 32'sd-0.08098602767931706, 32'sd-0.012251615492995013, 32'sd0.02392681618387769, 32'sd-0.10772458076697644, 32'sd-0.005822961793006944, 32'sd-0.14456409173514756, 32'sd-0.17273152544079753, 32'sd-0.012623183292623161, 32'sd0.007281352717217577, 32'sd0.04210517991798484, 32'sd-0.0018388243406382632, 32'sd0.08828437297986826, 32'sd0.00590818170318206, 32'sd-0.015701027707310952, 32'sd0.005809501542000224, 32'sd0.07744111904306476, 32'sd0.061208135134545816, 32'sd0.03140968024049573, 32'sd-0.057512664920927305, 32'sd0.04117485252636155, 32'sd-0.06597816435893958, 32'sd-0.09670011302008294, 32'sd0.000416435162904306, 32'sd0.022406314083483897, 32'sd-0.07557220423766296, 32'sd0.04006390069592561, 32'sd0.07870605146327458, 32'sd-0.02155639665999355, 32'sd-0.047157851652863264, 32'sd-0.11450099804707627, 32'sd-0.01955444953019277, 32'sd0.02737851184681912, 32'sd-0.07452751150652497, 32'sd-0.10257267462104293, 32'sd-0.2090236090364937, 32'sd-0.09628738197065144, 32'sd-0.07018120390776807, 32'sd-0.05116203105654296, 32'sd0.0950951653595234, 32'sd-0.061858811636911676, 32'sd-0.1122589465109182, 32'sd0.017628433056595665, 32'sd0.004323763889039877, 32'sd0.05798405537066887, 32'sd-0.01386085563702466, 32'sd0.013229331880803134, 32'sd-0.06016042203218695, 32'sd0.09624879662702696, 32'sd0.048815452975058224, 32'sd-0.014497940304514874, 32'sd0.03894680743130699, 32'sd0.1252919465539054, 32'sd-0.004997145824125132, 32'sd0.10546553890675703, 32'sd0.024248593920686245, 32'sd-0.08803354656690418, 32'sd-0.0754583661429914, 32'sd0.024546213720289152, 32'sd-0.06930880572197899, 32'sd-0.1696343235155373, 32'sd-0.05043346214920944, 32'sd-0.14348637774631776, 32'sd-0.15742163036969983, 32'sd-0.15344442337475186, 32'sd-0.12716953314109458, 32'sd0.00862289702931176, 32'sd0.030586907098854595, 32'sd-0.137304460372331, 32'sd0.00797329665822754, 32'sd0.10251442806742056, 32'sd-0.01596840526776232, 32'sd0.030186213247058922, 32'sd-0.0655239138490555, 32'sd0.008103291933967837, 32'sd-0.048215992985521906, 32'sd0.021786019430917403, 32'sd0.08946747937897936, 32'sd0.061923378150235873, 32'sd0.013267994105602011, 32'sd-0.019394397847502944, 32'sd0.005658483853468289, 32'sd-0.01548121960361249, 32'sd-0.02002047781412945, 32'sd-0.07181920937552148, 32'sd-0.143349348049387, 32'sd-0.080061677987652, 32'sd-0.1988663877878324, 32'sd-0.16613338876632222, 32'sd-0.23121690257215538, 32'sd-0.2064456597666313, 32'sd-0.26247402966400774, 32'sd-0.06366027778257012, 32'sd-0.09438526849797989, 32'sd-0.03998687567939442, 32'sd-0.09373690378945784, 32'sd-0.07209159273191675, 32'sd0.02494180116102909, 32'sd0.044036939136866744, 32'sd0.01485388455868846, 32'sd-0.05695476822699382, 32'sd0.04350614168699256, 32'sd-0.08868515567116796, 32'sd0.034122068209141036, 32'sd-0.05551103707267304, 32'sd-0.06582403792392319, 32'sd-0.10801857418142718, 32'sd-0.0512784574957826, 32'sd-0.02916462858351735, 32'sd-0.07352853557889406, 32'sd0.012794069800891362, 32'sd-0.14721970371693402, 32'sd-0.08931479432278137, 32'sd-0.11564413476548263, 32'sd-0.0506347159641238, 32'sd-0.19126346080190734, 32'sd-0.1605496737689509, 32'sd-0.10587813109061776, 32'sd-0.21329437097526824, 32'sd-0.1063563606343363, 32'sd-0.08634891975458595, 32'sd-0.11573745020675372, 32'sd0.01262986564475823, 32'sd-0.014842582527508374, 32'sd-0.0249799418442676, 32'sd0.009978773034537517, 32'sd0.03292271554144304, 32'sd-0.007228857423272188, 32'sd0.07120999316472078, 32'sd0.06055264021152542, 32'sd0.06958424851506534, 32'sd0.05749052282144603, 32'sd-0.012652268344494733, 32'sd0.02357810474671818, 32'sd-0.10572870743122234, 32'sd-0.0982623553222054, 32'sd0.038322021057803565, 32'sd-0.08021841149855531, 32'sd-0.09382698490476576, 32'sd-0.00037005694610635744, 32'sd-0.045833413512562246, 32'sd-0.12489686387263636, 32'sd-0.015612899712643132, 32'sd-0.08601303691013983, 32'sd-0.19263848128185207, 32'sd-0.12131826274461464, 32'sd0.004004776913331218, 32'sd-0.10101497016390815, 32'sd-0.1467757628402087, 32'sd-0.1899536759157815, 32'sd-0.12329435355268756, 32'sd0.0563237119315059, 32'sd0.026673308178391465, 32'sd-0.12960417103823893, 32'sd0.04198244308702771, 32'sd0.01780015628531619, 32'sd0.09537693138055789, 32'sd0.060900248477127626, 32'sd0.050638136383498455, 32'sd-0.06620548142093169, 32'sd-0.03553274399988392, 32'sd-0.00035066225464598915, 32'sd0.0632281043911391, 32'sd0.019668102973374454, 32'sd-0.12150268026266949, 32'sd-0.10264312770534538, 32'sd0.01004645505519857, 32'sd0.08542957861028862, 32'sd0.0006243914190410605, 32'sd0.004508713629915118, 32'sd-0.01696896721708873, 32'sd-0.07109135257776056, 32'sd-0.039333805951363286, 32'sd0.0026405075869762565, 32'sd0.0531824677649328, 32'sd-0.08023274867213924, 32'sd-0.1515888053714262, 32'sd-0.037874635707728435, 32'sd-0.0833882097660322, 32'sd0.03118230460997494, 32'sd0.10487534650918248, 32'sd0.07546069603750626, 32'sd0.081992654560513, 32'sd0.09775866351242031, 32'sd0.035151665872346326, 32'sd0.03562687282056573, 32'sd0.048230527371108736, 32'sd-0.0658230872270041, 32'sd0.017521907324922936, 32'sd0.04827794973407108, 32'sd-0.01572926418387795, 32'sd-0.07386997745390878, 32'sd0.016250380177230028, 32'sd-0.024419950637747104, 32'sd0.10406293230340168, 32'sd0.07541446412265465, 32'sd0.06932320517838338, 32'sd0.06647164912603634, 32'sd0.05139461560067343, 32'sd0.061004090254655106, 32'sd0.0885412917747229, 32'sd-0.060446981599241494, 32'sd0.046895559003625, 32'sd-0.10605559906027127, 32'sd-0.005019992467303274, 32'sd0.05531981602674288, 32'sd0.008241397104787978, 32'sd0.041944185251267106, 32'sd-0.005208903393277771, 32'sd-0.02891426014869028, 32'sd0.13238078595128935, 32'sd0.013938433730399878, 32'sd0.018088106474683292, 32'sd0.07330641549086479, 32'sd-0.07044274884065589, 32'sd0.043850538938653046, 32'sd-0.0336529541531002, 32'sd0.09686239030341683, 32'sd0.10768700795912328, 32'sd-0.03184371529651118, 32'sd0.032303126399104425, 32'sd-0.10507308781379686, 32'sd0.006322606053978278, 32'sd-0.023617268607567, 32'sd0.010040210519530695, 32'sd0.0900675445421232, 32'sd0.05943455262610136, 32'sd0.15559007310023615, 32'sd0.11723538548044896, 32'sd0.08078082779400542, 32'sd0.12022582299048439, 32'sd-0.03144340329025098, 32'sd0.04082368634935781, 32'sd0.03831257345178647, 32'sd-0.0856839520583942, 32'sd-0.007065774548375259, 32'sd0.0176280489949565, 32'sd0.05706457681304967, 32'sd0.03198232508476349, 32'sd-0.03204030354586118, 32'sd0.08987132448741153, 32'sd0.011935607735467046, 32'sd-0.022294121588870074, 32'sd-0.045530397605375354, 32'sd0.029047818563091462, 32'sd0.031452514589052474, 32'sd0.015564564637698283, 32'sd-0.009427450319638752, 32'sd-0.08411321590809126, 32'sd-0.09623699093759155, 32'sd-0.04085459365276043, 32'sd-0.018456538763483802, 32'sd-0.09314099471472548, 32'sd-0.014419721590934723, 32'sd0.17940040121196474, 32'sd0.13477137272284978, 32'sd0.11912968078884145, 32'sd0.019971724795459046, 32'sd0.015578160650058225, 32'sd-0.09917451421464102, 32'sd0.12700623916167209, 32'sd0.02897796416154919, 32'sd-0.03995755306260325, 32'sd-0.026111444379033028, 32'sd0.022621595171308725, 32'sd0.01605622198883062, 32'sd-0.037791386605624054, 32'sd0.03705410585815283, 32'sd-1.5460874996707152e-125, 32'sd0.027399518496306976, 32'sd0.013020943394141024, 32'sd0.10506680168452608, 32'sd0.025730263768972163, 32'sd-0.04635260612708881, 32'sd0.12296517384171092, 32'sd0.07472598916450313, 32'sd0.07025107734990658, 32'sd-0.14224903229598063, 32'sd-0.09102923104924637, 32'sd-0.020154546162860377, 32'sd-0.02360530332311356, 32'sd0.08549087138611372, 32'sd0.18466970971854352, 32'sd0.047959313217138935, 32'sd0.05830014220018921, 32'sd0.08471489522871613, 32'sd-0.05153454025713007, 32'sd0.0228035623138136, 32'sd0.05271856243253393, 32'sd-0.003567415489812124, 32'sd-0.04761684949155697, 32'sd0.07183867353080435, 32'sd0.03121544703802063, 32'sd-0.05003210010137572, 32'sd-0.12707603923853336, 32'sd-0.05856826488684208, 32'sd0.08508159143662247, 32'sd0.025071352863595395, 32'sd-0.009160518662513049, 32'sd0.008833267309582572, 32'sd0.050108488760229206, 32'sd-0.04321019563720045, 32'sd-0.003990032474798319, 32'sd-0.018334381735600896, 32'sd0.045989492802729584, 32'sd-0.044708682002358675, 32'sd-0.040066773223399424, 32'sd-0.04802549789201205, 32'sd0.02209272469011021, 32'sd0.034915136857443865, 32'sd0.06830472641610985, 32'sd0.07700392856904159, 32'sd0.13857140157980788, 32'sd0.1339197112861782, 32'sd0.056148566776655244, 32'sd0.03894882003965607, 32'sd-0.03433620599706988, 32'sd0.015294431475410241, 32'sd-0.06000637948614736, 32'sd0.04161313002803415, 32'sd0.013986974079390369, 32'sd0.14191487182176374, 32'sd0.025485018372958225, 32'sd-0.02332032740406527, 32'sd0.03229053885573909, 32'sd0.022914289934203375, 32'sd0.07667626153822268, 32'sd-0.06020172764590624, 32'sd0.059478793334805706, 32'sd-0.06319288924917708, 32'sd-0.02354996980446834, 32'sd0.056689239657732544, 32'sd0.1283329315132835, 32'sd-0.056419627841086235, 32'sd-0.02658408519380116, 32'sd-0.029418882027117708, 32'sd0.06825271547818255, 32'sd0.06155221964590857, 32'sd0.0917900460390681, 32'sd0.05865720077616888, 32'sd0.1441258530175501, 32'sd0.10941403726619907, 32'sd0.028682694239917494, 32'sd0.045690750540755005, 32'sd0.041972796923167556, 32'sd-0.03532942666681736, 32'sd-0.0021553062675502286, 32'sd0.09827445469307819, 32'sd-0.11430018740592865, 32'sd0.08865370051804258, 32'sd0.0695544116343968, 32'sd0.025049848827110872, 32'sd2.0329931496939776e-121, 32'sd0.025046698662129448, 32'sd0.07324143509494102, 32'sd0.015742415230509958, 32'sd-0.03451989154343586, 32'sd0.05071704632898456, 32'sd-0.02453986524551453, 32'sd0.08024000696392877, 32'sd0.07361489234253822, 32'sd0.04754494627639794, 32'sd0.04912491999004355, 32'sd0.12890863694922358, 32'sd0.06222811875088142, 32'sd0.04815394583392959, 32'sd0.10457160398908143, 32'sd0.042620044301152425, 32'sd0.05755059584392797, 32'sd-0.06408980287168459, 32'sd0.1038102715009231, 32'sd0.1059411051317766, 32'sd0.09681746584414776, 32'sd0.027756257031278514, 32'sd-0.017155106675915334, 32'sd-0.00790994098436735, 32'sd0.09894081850164303, 32'sd-0.08402690350797862, 32'sd-0.03541742518773503, 32'sd0.11741738661053443, 32'sd0.06666869027374316, 32'sd0.04426444233884565, 32'sd-0.003211982232021251, 32'sd-0.06085212561831092, 32'sd0.0015449168355293828, 32'sd0.11513233875131051, 32'sd0.06623374007380514, 32'sd0.06978742517418499, 32'sd-0.008673374666531172, 32'sd0.12655373140108542, 32'sd-0.021818905837313555, 32'sd-0.01977053694194235, 32'sd-0.009109020697677859, 32'sd0.05422475188164887, 32'sd0.043011294637273406, 32'sd0.01446531366320952, 32'sd-0.014820003499794116, 32'sd0.07323976410148184, 32'sd0.12555891253330634, 32'sd0.0689350383490246, 32'sd0.026731151156184088, 32'sd-0.004177988885721284, 32'sd0.02029563631168378, 32'sd-0.024494045998252733, 32'sd0.10291202978798297, 32'sd-0.0757203960807386, 32'sd0.012682501322048583, 32'sd0.013413012615047086, 32'sd0.04669547835123703, 32'sd-0.08707729305861212, 32'sd-0.026095571994545354, 32'sd-0.0005070923092125771, 32'sd0.11345964042407512, 32'sd0.08327132168888099, 32'sd-0.09083434008406427, 32'sd0.058567545379282764, 32'sd0.07468120957595215, 32'sd0.09388547721924921, 32'sd-0.09670780405863466, 32'sd0.012538050352181354, 32'sd0.03755309550873881, 32'sd-0.09543565402374724, 32'sd-0.05139242011734946, 32'sd-0.0751946290147897, 32'sd-0.01991733585304039, 32'sd-0.024211609606516093, 32'sd-0.08031628353436064, 32'sd-0.02817013465487019, 32'sd0.09695394919384795, 32'sd-0.01129981467401851, 32'sd0.016056558049446838, 32'sd-0.002993082509579374, 32'sd-0.03717622378416446, 32'sd-0.01184634970707225, 32'sd0.02389590309753105, 32'sd0.06759601278431561, 32'sd-2.6113398693960706e-124, 32'sd-0.04460188902818885, 32'sd-0.027686343176579906, 32'sd0.013438231265444904, 32'sd0.060736855973496914, 32'sd-0.07231581616808305, 32'sd0.03069998267054107, 32'sd-0.03008539690902754, 32'sd0.0034791317100061965, 32'sd0.0728130088656971, 32'sd-0.09502108419252028, 32'sd0.03523520258044093, 32'sd0.045801390715168845, 32'sd-0.045076591173503475, 32'sd-0.11767445504718944, 32'sd-0.08709540889217517, 32'sd-0.03588768639319811, 32'sd-0.1032211909396923, 32'sd-0.06650287948579274, 32'sd-0.08643595790051505, 32'sd-0.0003863610766019354, 32'sd0.012576382308334876, 32'sd0.07192812199770364, 32'sd0.022291401347395042, 32'sd-0.01457859419541391, 32'sd0.04534584333188955, 32'sd-0.016745896116576894, 32'sd-7.348282596970499e-115, 32'sd-2.3824439138329073e-121, 32'sd-8.602559370586781e-128, 32'sd0.06911022871756298, 32'sd0.003869340141201307, 32'sd0.1073226169932097, 32'sd-0.0019573312631278057, 32'sd-0.06941842420358517, 32'sd-0.029973069800578133, 32'sd0.05193161893485603, 32'sd0.0008754630742594064, 32'sd-0.034797593323543305, 32'sd-0.03866225051131717, 32'sd0.006389076116787019, 32'sd-0.14237826576035464, 32'sd-0.2899335388072497, 32'sd-0.2032587997390038, 32'sd-0.05226368970158463, 32'sd0.015518383172515698, 32'sd0.008322233859678351, 32'sd-0.028352613045689357, 32'sd0.01775199808453831, 32'sd0.009750303847998567, 32'sd0.012878225047280282, 32'sd0.023896612687292047, 32'sd-0.04041704255660727, 32'sd0.009996479660322372, 32'sd-0.012914227101722192, 32'sd1.6679038189782584e-116, 32'sd4.284868424958e-125, 32'sd-8.528231774407352e-125, 32'sd-0.06770380098502117, 32'sd-0.02904719994827475, 32'sd0.08735537103025362, 32'sd0.036211152417934114, 32'sd0.1109798688919277, 32'sd0.06813609404134115, 32'sd-0.018342056621361905, 32'sd0.06211566722596587, 32'sd0.07624103432757927, 32'sd-0.04553170737705818, 32'sd-0.02302973289236963, 32'sd-0.03165196888608371, 32'sd0.005256315617638478, 32'sd-0.054884506974483285, 32'sd0.048225236535005, 32'sd0.07914405046074545, 32'sd0.056121685686510256, 32'sd-0.1459671298932664, 32'sd-0.07707663860100333, 32'sd0.0905048989602846, 32'sd0.09891870001223603, 32'sd-0.0249134775907329, 32'sd0.01779274888259634, 32'sd0.07194370955068387, 32'sd0.0711458927292369, 32'sd8.161035306496798e-122, 32'sd1.7168158773846857e-123, 32'sd1.0269919365387187e-121, 32'sd-3.724240034482763e-126, 32'sd0.07047662005178378, 32'sd-0.012382040891748339, 32'sd0.0604782269146339, 32'sd0.01500556802140573, 32'sd-0.064289004597972, 32'sd-0.017659840117428632, 32'sd0.07447974825461526, 32'sd0.05599653130153232, 32'sd-0.042632460377512095, 32'sd0.06304524433414949, 32'sd0.06220199310946347, 32'sd0.10773342533876312, 32'sd0.13286619773810396, 32'sd-0.05339546294325269, 32'sd0.0013713668247855955, 32'sd0.04789832079405983, 32'sd0.034150922972168894, 32'sd-0.07381427059644918, 32'sd-0.005492740462061191, 32'sd0.05107423598975718, 32'sd-0.006222463745681788, 32'sd0.016515964182795648, 32'sd0.06541222937828868, 32'sd1.9315544459593482e-114, 32'sd-6.085878568819948e-127, 32'sd1.793753942179389e-123, 32'sd5.806633035312686e-121, 32'sd2.2645110129742927e-115, 32'sd1.6341889002256245e-121, 32'sd0.09441671545136787, 32'sd0.09955836966345416, 32'sd0.05705244606500251, 32'sd0.08783382188100608, 32'sd0.0060626910502522315, 32'sd0.06390660435051772, 32'sd0.10280819351231525, 32'sd0.12730860043983389, 32'sd0.1902492688701758, 32'sd0.15171829481315321, 32'sd0.12461685921710805, 32'sd0.08791215698398454, 32'sd0.10958444120046153, 32'sd-0.001070245996446652, 32'sd-0.007526146944545699, 32'sd-0.0029639102639999098, 32'sd-0.003924896107102719, 32'sd0.003823467423232518, 32'sd0.10690077697215454, 32'sd0.013322149972554908, 32'sd2.3270201473248344e-122, 32'sd-2.461081212637581e-123, 32'sd-4.6887618587519825e-120, 32'sd-1.796201645266979e-123},
        '{32'sd-3.1008274667221346e-123, 32'sd2.2850965366839163e-115, 32'sd-9.947707866201858e-126, 32'sd1.8246122010326334e-126, 32'sd-5.941127432204221e-131, 32'sd8.901414262368495e-127, 32'sd2.8161012467889146e-124, 32'sd2.5168769112229107e-124, 32'sd-5.179777469032377e-124, 32'sd2.7110254085209623e-125, 32'sd1.3453102677282444e-114, 32'sd1.7223758274047342e-125, 32'sd0.06040130676564822, 32'sd0.047207932742327686, 32'sd-0.06126910963975987, 32'sd-0.02445874083811529, 32'sd3.417664060853493e-125, 32'sd2.0655547399296683e-124, 32'sd1.1081111504786104e-121, 32'sd-3.726084217244693e-125, 32'sd-5.6572305262576335e-121, 32'sd4.32042261667573e-125, 32'sd-3.3411603533469446e-122, 32'sd1.0373673367871611e-126, 32'sd-5.29412646072206e-118, 32'sd-6.380587455608983e-118, 32'sd-2.853410490346156e-114, 32'sd2.5109256216681408e-126, 32'sd-3.641325209480865e-129, 32'sd-1.3315607583220018e-122, 32'sd2.057187606421218e-117, 32'sd-6.900823420669728e-123, 32'sd0.10835008070006276, 32'sd0.06014537280284235, 32'sd-0.04745944153755541, 32'sd-0.03508799825875686, 32'sd-0.02749608927388442, 32'sd0.049281224994650284, 32'sd0.05529148481791099, 32'sd-0.02901852974926035, 32'sd0.06077899257800889, 32'sd-0.03189559157473784, 32'sd0.011575370730342345, 32'sd0.008765599834884587, 32'sd0.04572346924136598, 32'sd0.04006310229335363, 32'sd0.06920834644954782, 32'sd-0.018042001865758484, 32'sd0.038991444547027784, 32'sd-0.008593519673196876, 32'sd-0.05080619570644615, 32'sd0.0055502509393081665, 32'sd7.009950263168324e-119, 32'sd-1.8132760899523774e-122, 32'sd-1.6945971796984408e-122, 32'sd6.451207335225858e-117, 32'sd-7.873593083378788e-129, 32'sd2.7469967895213266e-129, 32'sd0.010029491455967843, 32'sd-0.047493527012259076, 32'sd0.03993273768109472, 32'sd-0.015926354098452885, 32'sd-0.05056062057653142, 32'sd0.08025175414750994, 32'sd-0.008327750152939758, 32'sd0.017019524200057135, 32'sd0.022796209647457644, 32'sd-0.038392898380321096, 32'sd0.04288368873904994, 32'sd-0.07989361471562541, 32'sd-0.0334663883823628, 32'sd-0.014202174911780845, 32'sd-0.05547829770014854, 32'sd-0.017608679070858252, 32'sd-0.08645879918358396, 32'sd0.08244157906475912, 32'sd0.06756147889369968, 32'sd0.030582943996695602, 32'sd-0.03973086959474398, 32'sd0.03969922991526278, 32'sd-0.009995108812879416, 32'sd0.016319245293850405, 32'sd-2.0412077641265807e-122, 32'sd1.0913653414961354e-117, 32'sd-2.169097115305513e-125, 32'sd2.8421174481870286e-120, 32'sd-0.02007843612388996, 32'sd-0.0781745864381317, 32'sd0.13519537852828928, 32'sd-0.05231827547698842, 32'sd0.009827603260464104, 32'sd-0.011759885570275293, 32'sd-0.0009732108492030282, 32'sd-0.006974796366972298, 32'sd0.06725474031233428, 32'sd-0.025689198551000842, 32'sd-0.15805330409468216, 32'sd-0.04066552491432181, 32'sd0.047171686792829924, 32'sd0.029983233779208713, 32'sd0.04747407317051814, 32'sd-0.007609142559640947, 32'sd0.12846871342395105, 32'sd0.09643761627795398, 32'sd0.01777800605998052, 32'sd0.03144971569868458, 32'sd0.0012585251017742582, 32'sd0.006095305359125446, 32'sd0.05227198513531041, 32'sd-0.0702321809296506, 32'sd-0.05522048799084779, 32'sd1.30365833664537e-125, 32'sd-2.1060440611299864e-114, 32'sd0.04656806523765227, 32'sd0.0701941629618746, 32'sd0.03158732776055311, 32'sd0.024670327669848103, 32'sd-0.015685197233337864, 32'sd-0.00962775018018465, 32'sd-0.028950838351069905, 32'sd-0.15496659294635695, 32'sd-0.05951842364028277, 32'sd0.005100796532918886, 32'sd0.02754085513110485, 32'sd0.09704567371034259, 32'sd0.0074617256326978245, 32'sd0.05379353779216036, 32'sd-0.02231261086775469, 32'sd0.09820674723355981, 32'sd-0.07762622960048059, 32'sd0.029683194916042304, 32'sd0.06736966456887476, 32'sd0.058194305323749466, 32'sd-0.00017503671341439106, 32'sd0.010119654925530365, 32'sd-0.06806343409641921, 32'sd-0.0803558303022159, 32'sd0.004656330430271301, 32'sd0.006665122389559458, 32'sd8.639257354709183e-05, 32'sd-1.8480645981701383e-116, 32'sd-0.004443409571828919, 32'sd-0.08017187183766786, 32'sd-0.05203197125470375, 32'sd-0.09944518962187965, 32'sd-0.08607536009605724, 32'sd0.003285213742763822, 32'sd-0.03569623034598596, 32'sd-0.03605326516356289, 32'sd0.03739344227453221, 32'sd0.038934856953039526, 32'sd0.03975766939700659, 32'sd0.001513719697106667, 32'sd0.01193258465723166, 32'sd-0.08006555897034666, 32'sd-0.08509683793659077, 32'sd-0.05803758114074451, 32'sd0.10427239443468024, 32'sd0.01609938315658899, 32'sd0.04464258011537436, 32'sd-0.08434146793675543, 32'sd0.06221500120885994, 32'sd0.09760313013886651, 32'sd-0.04144666733211313, 32'sd0.07166250264184035, 32'sd-0.07759808346848429, 32'sd0.03219483001752919, 32'sd-0.05709581412828409, 32'sd5.837084479564791e-125, 32'sd-0.03152264311013917, 32'sd0.00243754450686287, 32'sd-0.030337203313102443, 32'sd0.010313170694932853, 32'sd0.052062848714803905, 32'sd-0.1412381481657696, 32'sd-0.03286756111135107, 32'sd-0.041125344380488836, 32'sd0.0055343603348049575, 32'sd0.04254475330520874, 32'sd0.1562538426759269, 32'sd0.02021670301226295, 32'sd0.035132742478268454, 32'sd-0.04664583716152497, 32'sd-0.14987017991761445, 32'sd-0.1754535709317356, 32'sd0.028782623553971234, 32'sd0.052525716137151214, 32'sd0.06994441478004913, 32'sd0.0753752230017163, 32'sd-0.1320439560548174, 32'sd0.025333110587638503, 32'sd0.06593406825408303, 32'sd-0.049475413475231704, 32'sd0.007391329131339558, 32'sd0.030408906004051304, 32'sd0.10128335356936, 32'sd0.01164986957091769, 32'sd0.05455287575417241, 32'sd0.020290925362663706, 32'sd-0.16757183757358102, 32'sd-0.04692559510693171, 32'sd-0.04176507470406195, 32'sd-0.1425758034713297, 32'sd0.017619058486375648, 32'sd0.08704871945011514, 32'sd0.10936230573839673, 32'sd0.022619846257977298, 32'sd0.04862426531396626, 32'sd-0.0996892378497157, 32'sd-0.04387198743449093, 32'sd0.04669855234933246, 32'sd-0.014072289271308283, 32'sd-0.15864574157477018, 32'sd-0.08105596388263081, 32'sd0.10878882409540445, 32'sd0.07239308751250412, 32'sd0.05271804447765471, 32'sd0.11391346521081559, 32'sd0.09051026222750003, 32'sd0.005998217335909052, 32'sd-0.08592218913888135, 32'sd-0.03819839166729573, 32'sd0.009049392224750458, 32'sd-0.017539998951231248, 32'sd-0.02183876503468907, 32'sd0.015712686298280435, 32'sd0.06939504723459043, 32'sd-0.07593111803468779, 32'sd-0.039832340551783085, 32'sd-0.11203920850135904, 32'sd0.027058566116980137, 32'sd0.05589495247570614, 32'sd0.057513173305332906, 32'sd0.1126262197174413, 32'sd-0.04209606539633977, 32'sd-0.06275600081804293, 32'sd-0.05741486691822434, 32'sd0.012413595359762868, 32'sd-0.02216532664953351, 32'sd0.09112656636432778, 32'sd-0.04187713040620113, 32'sd0.022031545338225628, 32'sd0.04975480482834752, 32'sd-0.045456980505893245, 32'sd-0.037955995155054295, 32'sd0.06511466790786798, 32'sd0.05940871287169927, 32'sd0.02158218522533095, 32'sd0.04409944951953474, 32'sd0.033770556680652104, 32'sd-0.04090519968384322, 32'sd-0.047400184158411275, 32'sd-0.05513663385700754, 32'sd-0.05919572185725988, 32'sd0.09317182975866727, 32'sd0.037851927041519, 32'sd-0.05788689867916514, 32'sd-0.13683005493228162, 32'sd-0.13092262709266456, 32'sd0.066995441445435, 32'sd0.14021802898057115, 32'sd-0.00871915040077496, 32'sd0.05606668842591097, 32'sd0.10041989738856201, 32'sd-0.11852219456224448, 32'sd-0.18081463301217443, 32'sd-0.0030034754819024266, 32'sd-0.12612504443914746, 32'sd0.011719730451259595, 32'sd-0.08719704884866862, 32'sd-0.14945662247226937, 32'sd-0.1508689944333582, 32'sd-0.18182491397744585, 32'sd-0.04344244628792335, 32'sd-0.04745439717218051, 32'sd-0.06723866688724954, 32'sd-0.15025787310302435, 32'sd-0.19657928963907148, 32'sd-0.01283277643472015, 32'sd-0.0562264312550615, 32'sd-0.037789312230355546, 32'sd-0.055476603963874695, 32'sd0.02944781144908582, 32'sd-0.009497009937980154, 32'sd-0.039146260189668144, 32'sd-0.09597080959642859, 32'sd-0.06582176161485793, 32'sd0.11460114841495507, 32'sd0.13657340386049657, 32'sd0.15838328512667194, 32'sd0.12551558720839698, 32'sd0.10907105455076524, 32'sd0.011174667182014628, 32'sd-0.21529957042764156, 32'sd-0.27748952421518647, 32'sd-0.13895174534120158, 32'sd0.08591234794485166, 32'sd-0.04922972847113717, 32'sd-0.03670203362901119, 32'sd-0.004682874660756374, 32'sd-0.044607995806091316, 32'sd-0.11643131580476533, 32'sd-0.09422954143260036, 32'sd-0.07528948358227118, 32'sd-0.021479876074953566, 32'sd-0.13023151291988944, 32'sd-0.000859910193077554, 32'sd0.03437961082574914, 32'sd0.06165189060646882, 32'sd0.14246478335449958, 32'sd-0.0015625532592735546, 32'sd0.0168378246661745, 32'sd0.010263885391135442, 32'sd-0.09675425725914039, 32'sd-0.07888393832917495, 32'sd0.12155385420082358, 32'sd0.1439514566168918, 32'sd0.20312031400578145, 32'sd0.19645396651560473, 32'sd0.053522587798066616, 32'sd-0.09432452930587476, 32'sd-0.12777543786742418, 32'sd-0.04373193383210286, 32'sd0.04947923345993372, 32'sd0.08918799910080359, 32'sd0.06589309998505034, 32'sd0.07049068008424961, 32'sd-0.019682375787744764, 32'sd-0.08407490917866975, 32'sd-0.06593202275039263, 32'sd-0.10000308424202707, 32'sd-0.12881815583108866, 32'sd0.028709762796680343, 32'sd-0.14641398247293666, 32'sd-0.0777978827997206, 32'sd-0.00715872511202142, 32'sd0.0019708928294123193, 32'sd-0.07156388731044422, 32'sd-0.09364790865730568, 32'sd0.03747867162874912, 32'sd-0.01611757109922972, 32'sd-0.09702026052135015, 32'sd-0.09207784091603774, 32'sd-0.023285445056491657, 32'sd0.1556954418216269, 32'sd0.26778765452744063, 32'sd0.045488133216973606, 32'sd0.048499295590275854, 32'sd-0.0334225956571992, 32'sd-0.15702785102461758, 32'sd-0.08126012454539616, 32'sd0.13954720896555384, 32'sd0.09160792961651866, 32'sd0.06614005828574965, 32'sd0.027943250281079503, 32'sd0.05436382781286001, 32'sd0.014311527907608826, 32'sd0.045146401278008626, 32'sd0.010819737767270942, 32'sd-0.09760957313777743, 32'sd0.012377210451674439, 32'sd0.045537233048758785, 32'sd-0.1425293083236841, 32'sd-0.023013740094970845, 32'sd-0.014974861919474232, 32'sd-0.027602650088067896, 32'sd3.9660549354015765e-05, 32'sd-0.019440259341307498, 32'sd0.024366817007508722, 32'sd-0.05633754503788712, 32'sd-0.05409223810367491, 32'sd0.0835341489199964, 32'sd0.04298517717023119, 32'sd0.2512501005329735, 32'sd0.12536195108504608, 32'sd-0.06629859115834381, 32'sd-0.07567964282534005, 32'sd-0.08984465947642939, 32'sd0.018295950912798335, 32'sd0.17316109562341267, 32'sd-0.05537228011195619, 32'sd-0.12084324424179323, 32'sd0.048033307771907986, 32'sd0.05035345691388908, 32'sd0.14473288868734915, 32'sd-0.05189946508926753, 32'sd0.06180830289149739, 32'sd0.08999228999370716, 32'sd0.05203235294598858, 32'sd0.11882793178691729, 32'sd-0.050825326898725896, 32'sd0.015447836109908708, 32'sd0.03379279173384949, 32'sd-0.03501050406190904, 32'sd0.017425789570601948, 32'sd-0.11123095286424725, 32'sd-0.05483728640509889, 32'sd0.037105220007106456, 32'sd-0.03712882702400782, 32'sd0.06589912294313613, 32'sd0.13996948374529292, 32'sd0.12176299311454361, 32'sd0.18732505050581255, 32'sd0.0929744832284864, 32'sd-0.03086865782288439, 32'sd-0.0251986014989245, 32'sd0.043229913029423014, 32'sd-0.11361356566639855, 32'sd0.01618078933964432, 32'sd0.0930789181268787, 32'sd0.06634266224792265, 32'sd-0.005234084684430251, 32'sd0.10092324753992447, 32'sd0.03576304176788649, 32'sd0.11844135308535338, 32'sd0.12045943617717321, 32'sd0.03859859411132783, 32'sd0.04253789013974186, 32'sd-0.06669881151029713, 32'sd-0.058085277890423996, 32'sd-0.07262209554242056, 32'sd-0.028433546257231764, 32'sd-0.09287820823920012, 32'sd-0.034034603246821546, 32'sd-0.03757662990787371, 32'sd0.020113764195257917, 32'sd-0.14821873645884004, 32'sd-0.0406947235403989, 32'sd0.12120481406015933, 32'sd0.17217167037181044, 32'sd0.20333469917615993, 32'sd0.12940351693865823, 32'sd0.19120019532531926, 32'sd0.023699427644405423, 32'sd-0.06552243505385372, 32'sd-0.11478867315929253, 32'sd-0.09592785397854885, 32'sd0.00358205692180189, 32'sd0.0148990502110667, 32'sd-0.02762926067123304, 32'sd0.1553057948796111, 32'sd0.07644954284104459, 32'sd-0.09834579098720954, 32'sd0.060165411021552206, 32'sd0.04237785058966004, 32'sd0.025879757320654253, 32'sd0.01460383576247296, 32'sd-0.07081244655890999, 32'sd0.024725989421162945, 32'sd0.010694169870419079, 32'sd-0.057734069920332906, 32'sd-0.04598524220786152, 32'sd0.08147501597665043, 32'sd-0.12062601655943232, 32'sd-0.17956119633059062, 32'sd-0.15118106828547015, 32'sd0.15623484218834457, 32'sd0.012067221314471408, 32'sd0.08588533047301863, 32'sd0.15378447811931173, 32'sd0.09640097931682806, 32'sd-0.0597099245238451, 32'sd-0.1734585470709183, 32'sd-0.030748080488206476, 32'sd0.008254937781135193, 32'sd0.007704794212323475, 32'sd-0.05705489090847397, 32'sd0.12814754161342248, 32'sd-0.018966027551738755, 32'sd-0.002885139449364238, 32'sd-0.10282565551555863, 32'sd0.017912848208537804, 32'sd-0.10134211372501584, 32'sd0.05493263674515202, 32'sd-0.10297117743976143, 32'sd0.0571561564575919, 32'sd3.8275936546492036e-121, 32'sd0.0033050514653580852, 32'sd0.031015101679980055, 32'sd0.0031136822879404254, 32'sd0.011646282168173056, 32'sd-0.13466689430110404, 32'sd-0.09095461654355931, 32'sd-0.16013502726393108, 32'sd0.03630643985116807, 32'sd-0.04000572945677692, 32'sd0.12804174178141975, 32'sd0.19538962955983596, 32'sd0.221484669055395, 32'sd0.08680341353515555, 32'sd-0.089550035316978, 32'sd-0.16959974703881786, 32'sd-0.1255499225579886, 32'sd-0.08097306493606153, 32'sd0.0025826245614921344, 32'sd0.09171903686239799, 32'sd-0.05238445546965393, 32'sd-0.05231902200472349, 32'sd-0.030814204185151465, 32'sd-0.001875575312930085, 32'sd0.05542641727116128, 32'sd0.0009383317739893401, 32'sd0.05343777501618592, 32'sd0.021463792985805252, 32'sd-0.027489115058602485, 32'sd-0.022941775578638784, 32'sd0.04060521100067226, 32'sd0.01247353354361198, 32'sd-0.029559008533064937, 32'sd-0.18220387148547945, 32'sd-0.15085651229336022, 32'sd-0.10082040402834629, 32'sd-0.06924444759140519, 32'sd0.13563500248125843, 32'sd0.060716462968038065, 32'sd-0.0737461582275175, 32'sd0.08301213616959666, 32'sd-0.00468920752817519, 32'sd-0.0994712271049089, 32'sd-0.0767740684758775, 32'sd-0.13416190030446848, 32'sd0.0265915159324904, 32'sd0.019115775278145255, 32'sd0.0812699511925784, 32'sd0.009422381672718855, 32'sd-0.03257577333498791, 32'sd-0.013590292729502103, 32'sd0.011404970709750247, 32'sd-0.029644787808646343, 32'sd0.010952005878126688, 32'sd0.0599754040373328, 32'sd-0.01894998589578998, 32'sd-0.03657205541179041, 32'sd-0.056714047938790264, 32'sd-0.05191820280168799, 32'sd-0.0738053452609465, 32'sd-0.07192007285032367, 32'sd-0.010742301927311177, 32'sd-0.03214085352416777, 32'sd-0.06847886040439284, 32'sd-0.08573369964009465, 32'sd-0.03603266556214545, 32'sd-0.07627827424226812, 32'sd-0.0183354322534887, 32'sd0.019192500677826137, 32'sd0.10290029866313512, 32'sd0.0034871437122487386, 32'sd-0.14347927643716935, 32'sd-0.1824042435352711, 32'sd0.010897890204588456, 32'sd0.1348451632394027, 32'sd0.025409127370787814, 32'sd-0.014678903206262273, 32'sd-0.15973613747672913, 32'sd0.05712948408456416, 32'sd0.06261987728779633, 32'sd0.050115484665931284, 32'sd-0.027952626831453473, 32'sd-0.03364837071147684, 32'sd-0.11652567618435211, 32'sd1.6824737488983968e-123, 32'sd-0.027508970100342336, 32'sd-0.051645443868724494, 32'sd-0.04560096870576313, 32'sd-0.024718561251416832, 32'sd-0.07169162928087608, 32'sd-0.044749575791089374, 32'sd-0.2012157594797257, 32'sd-0.057109136014835915, 32'sd-0.11262196061039743, 32'sd-0.12720826928047965, 32'sd0.04576183783262254, 32'sd0.04398943570144351, 32'sd0.04375833701217174, 32'sd-0.04438957286916606, 32'sd-0.07247786924389335, 32'sd0.045440109840578086, 32'sd0.11754731486165049, 32'sd0.14043035253060682, 32'sd0.025438290937221896, 32'sd-0.051104133879143115, 32'sd-0.0431189498235149, 32'sd0.021618791333149402, 32'sd-0.02342323619326005, 32'sd-0.03723527539000723, 32'sd-0.021361806828645816, 32'sd-0.08576055302296563, 32'sd0.03855603792356229, 32'sd-0.03955413153551402, 32'sd-0.02815966633290465, 32'sd0.019820630971776783, 32'sd-0.09666495655075154, 32'sd-0.010089609432243275, 32'sd0.08073640425352688, 32'sd-0.11439662257077715, 32'sd-0.18923580288115202, 32'sd-0.0970757413549004, 32'sd-0.002656390340543576, 32'sd-0.10927660194995453, 32'sd-0.06307454908987195, 32'sd0.15287537662820586, 32'sd-0.004705058716544457, 32'sd0.02688018069735795, 32'sd-0.09913123517228141, 32'sd-0.057901423427054004, 32'sd0.07191462104405799, 32'sd0.1332308949078866, 32'sd0.006070671898871812, 32'sd0.08739020875754419, 32'sd-0.030480241915748527, 32'sd0.08096017001660215, 32'sd0.010914686840493794, 32'sd-0.06610167314546288, 32'sd-0.022243318061789138, 32'sd0.0459538546483412, 32'sd-0.07178449289322256, 32'sd-0.04097754586178916, 32'sd0.08537660701067876, 32'sd0.050488676239858386, 32'sd0.008027692391049479, 32'sd-0.04892633456482116, 32'sd0.017279622193187603, 32'sd-0.16313756245735156, 32'sd-0.18622058261319577, 32'sd-0.14032061227860557, 32'sd-0.07178815512505127, 32'sd0.05239851310799167, 32'sd0.0014714699145862062, 32'sd0.014667993393916117, 32'sd-0.061988461828930905, 32'sd-0.0031626471845040377, 32'sd0.0737663598031634, 32'sd0.14485402919232213, 32'sd0.06506111585794476, 32'sd0.07188161755792, 32'sd0.0648102991593026, 32'sd-0.03285325801299435, 32'sd0.010941754688220468, 32'sd-0.1229052115291635, 32'sd-0.06875974067139337, 32'sd-0.08314910148357123, 32'sd0.04302718641043036, 32'sd-0.030201237892049173, 32'sd0.04401556033234183, 32'sd-1.1109774148466724e-119, 32'sd0.011780896868805627, 32'sd-0.06838607054360436, 32'sd0.07455996291757123, 32'sd-0.05466763415405865, 32'sd0.0825772919633506, 32'sd-0.04070102739682267, 32'sd-0.04843874410083334, 32'sd-0.06042740279876114, 32'sd0.003456331774398446, 32'sd0.03217435457002352, 32'sd-0.03206585411955171, 32'sd0.06107565082483633, 32'sd0.017020441675805405, 32'sd0.054558862864524556, 32'sd0.11529778396823565, 32'sd0.16207586102466107, 32'sd0.08028347040373572, 32'sd-0.03676421440278588, 32'sd-0.11132504918078062, 32'sd-0.10568189828497472, 32'sd0.006523612448784171, 32'sd-0.1640814736189574, 32'sd0.016707099376866937, 32'sd0.03173708999247779, 32'sd0.05009703596990667, 32'sd0.03822286892453172, 32'sd-4.658395507336909e-123, 32'sd-1.4208776912847905e-118, 32'sd6.138945361213193e-126, 32'sd0.014570361969588252, 32'sd-0.008943818340078872, 32'sd-0.060009979711937264, 32'sd-0.060463995946157444, 32'sd-0.0877673987141074, 32'sd0.027078581901233776, 32'sd0.005852631730151635, 32'sd-0.019967104376369827, 32'sd-0.04328506565202905, 32'sd0.052426675145114454, 32'sd-0.06682693005131203, 32'sd0.02175363364385039, 32'sd-0.023147491691426183, 32'sd-0.016884196260561705, 32'sd-0.022652574828918026, 32'sd-0.10232146483437818, 32'sd-0.14563155085736007, 32'sd-0.028001890579207878, 32'sd0.011303021112900128, 32'sd0.024445005327075296, 32'sd-0.02072911138021722, 32'sd-0.018453415094550136, 32'sd-0.024579539949903292, 32'sd-0.09116923983275035, 32'sd-0.026082734834144708, 32'sd-3.592811951708722e-116, 32'sd1.9070925615006137e-114, 32'sd1.0761996235546008e-118, 32'sd0.017625618689826435, 32'sd0.03748151365577539, 32'sd-0.011598343856757985, 32'sd-0.042590156847339716, 32'sd0.04181087861107716, 32'sd0.006477154689445872, 32'sd0.013837313892589641, 32'sd0.16624948118669988, 32'sd-0.008792756728585049, 32'sd-0.08397592814713845, 32'sd-0.1449796563069975, 32'sd-0.12589521534417678, 32'sd-0.011438661199076643, 32'sd-0.0804466072095679, 32'sd-0.013154463588830061, 32'sd0.09935701007766948, 32'sd0.1169052050260296, 32'sd-1.738407630041558e-05, 32'sd-0.035488757044328786, 32'sd-0.028974589628600108, 32'sd0.06410775126307691, 32'sd0.04188425473900251, 32'sd-0.05704216734638261, 32'sd-0.052477460221413905, 32'sd0.025679479805476198, 32'sd1.5386758798958606e-120, 32'sd3.597872618653621e-119, 32'sd1.0432679315581715e-115, 32'sd2.546627474010807e-115, 32'sd-0.009031189132088786, 32'sd-0.02686048973342578, 32'sd-0.00874571839213391, 32'sd0.04960590015388188, 32'sd0.03741534487392712, 32'sd0.07148803812112717, 32'sd0.019592906500647784, 32'sd0.03558788178799626, 32'sd0.06506876315420387, 32'sd-0.00499756721091063, 32'sd0.0401945452784605, 32'sd-0.024677006648999994, 32'sd-0.15445260416596393, 32'sd-0.10619206761029086, 32'sd-0.023043954180722023, 32'sd-0.002013083597711654, 32'sd-0.004112348562652637, 32'sd-0.06040717830230203, 32'sd0.024807831482773674, 32'sd0.05187695623782118, 32'sd0.07401634706855699, 32'sd-0.02890882698598563, 32'sd-0.02645398184343196, 32'sd-4.380985027692734e-121, 32'sd2.912494215340664e-127, 32'sd8.329127219761118e-118, 32'sd-1.8280891655272203e-117, 32'sd-9.01648349592374e-120, 32'sd2.4968616843477513e-124, 32'sd-0.043096537390550374, 32'sd-0.026658689951139427, 32'sd0.09739337308601886, 32'sd0.027695034267389344, 32'sd0.0035592615038518302, 32'sd-0.040133235881545375, 32'sd-0.014051668389033467, 32'sd0.06983428866922942, 32'sd0.09302896379115802, 32'sd0.09319300813364158, 32'sd-0.0039692625725933186, 32'sd-0.04010685529111535, 32'sd-0.06212867339239513, 32'sd-0.01411131453536655, 32'sd-0.07746534667635221, 32'sd-0.04782933322903003, 32'sd0.006830617605585998, 32'sd-0.06604075765954252, 32'sd-0.07838050127852882, 32'sd0.020569362446734598, 32'sd1.3413755706898356e-122, 32'sd-2.2679800262421764e-120, 32'sd-8.294587375117341e-122, 32'sd-1.5097063185143577e-123},
        '{32'sd-1.192353315440166e-118, 32'sd5.41127985039343e-126, 32'sd6.995519029253768e-123, 32'sd-1.616114341160768e-116, 32'sd-6.873133440181915e-128, 32'sd4.223203288388636e-128, 32'sd9.652098383422728e-121, 32'sd1.5376468187587064e-121, 32'sd6.555670743200737e-120, 32'sd9.957919751545956e-124, 32'sd-4.067292866569673e-124, 32'sd-3.256623771335323e-120, 32'sd-0.09048443912656269, 32'sd0.009175019571669442, 32'sd-0.025975999550947773, 32'sd-0.0023320181121335866, 32'sd3.2140827802820636e-121, 32'sd1.6797330804930003e-127, 32'sd2.5609499589589575e-124, 32'sd2.0720306039277215e-127, 32'sd-1.9712418282890098e-118, 32'sd-5.637221752618692e-125, 32'sd1.3415445474148676e-117, 32'sd-2.0233574854632917e-121, 32'sd6.545769260613753e-115, 32'sd-1.764176336022428e-123, 32'sd-7.885957551189971e-118, 32'sd-6.361202856662134e-124, 32'sd8.670610359592356e-121, 32'sd3.242967537034593e-123, 32'sd4.2110999186464783e-125, 32'sd3.289065188225552e-119, 32'sd0.0446000393546715, 32'sd0.04599785932450842, 32'sd-0.01941436197133868, 32'sd-0.056515346296795194, 32'sd-0.11436293300477561, 32'sd-0.03223908311148313, 32'sd0.10320789502097132, 32'sd0.07573934466506158, 32'sd0.09815724177247266, 32'sd0.08716529317147294, 32'sd0.12387920516756995, 32'sd0.10213177893101019, 32'sd0.007836390661902358, 32'sd0.04389732281590051, 32'sd0.09320447963216891, 32'sd0.018381645393935716, 32'sd0.036637546756056016, 32'sd0.0014569049343840226, 32'sd-0.00249331986327629, 32'sd0.022983897933155827, 32'sd-3.8158210824756296e-119, 32'sd-6.613859262232297e-124, 32'sd-6.937541419595263e-122, 32'sd1.0447264476960704e-120, 32'sd3.5638641987008284e-118, 32'sd-1.073714492586804e-124, 32'sd0.07381230399944338, 32'sd-0.015365199444135648, 32'sd0.07215521244464651, 32'sd-0.016773663765130693, 32'sd0.025532034261677158, 32'sd0.0033887636031137017, 32'sd0.04713374881415756, 32'sd-0.015177944066595306, 32'sd-0.02037148518226103, 32'sd-0.029060538059423643, 32'sd-0.10232106980109966, 32'sd0.01627571954836072, 32'sd0.13724941937424368, 32'sd0.06933764384493879, 32'sd0.024738623843061223, 32'sd0.047147768970591676, 32'sd-0.04458962702305729, 32'sd0.0010059957388444882, 32'sd0.04152292622189458, 32'sd0.06086955406241168, 32'sd0.049440673941085284, 32'sd0.05967350345214282, 32'sd0.0561872647344918, 32'sd0.0025223716340940167, 32'sd-3.1090530862936555e-120, 32'sd-2.5199359102760126e-124, 32'sd-6.401627639684468e-115, 32'sd3.6919796657344294e-127, 32'sd-0.029780594174057373, 32'sd0.029511396585892326, 32'sd-0.04443427127563953, 32'sd-0.006422844551868666, 32'sd-0.08483564236183927, 32'sd-0.043621311752470394, 32'sd-0.028857982257160276, 32'sd0.007257679182182312, 32'sd0.06741286057577725, 32'sd0.025641767534792616, 32'sd-0.06594444056543322, 32'sd0.10734808781810513, 32'sd0.08195070736355384, 32'sd0.0008402273495596037, 32'sd0.04627426297774361, 32'sd0.10442926873303104, 32'sd0.0774773237594162, 32'sd-0.010353985966235577, 32'sd0.0933413220680903, 32'sd0.03558654748486661, 32'sd0.04760503805984062, 32'sd-0.04629550045592937, 32'sd0.04006489681292091, 32'sd-0.05245757651762596, 32'sd0.0049910179715506155, 32'sd-4.323643869772065e-125, 32'sd2.8188370089330337e-122, 32'sd0.07202797601784287, 32'sd0.033950175785334, 32'sd-0.02302211281463805, 32'sd-0.13756649931394582, 32'sd-0.011002512978899117, 32'sd0.06047899158818597, 32'sd0.03814350614859645, 32'sd-0.0342354780099625, 32'sd0.1342276402252278, 32'sd0.07281512570994184, 32'sd0.006496975843566132, 32'sd-0.028270852013440952, 32'sd0.010544702569207046, 32'sd-0.015714721389836987, 32'sd-0.07790235921612224, 32'sd0.0299398129155316, 32'sd-0.07920231428925781, 32'sd0.013397918121849648, 32'sd0.07024465874548068, 32'sd0.14211650753469007, 32'sd-0.01803770068699998, 32'sd0.03418735661450519, 32'sd0.102759092654622, 32'sd-0.02744686038349014, 32'sd0.016361948717429145, 32'sd0.011272275071122223, 32'sd0.0494013752136692, 32'sd2.709124030907133e-115, 32'sd0.0219603621448606, 32'sd0.07923158822678024, 32'sd0.06635703309968706, 32'sd-0.010057204036160946, 32'sd-0.11404422230372549, 32'sd-0.028571042131716216, 32'sd-0.12140976378423962, 32'sd0.06409705897202621, 32'sd-0.0019299350576941455, 32'sd0.0752334535681844, 32'sd-0.010096728267433613, 32'sd-0.025386516882412814, 32'sd-0.019681691082425783, 32'sd-0.015836060593536875, 32'sd-0.010781754946971997, 32'sd-0.17240875991777363, 32'sd-0.12370844223641064, 32'sd-0.07053698906226168, 32'sd-0.011008287174372985, 32'sd-0.12710809880139198, 32'sd-0.1184561651646882, 32'sd-0.00999763770002498, 32'sd0.06690567067053674, 32'sd0.011434662123007625, 32'sd0.050057820804521966, 32'sd0.056044811159837275, 32'sd0.010582554896101343, 32'sd4.0408176186222243e-125, 32'sd0.050896631387871816, 32'sd0.03883643607857937, 32'sd0.04339718268330633, 32'sd0.08703185057003864, 32'sd0.040030004588330614, 32'sd0.08023601055096126, 32'sd0.08693920175901171, 32'sd-0.033377869038994076, 32'sd-0.0549319667372493, 32'sd-0.03811559885344072, 32'sd0.02687673314462735, 32'sd-0.0785871410737602, 32'sd-0.011420028733196511, 32'sd-0.08649501486532278, 32'sd-0.03329234689613403, 32'sd0.045503334082205575, 32'sd-0.046775398217230306, 32'sd-0.012648770518847496, 32'sd-0.08186379445056598, 32'sd-0.03156732851546979, 32'sd0.002168540944971431, 32'sd-0.030936528874751682, 32'sd0.04128641265831686, 32'sd-0.008523409692669341, 32'sd0.04311225870510337, 32'sd0.046625472615902656, 32'sd-0.06206327815387318, 32'sd0.05668265808587601, 32'sd0.00020929539691975373, 32'sd-0.0364927445678899, 32'sd-0.0834110964767149, 32'sd0.06575338364668752, 32'sd0.08959840436843045, 32'sd0.020906273238302464, 32'sd0.06192602268573528, 32'sd0.004505477981838457, 32'sd0.004411906171319657, 32'sd-0.04566651414331741, 32'sd-0.07818378446169855, 32'sd-0.004595676886111036, 32'sd-0.14074493327997156, 32'sd-0.1425235153151492, 32'sd0.02898468892588098, 32'sd0.08006112877565853, 32'sd0.05372679326544087, 32'sd0.017417043203059344, 32'sd-0.02190871192721524, 32'sd-0.02701045765562527, 32'sd0.01591306342829289, 32'sd0.018143746138359375, 32'sd0.025971513282426802, 32'sd0.11349859957018939, 32'sd-0.06147426773227484, 32'sd0.03592127337368238, 32'sd-0.010111304999196687, 32'sd0.010097183725430257, 32'sd0.0445702621542717, 32'sd0.015321395646053181, 32'sd0.050848743313361415, 32'sd0.07843124731551616, 32'sd0.03908278738574318, 32'sd-0.00026626921696792515, 32'sd0.12698925861842278, 32'sd0.1331682393329519, 32'sd0.10359176500631015, 32'sd0.0687088113916801, 32'sd0.04662454663622151, 32'sd-0.04942845509223248, 32'sd-0.1757383159678911, 32'sd0.017985727355913153, 32'sd0.11444121028548762, 32'sd0.23269474505478613, 32'sd0.04235099890918283, 32'sd0.009389350978254956, 32'sd0.01334457003145188, 32'sd-0.021170845297913406, 32'sd0.01651768063181013, 32'sd-0.013994335237229249, 32'sd-0.02485440388853413, 32'sd0.11189342699668052, 32'sd-0.09948526443612488, 32'sd-0.07139597005569233, 32'sd0.006069471372597109, 32'sd0.11186059275372114, 32'sd0.09166752304075348, 32'sd-0.0036946004502660594, 32'sd0.00582484830107439, 32'sd0.06471398648112325, 32'sd0.05966136394341815, 32'sd-0.043092633915766294, 32'sd0.029619583179731554, 32'sd0.13339660172878312, 32'sd0.02728391191309229, 32'sd0.11062901468949968, 32'sd-0.06336883819488869, 32'sd-0.2187081406477263, 32'sd-0.08034800918185812, 32'sd0.05686838994763913, 32'sd0.031018309736788482, 32'sd0.11088826349267844, 32'sd-0.0632313044089132, 32'sd0.05703873191590675, 32'sd0.1432177253106349, 32'sd0.1904017262802557, 32'sd0.02762835011729217, 32'sd0.039621982459496816, 32'sd0.07384916806181845, 32'sd-0.006725167544869182, 32'sd0.07315624458286529, 32'sd-0.03751943804630957, 32'sd-0.0019096198545200118, 32'sd0.1008268872073891, 32'sd-0.007769720496813974, 32'sd0.09128236049292958, 32'sd-0.06968415942701378, 32'sd0.1342653572433716, 32'sd0.06700095941638404, 32'sd-0.031083265602859147, 32'sd-0.029402271352255156, 32'sd0.05466295236785856, 32'sd0.06798725044220504, 32'sd0.12541875984605558, 32'sd0.13322171817113518, 32'sd-0.09132464447373796, 32'sd-0.09768861555773316, 32'sd-0.14072174529252326, 32'sd-0.022617186118526412, 32'sd0.07010586689173257, 32'sd0.001630007660912777, 32'sd0.12411116965093179, 32'sd0.09641905249919477, 32'sd0.11021862050514165, 32'sd0.06485733657525038, 32'sd0.08490476609150428, 32'sd0.023130000710903566, 32'sd0.031781323324418624, 32'sd-0.032479077243920615, 32'sd-0.045851524619820415, 32'sd-0.09188304517173133, 32'sd0.008081738274750486, 32'sd0.0018236106871009042, 32'sd-0.03627827759286548, 32'sd-0.011208933417480837, 32'sd0.03754667325715674, 32'sd0.0033121968015219863, 32'sd0.004660271430857343, 32'sd-0.0270917882127295, 32'sd0.0965697447409473, 32'sd0.19429657957626048, 32'sd0.10213913892444526, 32'sd0.14615998845457112, 32'sd-0.08245048142222518, 32'sd-0.20824808016112256, 32'sd-0.08099938460420704, 32'sd-0.09996204417089045, 32'sd-0.010765825330517339, 32'sd0.12568980175426706, 32'sd-0.010577951173045025, 32'sd0.021428589514574853, 32'sd0.10216145394716392, 32'sd-0.03071886657933299, 32'sd0.05191678027617735, 32'sd-0.017276066464505708, 32'sd0.04399720540171385, 32'sd0.01800647204996631, 32'sd-0.003031324915113224, 32'sd0.018186933626574843, 32'sd0.03618979891088467, 32'sd0.04719131369149304, 32'sd0.0758069400040811, 32'sd-0.028248844023316122, 32'sd-0.03647053650870769, 32'sd0.07938982330386177, 32'sd0.053833010892587026, 32'sd0.13503561518930446, 32'sd0.04158938906190219, 32'sd0.18215497980476242, 32'sd0.2432847927298892, 32'sd0.04543771366776882, 32'sd-0.021201640339201726, 32'sd-0.2427276029652166, 32'sd-0.36812410706610166, 32'sd-0.12146048428110535, 32'sd0.13242570701146394, 32'sd-0.005634926113273284, 32'sd0.06395754252460062, 32'sd-0.07921672851878307, 32'sd0.007518979897660356, 32'sd0.012508501006588017, 32'sd0.021509213769028722, 32'sd0.10137193921490308, 32'sd0.0550060055865133, 32'sd0.010364515908606393, 32'sd0.13752147741644027, 32'sd0.09138643073366884, 32'sd0.058893022838489774, 32'sd0.02871400290181819, 32'sd0.022726812381680214, 32'sd0.03760477415842812, 32'sd0.012025408590123503, 32'sd0.0838180094154091, 32'sd0.12610815050705357, 32'sd0.15065461472681185, 32'sd0.24631376792601642, 32'sd0.13000598410326025, 32'sd0.25844888084902484, 32'sd0.11038124128117971, 32'sd-0.20298764617168788, 32'sd-0.2941105186795784, 32'sd-0.35686368473908353, 32'sd-0.07437372574627801, 32'sd-0.012805063533355443, 32'sd-0.02574449452133897, 32'sd0.015013225507344468, 32'sd-0.019145381421942286, 32'sd0.03948113478221664, 32'sd0.11178497761031411, 32'sd0.0714520427762624, 32'sd0.13979174932698607, 32'sd0.016544282886638076, 32'sd0.05979014269661751, 32'sd0.11661035802825741, 32'sd-0.10733318753485012, 32'sd0.02316679029778629, 32'sd0.08313099477991302, 32'sd0.08398084590429414, 32'sd0.036129910019058104, 32'sd0.027201936974810968, 32'sd0.12155313912005278, 32'sd0.11865592771782368, 32'sd0.1749682483776781, 32'sd0.09635519487887165, 32'sd0.21440892102099068, 32'sd0.15641252077866055, 32'sd0.0020536763530991705, 32'sd-0.08176756051460853, 32'sd-0.2698624382869181, 32'sd-0.1948003866708614, 32'sd-0.12407042403848736, 32'sd0.03596974033806083, 32'sd-0.033572666868248, 32'sd0.04090571517403072, 32'sd-0.0821271316862217, 32'sd0.00690980782979179, 32'sd0.02024499930636799, 32'sd0.0889630488515173, 32'sd0.07318058192856677, 32'sd-0.002456404224195525, 32'sd0.051578964683603616, 32'sd-0.04516403933264609, 32'sd0.018189532005908667, 32'sd0.08643697128941297, 32'sd-0.05490528880460223, 32'sd0.02824062795836869, 32'sd-0.06317263773256444, 32'sd-0.09878643877725288, 32'sd0.033269602573623554, 32'sd0.10293057101770033, 32'sd0.11307954710296582, 32'sd0.02742177352506899, 32'sd0.1257836516286322, 32'sd-0.050733887413185026, 32'sd-0.14202247780892374, 32'sd-0.2471538518508078, 32'sd-0.2659967515448463, 32'sd-0.22006958642072563, 32'sd-0.12715115039059513, 32'sd-0.11439374389566999, 32'sd-0.16322704496529705, 32'sd-0.06462884975655843, 32'sd0.021735736771498072, 32'sd-0.024242661253378622, 32'sd0.030750219493405357, 32'sd0.05246183579819695, 32'sd0.059404231664598184, 32'sd-0.08242942729025166, 32'sd0.08207075187882072, 32'sd-0.006879797633230326, 32'sd0.027291418017896925, 32'sd0.031204663178240152, 32'sd0.0429819169103119, 32'sd0.013654511567387779, 32'sd0.04715114643279134, 32'sd-0.02336259065509511, 32'sd-0.012755808783930157, 32'sd0.14183059361909844, 32'sd0.1062291927770183, 32'sd0.1365000207828451, 32'sd-0.0965803273662606, 32'sd-0.10056278203305624, 32'sd-0.2366186870177421, 32'sd-0.3342919053715811, 32'sd-0.2650921748985043, 32'sd-0.1043526729916079, 32'sd0.022073918150443485, 32'sd-0.13548781553113623, 32'sd-0.09172397938798613, 32'sd-0.04471707656647152, 32'sd-0.0328130409852944, 32'sd0.053611745867745524, 32'sd0.09161454498045947, 32'sd0.06227355873118946, 32'sd-0.077848167282392, 32'sd-0.06015766688448124, 32'sd0.14121615937931817, 32'sd-0.008313220877917263, 32'sd0.04281120032275044, 32'sd-4.7717526423602434e-117, 32'sd-0.04000759277307284, 32'sd0.06400011289633496, 32'sd0.06851150475806221, 32'sd0.12188122911450956, 32'sd0.10273410022711693, 32'sd0.06965319164437181, 32'sd0.04611811561485771, 32'sd0.004217123863249606, 32'sd0.0470210131023259, 32'sd-0.1725693082804886, 32'sd-0.2554181739647573, 32'sd-0.21797253821387214, 32'sd-0.16952396317969207, 32'sd-0.03719972195133521, 32'sd-0.04793587717902216, 32'sd0.0619248108780512, 32'sd-0.06938368617876728, 32'sd0.07120500161704905, 32'sd0.07250636649192949, 32'sd0.008541661331514095, 32'sd0.040275111243816684, 32'sd-0.06560580253939517, 32'sd0.005304873664710224, 32'sd0.052839743860067734, 32'sd0.07053246940129625, 32'sd-0.009798195992384918, 32'sd-0.04576278253397565, 32'sd0.042781558128625816, 32'sd-0.0626250482570157, 32'sd0.007018761318813921, 32'sd0.007918133187758952, 32'sd0.02593423173001867, 32'sd-0.008492395976821292, 32'sd-0.011746027182958111, 32'sd0.008706888999813771, 32'sd0.05995148823414959, 32'sd0.03742480329865113, 32'sd0.02755993131769571, 32'sd-0.16823824219264308, 32'sd-0.242874622900466, 32'sd-0.06660056695770689, 32'sd-0.02611959526514168, 32'sd-0.06674937453053786, 32'sd-0.023341904321311214, 32'sd-0.007411531930421753, 32'sd0.09994173704244634, 32'sd0.00906711761072423, 32'sd0.07395624652534372, 32'sd0.005410618702606594, 32'sd-0.025919295708191768, 32'sd-0.06620177915822427, 32'sd0.11288987581822796, 32'sd0.05096031502738434, 32'sd-0.08722417897661566, 32'sd0.044711230298527124, 32'sd0.027199247767132295, 32'sd0.06206158241015797, 32'sd0.02698012007834033, 32'sd0.060239371360588406, 32'sd0.028085000472674693, 32'sd2.5407397833651455e-05, 32'sd-0.007799591199393713, 32'sd-0.010343941426805435, 32'sd-0.026136696195342684, 32'sd0.001474711813037847, 32'sd-0.0007177547995430355, 32'sd-0.15391383524670801, 32'sd-0.026655649006412818, 32'sd0.0011186184615830338, 32'sd0.09815665832320934, 32'sd-0.0689921292106513, 32'sd-0.11774823818908373, 32'sd-0.1296577746393433, 32'sd0.10980767942924582, 32'sd-0.06593965059328782, 32'sd-0.055820361628635906, 32'sd-0.07518745352099396, 32'sd-0.07637767298725835, 32'sd-0.027905716183590914, 32'sd0.06840722553001193, 32'sd0.0018721073561822578, 32'sd-0.07051351973512657, 32'sd-0.012615726192259893, 32'sd-5.123638894626229e-126, 32'sd0.0940560423432582, 32'sd0.018446373543169803, 32'sd0.07332365316798387, 32'sd-0.06156340456075932, 32'sd0.019215331046216234, 32'sd0.0008916004958496987, 32'sd0.07291577995791074, 32'sd-0.017143837546157763, 32'sd-0.0367154947283861, 32'sd0.044583680067901914, 32'sd-0.09926650128901866, 32'sd-0.033875433900247255, 32'sd0.016802704132291228, 32'sd-0.09177537052395386, 32'sd-0.017751551482985704, 32'sd0.027546472362604144, 32'sd0.05295486741576412, 32'sd0.08704065682238556, 32'sd0.06158476556625757, 32'sd-0.00042108550418262406, 32'sd-0.012977208492908175, 32'sd-0.028957459698183696, 32'sd-0.22043532767153326, 32'sd-0.08599267744767666, 32'sd0.01445723226282388, 32'sd0.07616118859586776, 32'sd-0.018022071984561818, 32'sd0.04358691378131359, 32'sd0.07154908283258131, 32'sd0.03235888819465323, 32'sd0.028866034052883568, 32'sd-0.0026942262375948185, 32'sd0.007809273140133296, 32'sd-0.08873885869314484, 32'sd0.03662037765683101, 32'sd0.04429094460011727, 32'sd-0.023034774278645417, 32'sd0.014431002595119664, 32'sd0.12858544676271053, 32'sd0.042093073835006475, 32'sd-0.03378115503883833, 32'sd-0.09677287334712856, 32'sd-0.0336128702652516, 32'sd0.021598656175035084, 32'sd-0.05541568018970016, 32'sd0.0482854795909589, 32'sd-0.008042395670758115, 32'sd-0.06527424924340146, 32'sd-0.0009992222244930003, 32'sd0.030532018487612247, 32'sd-0.08161741502978695, 32'sd0.03768815044780025, 32'sd0.07440965714777988, 32'sd0.038846116839595005, 32'sd0.026076855811417096, 32'sd-0.02062066868168265, 32'sd0.05099339059890768, 32'sd0.05894745156933516, 32'sd-0.08569075131203889, 32'sd0.017710747317709327, 32'sd0.02580358759207205, 32'sd-0.007793684948926728, 32'sd-0.05157868236441297, 32'sd0.06711920545390157, 32'sd-0.05572855900431773, 32'sd0.04537305145091285, 32'sd0.0025719349513926492, 32'sd-0.013402106376791909, 32'sd0.08381356192728112, 32'sd0.0007006079954314161, 32'sd-0.05458144106508454, 32'sd0.00396181818474918, 32'sd0.02560740717975456, 32'sd-0.0685508467797765, 32'sd-0.08945283973072062, 32'sd-0.01947456479717129, 32'sd0.02830014645340859, 32'sd-0.05242611876738471, 32'sd-0.014821745459392771, 32'sd-0.07246081209341602, 32'sd0.10942653927524673, 32'sd0.03671316638599038, 32'sd0.030658206247542154, 32'sd3.761453895050323e-115, 32'sd0.04155189088473439, 32'sd-0.06436011443756735, 32'sd-0.03652717258664788, 32'sd0.07138431288176403, 32'sd0.038149287986730236, 32'sd0.08419690107654006, 32'sd0.012595836382870368, 32'sd0.09909976702591043, 32'sd0.06614337291262701, 32'sd-0.0012766117850721715, 32'sd-0.06546223479024628, 32'sd0.032691596904791266, 32'sd0.03279054005006891, 32'sd0.006778595908027124, 32'sd-0.03039993959477889, 32'sd-0.022306574481220857, 32'sd0.023483204610962028, 32'sd-0.022168939333865878, 32'sd-0.0408421893705582, 32'sd0.06697781020134365, 32'sd0.026896969183550078, 32'sd0.04621985086645423, 32'sd0.026251106977805482, 32'sd0.005284360346199343, 32'sd0.06758443320256582, 32'sd0.03923670896424269, 32'sd-2.9430812475326986e-126, 32'sd-1.6317020931552796e-125, 32'sd-3.1478824771452813e-114, 32'sd0.033960642407572815, 32'sd0.061639963130848296, 32'sd0.0778205889753506, 32'sd0.12902530192978556, 32'sd0.053346005474496, 32'sd-0.03194851562716246, 32'sd0.004019362368006849, 32'sd0.04574573257526248, 32'sd-0.08458773506866747, 32'sd-0.02794914651330018, 32'sd0.07048622374331538, 32'sd-0.033415488968503756, 32'sd-0.07976103927295174, 32'sd0.008130170640631724, 32'sd-0.029883047980178275, 32'sd0.03061688733624397, 32'sd0.009181363501436978, 32'sd-0.055128508690938265, 32'sd-0.07397446696229833, 32'sd0.09035308215918593, 32'sd-0.058958554426916866, 32'sd-0.09903782505655788, 32'sd0.06560491340565608, 32'sd0.060923310020367695, 32'sd0.05827109466464567, 32'sd8.951786111136053e-123, 32'sd1.144308579232308e-124, 32'sd3.6635620296470515e-116, 32'sd-0.02066543663321504, 32'sd0.0004075068897153921, 32'sd0.06903115126883023, 32'sd0.03577067717321428, 32'sd0.05014418264772733, 32'sd-0.06547074530801275, 32'sd0.09787161398051789, 32'sd0.02782671303448666, 32'sd-0.01306034048476258, 32'sd0.04819992625453643, 32'sd0.11382922354561005, 32'sd0.04064415067142385, 32'sd0.018479250089304164, 32'sd-0.007056799447247297, 32'sd0.17858734289687545, 32'sd0.023092408106247707, 32'sd0.020762738035405508, 32'sd-0.10769756393981, 32'sd-0.06681218295699999, 32'sd0.016137361717672796, 32'sd0.04953686095186136, 32'sd0.06946431348229581, 32'sd-0.03520321238996876, 32'sd-0.002967615166082954, 32'sd0.02229717572301041, 32'sd-4.403384947834011e-118, 32'sd4.721139683606998e-117, 32'sd1.0394186298386922e-121, 32'sd2.0244322061944948e-117, 32'sd0.005703106699778489, 32'sd-0.05185098869622929, 32'sd0.08379193977452146, 32'sd0.007973762788553086, 32'sd0.007900002015730432, 32'sd0.06345952630450419, 32'sd-0.05288879291207761, 32'sd-0.07853896699179617, 32'sd-0.044670593935445355, 32'sd0.04925598462410363, 32'sd0.054936295650534775, 32'sd-0.04281264788162321, 32'sd-0.046757904782861036, 32'sd0.03252147054691895, 32'sd0.07240897382853288, 32'sd-0.04011630818521445, 32'sd0.08327940063630157, 32'sd0.09378596250875909, 32'sd-0.007027415544991831, 32'sd0.050635597806338875, 32'sd-0.03067716178039857, 32'sd0.11280770351296157, 32'sd0.08845059210706208, 32'sd-5.187442048642249e-130, 32'sd-2.566329021532114e-126, 32'sd1.2508268123086093e-117, 32'sd-7.494424509136232e-115, 32'sd-7.959951264266458e-117, 32'sd-4.3670508976326e-117, 32'sd0.1055109086121086, 32'sd0.055215832448343494, 32'sd-0.0017745827850329033, 32'sd0.037168148379559916, 32'sd-0.011303098637667623, 32'sd0.001712717705105268, 32'sd0.06208556577359966, 32'sd0.04058668841863585, 32'sd0.09166341618500769, 32'sd0.01807058290135168, 32'sd-0.001029207464457414, 32'sd0.0114113668893578, 32'sd0.00022618367459129133, 32'sd0.011141607912210225, 32'sd-0.04822057122649767, 32'sd0.0018546166781968666, 32'sd-0.11505811421358393, 32'sd-0.0326186376643908, 32'sd0.03371685458720627, 32'sd0.039075421044702616, 32'sd1.9730137293607463e-127, 32'sd-3.2884186332430047e-121, 32'sd3.589892060947724e-114, 32'sd-8.495895957915283e-117},
        '{32'sd2.677653543914882e-117, 32'sd-7.106830720264755e-115, 32'sd1.392404007670309e-118, 32'sd-1.072865713636163e-127, 32'sd-5.772179737480629e-121, 32'sd1.7486896134429178e-118, 32'sd-2.2600540744823265e-125, 32'sd-5.58286948397376e-117, 32'sd-9.883945712616118e-116, 32'sd1.0273207504070928e-119, 32'sd-2.968020249133398e-129, 32'sd2.9510874722568516e-116, 32'sd-0.02125775082926843, 32'sd-0.010345416749860168, 32'sd0.027444297477680683, 32'sd-0.047777968427063444, 32'sd-8.383310705960898e-120, 32'sd6.960639632516714e-121, 32'sd-6.828488350054217e-124, 32'sd6.351935782479691e-118, 32'sd-3.4827071406079536e-115, 32'sd-5.065702177410239e-118, 32'sd1.3620889850471176e-118, 32'sd2.962710376272047e-116, 32'sd-3.619832875937276e-127, 32'sd-5.426247241483566e-126, 32'sd8.86410021461497e-127, 32'sd4.71005263718144e-117, 32'sd7.171970700891771e-115, 32'sd-6.522524598729335e-115, 32'sd2.5210641819165007e-115, 32'sd2.7670076781586558e-118, 32'sd-0.04502335897906436, 32'sd0.044763166818725476, 32'sd-0.02696670641142908, 32'sd-0.03821569202052109, 32'sd-0.03958348518263375, 32'sd0.006878081351787716, 32'sd0.03250643425436866, 32'sd-0.009450637636161998, 32'sd0.043818346607386434, 32'sd0.0008660477038229297, 32'sd0.11222314234820663, 32'sd0.00614663809723698, 32'sd-0.024886610983182154, 32'sd0.04981271174734008, 32'sd-0.004106054210809705, 32'sd-0.07483966945002028, 32'sd-0.004814583191509263, 32'sd-0.06701063957364121, 32'sd-0.08092577888313134, 32'sd0.04047701671366375, 32'sd4.8623869608274966e-123, 32'sd-1.4352847577228193e-118, 32'sd-4.5096466997901276e-128, 32'sd1.1038105667751723e-121, 32'sd-1.0032944392842965e-117, 32'sd1.3610527970142764e-124, 32'sd0.006374317819252494, 32'sd-0.03362746273165223, 32'sd0.03443842488058966, 32'sd-0.05505317284685285, 32'sd-0.057190051140039014, 32'sd0.04476632243239486, 32'sd0.0336721910541971, 32'sd-0.01630277169708004, 32'sd0.0664532900269434, 32'sd0.07218990956078343, 32'sd-0.0511721677662933, 32'sd0.06406369252944268, 32'sd0.017580051926387348, 32'sd-0.02732204822502549, 32'sd-0.09109666487663189, 32'sd-0.05143630113678492, 32'sd-0.10069283198608008, 32'sd-0.1113919301970478, 32'sd-0.13099480040391465, 32'sd-0.024350573206599807, 32'sd-0.00965643974504462, 32'sd-0.028294106933958604, 32'sd-0.055062963892533554, 32'sd-0.049892021090098194, 32'sd-8.80336921877868e-121, 32'sd-5.269270095937025e-118, 32'sd-7.268475908541453e-129, 32'sd6.883645344688802e-126, 32'sd0.020910562409119055, 32'sd0.05112176013384408, 32'sd0.02729011990282438, 32'sd-0.08723838037005975, 32'sd-0.04381740307906789, 32'sd-0.09834450535165663, 32'sd-0.009507294781849578, 32'sd0.05802099367063603, 32'sd-0.012922531091171077, 32'sd-0.1942819593276375, 32'sd-0.04728004826977227, 32'sd-0.015095159126711949, 32'sd-0.06675166283936855, 32'sd0.03295213911266334, 32'sd0.06321197835011196, 32'sd0.035602801576198814, 32'sd0.026182408885647372, 32'sd-0.00035873191377764057, 32'sd-0.047415677653298495, 32'sd-0.024882032409263843, 32'sd0.02275654633823438, 32'sd-0.007656820681403227, 32'sd-0.09666804708681168, 32'sd-0.00402429141406401, 32'sd-0.006915826645587335, 32'sd-1.504399950369743e-122, 32'sd3.037669852174705e-122, 32'sd-0.044425975470973524, 32'sd-0.033560802597461054, 32'sd-0.057212854644899405, 32'sd-0.02720661008712111, 32'sd0.012959763571355542, 32'sd0.028305435142509352, 32'sd-0.019166366744246644, 32'sd-0.06502505372871024, 32'sd-0.04295047325664595, 32'sd-0.04502020089869754, 32'sd0.012173223330083234, 32'sd0.06259756170543257, 32'sd0.04888700095213144, 32'sd0.11479791123771062, 32'sd-0.00974297248303704, 32'sd0.05459440745259733, 32'sd0.006134822838387269, 32'sd0.11130164674174188, 32'sd0.11421116900378393, 32'sd0.09503569612563482, 32'sd-0.05685706730758359, 32'sd-0.024997678477989355, 32'sd-0.02721777257990325, 32'sd-0.06659360964412908, 32'sd-0.077724454990781, 32'sd-0.00516327042459411, 32'sd0.02146584208259211, 32'sd9.816333323363095e-126, 32'sd0.003895797525750016, 32'sd0.010848542674800923, 32'sd-0.07461605920062551, 32'sd-0.05561917825784803, 32'sd0.09420970693436474, 32'sd0.05318582333781523, 32'sd-0.1393819574211861, 32'sd-0.043517065361679506, 32'sd0.041739480298773786, 32'sd-0.029359284455753767, 32'sd0.10866570184377469, 32'sd0.01702691862675643, 32'sd0.057003328459494434, 32'sd0.10861360625042553, 32'sd0.07240064499355849, 32'sd0.03811281354488013, 32'sd0.12722553373878834, 32'sd0.06624285223502362, 32'sd-0.04656544504892906, 32'sd0.07765312777464571, 32'sd0.029051386603869602, 32'sd0.01868972219072041, 32'sd-0.030389880357482642, 32'sd-0.08941882875017004, 32'sd0.0769361154069468, 32'sd0.1043378132459285, 32'sd-0.002216352678920894, 32'sd9.431806316846874e-124, 32'sd-0.002404095049793946, 32'sd-0.04076161960307996, 32'sd0.05309970174247419, 32'sd0.032533640136288226, 32'sd-0.07114190978735951, 32'sd-0.03864115910220961, 32'sd0.02093892095638864, 32'sd-0.07987540453385643, 32'sd-0.03077464509354489, 32'sd0.012317220985127381, 32'sd0.11062769583522637, 32'sd0.10308938012179249, 32'sd0.020043231062131683, 32'sd-0.056596346436960605, 32'sd0.08492724639214776, 32'sd0.14822939133418875, 32'sd0.19897149211615517, 32'sd0.039473279029624636, 32'sd0.14303202283659974, 32'sd0.052887791484155344, 32'sd0.06962871830086116, 32'sd0.045342168239567306, 32'sd0.026314022323855796, 32'sd-0.06727069771536448, 32'sd-0.05388399074067304, 32'sd-0.0246006787269883, 32'sd-0.027452452478287138, 32'sd-0.02017317742593204, 32'sd-0.0002662018181097276, 32'sd0.040800166851127265, 32'sd-0.004516523033398455, 32'sd0.02600179752828097, 32'sd-0.021769123175206618, 32'sd-0.04322390600794488, 32'sd-0.07976908847590315, 32'sd-0.17467512037947755, 32'sd-0.04385709589063767, 32'sd0.07388754816403309, 32'sd0.04818493416913989, 32'sd0.021206623784623353, 32'sd-0.013250535175545891, 32'sd-0.06415035861783533, 32'sd-0.026935993111554587, 32'sd0.01659657415516142, 32'sd0.08659105707036263, 32'sd0.08465681407551737, 32'sd0.06610641109346407, 32'sd0.08215216811362598, 32'sd0.09449234905712461, 32'sd-0.016757764893779614, 32'sd0.02955800244818472, 32'sd-0.04407300614887237, 32'sd0.025343973376192288, 32'sd-0.02917146957491494, 32'sd-0.025725207573385866, 32'sd0.04010297993314046, 32'sd-0.026006889617028756, 32'sd0.07261647215826797, 32'sd-0.041745252605817275, 32'sd-0.03382290808586418, 32'sd-0.07314834718874386, 32'sd-0.0694910506984923, 32'sd-0.02011425542070566, 32'sd0.03503955078007301, 32'sd0.12017505352867221, 32'sd0.08342362857835338, 32'sd0.06098039964813702, 32'sd0.0022887947841581944, 32'sd-0.003399750672467412, 32'sd-0.005110737278646408, 32'sd0.014119002693946336, 32'sd0.013164111161576968, 32'sd0.07691289125405969, 32'sd0.08797459792621208, 32'sd0.13197280880713425, 32'sd0.13398506568523724, 32'sd-0.0008199771460617369, 32'sd0.004187853958048746, 32'sd0.07555873485853379, 32'sd-0.03926296583986669, 32'sd-0.030166667947295594, 32'sd-0.08573973462091405, 32'sd0.04388083545901003, 32'sd-0.020724614676508508, 32'sd-0.048087984096148804, 32'sd0.09874894675476528, 32'sd0.15681819046131298, 32'sd0.0279651845417946, 32'sd0.10016827090026079, 32'sd0.12788330344242174, 32'sd0.06114052481283846, 32'sd0.13654630158977465, 32'sd0.11661690334780765, 32'sd0.06791143685585414, 32'sd-0.13677251701654455, 32'sd-0.1860833077191057, 32'sd-0.10620392085834113, 32'sd-0.09548293732995174, 32'sd-0.021963671562055864, 32'sd0.013744234308382956, 32'sd-0.11269599178094948, 32'sd0.0740693077155197, 32'sd0.04515639756120965, 32'sd0.0539561145539013, 32'sd-0.004381394550397832, 32'sd-0.0013320913373747625, 32'sd-0.004043282516541838, 32'sd0.0538617305627749, 32'sd0.009995370485576116, 32'sd0.03126542024118634, 32'sd-0.03129039040859777, 32'sd-0.05136927528354561, 32'sd0.04085284808746502, 32'sd0.07507821702806738, 32'sd0.07192701563395677, 32'sd0.0671079404908888, 32'sd0.18064166795337733, 32'sd-0.005533163443330728, 32'sd0.14081748820009557, 32'sd0.1356381471463155, 32'sd-0.03475714010432818, 32'sd-0.02497698350662839, 32'sd-0.0639652169420526, 32'sd-0.0752533027215322, 32'sd-0.17355157459997966, 32'sd-0.0737801852359139, 32'sd0.035754784151510455, 32'sd-0.04415030423514028, 32'sd0.02468130723624238, 32'sd0.09956372193211957, 32'sd-0.05027515658684082, 32'sd0.036908937798335595, 32'sd-0.008311302239971372, 32'sd0.11315219585481802, 32'sd0.07267691008177289, 32'sd-0.01697672443327572, 32'sd0.04610417260282117, 32'sd0.04083181966877348, 32'sd0.04741315634693297, 32'sd0.004053946159212988, 32'sd-0.0976682128339102, 32'sd-9.202104897578941e-05, 32'sd0.09187056732251363, 32'sd-0.05776179096852086, 32'sd0.08912124156376973, 32'sd0.05277068098330651, 32'sd0.12437729126529705, 32'sd0.015815505490429226, 32'sd-0.004567962714263179, 32'sd-0.01317234620555647, 32'sd0.08939701464078148, 32'sd0.03926133658235902, 32'sd0.04353826368554149, 32'sd-0.1294648185023904, 32'sd-0.09279323266202352, 32'sd-0.0432723815621702, 32'sd-0.11638374156813887, 32'sd-0.14771819095574923, 32'sd0.0024435133449906576, 32'sd0.062220630322352734, 32'sd0.1547329172286158, 32'sd0.13501606185854445, 32'sd0.1278852129667534, 32'sd-0.023006309627147947, 32'sd-0.021337199528627976, 32'sd0.013032516688715318, 32'sd0.10176676445999999, 32'sd-0.0004795365514590602, 32'sd-0.04814293826186458, 32'sd-0.02289468087672801, 32'sd0.11189415128137503, 32'sd-0.08507268767798949, 32'sd-0.04833711729703912, 32'sd0.14243143934469418, 32'sd0.07215002476249752, 32'sd-0.09927021536778032, 32'sd0.0106727810864549, 32'sd0.06582835847896877, 32'sd0.11261286009817863, 32'sd0.07117066940177827, 32'sd-0.10510782415531528, 32'sd-0.11858858909044435, 32'sd-0.19356839034094808, 32'sd-0.14864145483468663, 32'sd0.011885736638938157, 32'sd-0.12078805441327976, 32'sd-0.04296061076090002, 32'sd0.1294624466845361, 32'sd0.054531398631483846, 32'sd0.09374805523700534, 32'sd0.08131279046842693, 32'sd0.02797924651579577, 32'sd0.02767040027721525, 32'sd-0.08715939999362465, 32'sd0.07019167299742769, 32'sd0.02342296612552738, 32'sd0.00714363137149837, 32'sd0.03162041148767968, 32'sd0.13495918529006048, 32'sd-0.03544747874882038, 32'sd-0.04192352004648119, 32'sd0.020348792613582755, 32'sd-0.09585745080564231, 32'sd0.05310792518818399, 32'sd-0.01527557637196926, 32'sd-0.03237512059761369, 32'sd-0.008773638325657494, 32'sd-0.05287164731786346, 32'sd0.0127222417178282, 32'sd-0.055937505160215104, 32'sd-0.05014309651112468, 32'sd0.017494443132886252, 32'sd-0.0686599711802871, 32'sd-0.07632397761611255, 32'sd0.025074921869735728, 32'sd0.10616941807871445, 32'sd0.18803395903008968, 32'sd0.08240928831512812, 32'sd0.009758443090307859, 32'sd-0.11217783042547018, 32'sd-0.07723161467751709, 32'sd-0.09386483025235227, 32'sd0.09086656699979787, 32'sd0.012362947768190696, 32'sd-0.012407573406707858, 32'sd-0.09366377398700881, 32'sd-0.04257370573423977, 32'sd0.08477516649398403, 32'sd-0.0035198843225579283, 32'sd-0.08878160862561903, 32'sd0.01924364738410836, 32'sd-0.17703601651696899, 32'sd-0.1760756862016698, 32'sd-0.0834790773703291, 32'sd-0.08307802048137958, 32'sd-0.08477826084272347, 32'sd0.09271091526622041, 32'sd-0.0018106858411164192, 32'sd0.05313430678977553, 32'sd0.06190761257054988, 32'sd-0.060353558447422836, 32'sd-0.11113241265542463, 32'sd-0.05443883751010968, 32'sd-0.02442929092598637, 32'sd0.06444796864015408, 32'sd0.004145368884960405, 32'sd-0.0569345648949319, 32'sd-0.13505682834158336, 32'sd0.077028552526491, 32'sd0.13370401232630338, 32'sd-0.002763697432208023, 32'sd-0.00988217619665145, 32'sd-0.03780184301933216, 32'sd-0.016421407872611964, 32'sd0.06556619052709596, 32'sd0.008764077805262829, 32'sd0.0145465227753156, 32'sd-0.009653084803384714, 32'sd-0.02921480348486217, 32'sd-0.05767780823885639, 32'sd0.0567869908787249, 32'sd-0.03834288877678489, 32'sd0.03318467351831847, 32'sd0.043648141667423826, 32'sd0.030084465363735272, 32'sd-0.062337868552173034, 32'sd-0.01474663782685105, 32'sd-0.03893595532391364, 32'sd-0.086533185551858, 32'sd-0.08899915436527706, 32'sd-0.07313079273856499, 32'sd0.043451924736543836, 32'sd0.09284706001700498, 32'sd0.0049701797151810835, 32'sd-0.14283890543470487, 32'sd-0.014398691859016424, 32'sd-0.12744768924191965, 32'sd0.012195359736614151, 32'sd0.021564798702671, 32'sd0.025997490563315292, 32'sd0.04877942041679047, 32'sd-0.055486172667910116, 32'sd0.10673577599276234, 32'sd0.036747679473520686, 32'sd-0.0890585075374857, 32'sd0.06534751771511653, 32'sd-0.08183173160381475, 32'sd0.0943231246891301, 32'sd-0.01604404114137842, 32'sd0.042750964802310144, 32'sd0.07105477879866694, 32'sd0.16982738851540924, 32'sd0.16011472387715175, 32'sd-0.11258381170518972, 32'sd0.012131160308808642, 32'sd0.03829442349031885, 32'sd-0.10908445547916475, 32'sd-0.09747281833085107, 32'sd0.008491182810713102, 32'sd-0.08469079585484185, 32'sd0.00928080015567, 32'sd-0.032422494014620884, 32'sd-0.014270365061405301, 32'sd0.05486622815999055, 32'sd0.05088404910682659, 32'sd-0.05183941136707481, 32'sd0.001211030869810737, 32'sd-1.2752247190938237e-117, 32'sd0.03609661967645554, 32'sd0.03964409058695229, 32'sd0.09037775330605108, 32'sd0.09595465012467637, 32'sd-0.027504610016208013, 32'sd0.08123975254818099, 32'sd0.007455909853815464, 32'sd0.035240630996753695, 32'sd0.00581653455980726, 32'sd0.061254986815182356, 32'sd0.224446700241921, 32'sd0.1953120869173575, 32'sd0.1400489677049725, 32'sd-0.03656214993182585, 32'sd-0.22317319189584747, 32'sd-0.20229065207173128, 32'sd-0.15568763754706216, 32'sd-0.18229374197144033, 32'sd-0.09525472980937874, 32'sd-0.021213056351024568, 32'sd-0.15607516271025362, 32'sd-0.07822778753253594, 32'sd0.047724441994888143, 32'sd-0.0421429358361518, 32'sd0.033745161603378045, 32'sd0.06739064267085336, 32'sd-0.0008000355400614814, 32'sd-0.04146863557821662, 32'sd0.016352091558051094, 32'sd0.026838663796430084, 32'sd-0.008876669440671132, 32'sd0.015672238306297936, 32'sd-0.01873314404597339, 32'sd0.05577803531275746, 32'sd-0.013294535996622683, 32'sd0.008174290217038164, 32'sd0.12278272007363443, 32'sd0.12985405232107766, 32'sd0.24574012934277115, 32'sd0.10492518334667382, 32'sd-0.057328178764897444, 32'sd-0.20251321182584658, 32'sd-0.3244273134780105, 32'sd-0.1986609434763399, 32'sd-0.028140863066996234, 32'sd-0.009443964826403604, 32'sd-0.1765081080636702, 32'sd-0.10315391679250958, 32'sd-0.11385294385694271, 32'sd0.027752141306915955, 32'sd-0.021925773034225087, 32'sd0.08620152300501799, 32'sd-0.048671138358171495, 32'sd0.02548613565744002, 32'sd-0.06750093913939208, 32'sd-0.0401481631421949, 32'sd-0.03389662160808467, 32'sd-0.04268570074605433, 32'sd-0.09551353466963522, 32'sd0.040165114488152916, 32'sd-0.10468287484140636, 32'sd0.02707550072887815, 32'sd-0.003084120017552625, 32'sd0.05255432820961623, 32'sd0.12828705709334484, 32'sd0.17037324087117295, 32'sd0.16874091334463184, 32'sd0.07701724770373596, 32'sd0.04876631926545816, 32'sd-0.29896491302512396, 32'sd-0.20456287430832762, 32'sd-0.0593068393421341, 32'sd0.03326012035126563, 32'sd-0.08223682070643451, 32'sd-0.1735384831627573, 32'sd-0.0367432603774685, 32'sd-0.038227841332396144, 32'sd0.043868449746982605, 32'sd0.0699659941233161, 32'sd0.007729023391518486, 32'sd0.007548641858489323, 32'sd0.011725576882703759, 32'sd0.009165068572990303, 32'sd4.900789953429212e-118, 32'sd-0.08356717015721908, 32'sd0.10116784706275785, 32'sd0.08237168508824387, 32'sd0.016235350559166948, 32'sd-0.0015849035915292498, 32'sd0.08309395561820641, 32'sd0.11802078434376902, 32'sd0.23211195728306713, 32'sd0.14535027780706672, 32'sd0.13281484931432852, 32'sd0.16706855728141692, 32'sd0.05847576947623681, 32'sd-0.07473420667667051, 32'sd-0.3318813779491382, 32'sd-0.05225504416970567, 32'sd0.05308792629097195, 32'sd0.028684047443906926, 32'sd0.03324091641966281, 32'sd0.01240150582386189, 32'sd-0.07053643301464188, 32'sd0.0319448691544346, 32'sd-0.09788515529855737, 32'sd0.001697507489794053, 32'sd0.0982405227108206, 32'sd0.053040728786189595, 32'sd0.05951143242884155, 32'sd0.052785504326477786, 32'sd-0.042494768063330024, 32'sd-0.04341430393700797, 32'sd0.031426434828069755, 32'sd-0.0013368257932802594, 32'sd0.04166032170138922, 32'sd0.04660114412301566, 32'sd0.09076808699254238, 32'sd0.04436366116045805, 32'sd0.05834301713500153, 32'sd0.12245408358399688, 32'sd0.13007392866530612, 32'sd0.08168240202393989, 32'sd-0.02197810384700588, 32'sd-0.2551569714405116, 32'sd-0.1524807091222531, 32'sd-0.0701901402716346, 32'sd0.03466134088794607, 32'sd0.0983629779947664, 32'sd0.036758121900164566, 32'sd-0.013596970329658183, 32'sd-0.043088285820359944, 32'sd0.06319913943317712, 32'sd-0.010350988317564062, 32'sd-0.12781427899398806, 32'sd0.036735551828882294, 32'sd0.014552372916266028, 32'sd0.09720221525383439, 32'sd-0.006990953541602664, 32'sd-0.02912599727799919, 32'sd0.022995874966789998, 32'sd-0.03499444633358109, 32'sd-0.08604571357175217, 32'sd-0.0350100141859959, 32'sd0.04362559866133532, 32'sd0.15184620898419451, 32'sd0.09084934887186441, 32'sd0.09007312976515008, 32'sd0.14329061271040547, 32'sd0.12646136695199664, 32'sd-0.046768562091176386, 32'sd-0.09224926874145431, 32'sd-0.1616197234554513, 32'sd-0.04719867664394454, 32'sd-0.028972178905752495, 32'sd-0.11324430733526729, 32'sd0.08611012690994704, 32'sd0.1261476450495391, 32'sd0.019625391035763776, 32'sd0.1142677244446694, 32'sd0.0038970491361109984, 32'sd0.03476469192823061, 32'sd-0.13515189124720442, 32'sd-0.09770481418069994, 32'sd-0.003923302687368484, 32'sd0.04942955850377278, 32'sd0.08729264644787578, 32'sd-4.482593594306065e-122, 32'sd-0.012840338721857145, 32'sd-0.07359352877984378, 32'sd-0.13331555925208258, 32'sd-0.004959886076677798, 32'sd0.018421399986210178, 32'sd0.042463694652497025, 32'sd0.11433933316206356, 32'sd0.14386299218410345, 32'sd0.11731851813315766, 32'sd0.04186752151878695, 32'sd0.06525854198986568, 32'sd-0.045047501003869124, 32'sd-0.05421150677860571, 32'sd-0.08985874066409696, 32'sd-0.06421335518057297, 32'sd-0.0830740562537646, 32'sd-0.09377671926879338, 32'sd-0.028081490992097932, 32'sd0.079878876566854, 32'sd-0.07925171924951926, 32'sd-0.016812483026094144, 32'sd0.014374017388095194, 32'sd-0.11276704573110125, 32'sd-0.0437103238103661, 32'sd-0.00861171695268284, 32'sd0.02356073125014668, 32'sd1.372374769019601e-126, 32'sd1.614684051538121e-125, 32'sd-3.793319031954516e-125, 32'sd-0.02233265382638865, 32'sd-0.04460065028733808, 32'sd-0.047779247830081376, 32'sd0.03666624879729414, 32'sd0.01667118181611972, 32'sd0.07697987538206794, 32'sd0.10495792052373981, 32'sd0.05948842665444706, 32'sd0.06528039908185311, 32'sd0.04985069826460005, 32'sd0.14238249415333615, 32'sd0.03844206300813365, 32'sd-0.03752585218392634, 32'sd-0.13522905062320065, 32'sd-0.21221050317641238, 32'sd-0.11462348327853425, 32'sd0.0343597023611912, 32'sd0.10000622762032926, 32'sd-0.03939107594728145, 32'sd0.015307862065737109, 32'sd0.0421166380221678, 32'sd-0.03794706028807291, 32'sd0.012955396954165255, 32'sd0.10178805585235266, 32'sd-0.029407041221482653, 32'sd-9.569261780907407e-120, 32'sd-6.081228565252419e-121, 32'sd-7.542847729639115e-115, 32'sd-0.007349772237802711, 32'sd0.025195997225468707, 32'sd0.01077944268909253, 32'sd-0.03632955563991611, 32'sd0.05523406011715153, 32'sd0.06874242067886298, 32'sd0.03813169558674135, 32'sd0.16412803929345388, 32'sd0.06119994869568024, 32'sd-0.0823526777521528, 32'sd0.0072435043287075425, 32'sd-0.029328797529177997, 32'sd0.035352509533140224, 32'sd-0.13704791686586146, 32'sd-0.18290456572152522, 32'sd-0.11511840094599778, 32'sd-0.056003796188391575, 32'sd0.021823721075331967, 32'sd0.011633881224025902, 32'sd0.09469520257583292, 32'sd-0.012447662724234908, 32'sd0.0666603542461356, 32'sd0.04354646383586884, 32'sd-0.06418452004605016, 32'sd0.05393139895216502, 32'sd6.385270904701481e-121, 32'sd3.287839393304288e-123, 32'sd6.836531927596138e-125, 32'sd5.07165230634313e-115, 32'sd-0.03335974954018959, 32'sd0.07756410319414796, 32'sd0.0545236054556541, 32'sd0.022022666622831207, 32'sd0.035125427876109706, 32'sd0.03854796218084564, 32'sd-0.02488692092632419, 32'sd-0.012913472263388778, 32'sd-0.1533702245223698, 32'sd-0.06718207387855879, 32'sd0.002399792047491628, 32'sd0.023224785837394082, 32'sd0.00557227501766155, 32'sd-0.05648779593307837, 32'sd-0.001544178079579971, 32'sd0.011159572697690518, 32'sd0.0641400193778383, 32'sd0.05681223865427268, 32'sd0.029810708703691225, 32'sd0.01242715208410419, 32'sd-0.020503923809859836, 32'sd0.009113969198863514, 32'sd-0.045618660387844574, 32'sd-8.708586057075031e-127, 32'sd1.0049812003033534e-121, 32'sd6.134176901493539e-126, 32'sd2.3042871207074873e-121, 32'sd9.901290186162369e-117, 32'sd6.710603718343607e-123, 32'sd0.019887022749645638, 32'sd-0.038136607437021915, 32'sd-0.010273366718984458, 32'sd-0.02857955070031975, 32'sd-0.08172812090435409, 32'sd-0.05349528192431158, 32'sd0.026336083647773078, 32'sd-0.030476929853723682, 32'sd0.04392545929286649, 32'sd0.0050351374445767915, 32'sd0.06670669615166785, 32'sd-0.033347442007310796, 32'sd0.02795669635012317, 32'sd-0.07896352394369847, 32'sd-0.04153112850153259, 32'sd0.031593423245296945, 32'sd-0.08570532019259207, 32'sd0.016664290251543867, 32'sd0.0756062130411495, 32'sd0.08047179335815065, 32'sd-1.3993807134924713e-118, 32'sd-7.25380180187684e-124, 32'sd2.4617042044674487e-124, 32'sd-1.2241402939738204e-128},
        '{32'sd-8.638063425991461e-120, 32'sd-3.2615058974203325e-120, 32'sd-1.7712603994863375e-121, 32'sd1.6639525260084647e-121, 32'sd2.07259769893924e-126, 32'sd2.1709806359799463e-120, 32'sd-4.820840882507423e-124, 32'sd1.5701050637280052e-115, 32'sd5.636691143346806e-116, 32'sd-8.700790856583702e-125, 32'sd-2.909339509231377e-122, 32'sd-8.198349027812175e-120, 32'sd-0.020377205019892763, 32'sd-0.012188267275277479, 32'sd0.07721888447447058, 32'sd0.1112525029225015, 32'sd1.1092674908098544e-121, 32'sd3.065891822747712e-126, 32'sd-1.7003777236593638e-126, 32'sd-6.135124542095124e-119, 32'sd-1.9623272558414375e-117, 32'sd-3.646356829561973e-122, 32'sd-1.0471566961676454e-119, 32'sd-7.31975682562529e-125, 32'sd-7.100587333189956e-122, 32'sd-7.313971588203575e-127, 32'sd8.404679306652828e-120, 32'sd-1.1780326331407113e-118, 32'sd1.513170092461186e-123, 32'sd1.559000881630326e-125, 32'sd2.76662687157994e-123, 32'sd6.83473904677963e-117, 32'sd-0.06969878383597221, 32'sd0.013519127647470056, 32'sd0.0938797889833528, 32'sd0.0014411921845697228, 32'sd0.02225445986956376, 32'sd-0.023605982497494, 32'sd-0.02784531128683476, 32'sd0.10900149623714521, 32'sd0.05739495369279635, 32'sd0.0569590437808324, 32'sd-0.10322838588950978, 32'sd-0.01129313180048012, 32'sd0.07831488894073611, 32'sd-0.021000660577636953, 32'sd-0.08303888376244993, 32'sd-0.05008011591420132, 32'sd-0.04266626397150908, 32'sd-0.03036477975748671, 32'sd0.009025428901228765, 32'sd-0.005741415431800175, 32'sd-6.473816643875967e-126, 32'sd-6.210902442759774e-120, 32'sd9.012455840269903e-122, 32'sd9.333943821434854e-128, 32'sd1.0267566365604049e-123, 32'sd-3.788821093277954e-122, 32'sd0.00733647793790713, 32'sd-0.015960784326811514, 32'sd0.0025380841495552466, 32'sd0.10786945240151606, 32'sd-0.023785619730808734, 32'sd0.0013894590212263868, 32'sd0.006502910786033232, 32'sd-0.03134033107141097, 32'sd0.027679578150439817, 32'sd0.14858821793022553, 32'sd0.08664446733068609, 32'sd0.027073334750364702, 32'sd-0.012120933421113712, 32'sd-0.11224598740197786, 32'sd-0.024399507918448797, 32'sd-0.013325183834981118, 32'sd-0.06373212626803289, 32'sd-0.10953580723458482, 32'sd-0.1498387438399862, 32'sd-0.09295428318645699, 32'sd-0.010234142504197801, 32'sd-0.024797206387825486, 32'sd-0.040966828628275304, 32'sd0.016114847883365736, 32'sd9.627562483399069e-116, 32'sd-1.897693861849228e-123, 32'sd-1.943418922312561e-116, 32'sd2.54091823496951e-115, 32'sd0.04742401359030107, 32'sd0.06492782553807681, 32'sd-0.03400202903294061, 32'sd0.045514720732418114, 32'sd0.008212282689774288, 32'sd-0.024876014505083373, 32'sd0.13399601480860887, 32'sd0.1137120164599676, 32'sd0.027662680386745298, 32'sd0.12426162966130519, 32'sd0.1745950165383245, 32'sd-0.059757507241804377, 32'sd0.05164669323290414, 32'sd0.07790376357911244, 32'sd-0.027578668840273917, 32'sd0.02751979478501341, 32'sd0.07378099280207964, 32'sd-0.041372680978940035, 32'sd0.08014647086146155, 32'sd-0.07597725294194803, 32'sd-0.06504641903621904, 32'sd-0.11597882546047933, 32'sd0.026317438617727743, 32'sd0.027041100331960354, 32'sd-0.020202399100635572, 32'sd-1.3041116267039224e-122, 32'sd3.149246210216937e-123, 32'sd-0.02248323977864846, 32'sd0.050282332038024256, 32'sd-0.035520245834386614, 32'sd0.034495515842542075, 32'sd0.01751422913631555, 32'sd0.0674819334758894, 32'sd0.06826221103582213, 32'sd0.055830975842735206, 32'sd0.06240922990059711, 32'sd0.020547083733618108, 32'sd0.1438452132451908, 32'sd0.11738628287565521, 32'sd0.04467414193248404, 32'sd0.005538713511477656, 32'sd0.07695829491648487, 32'sd-0.0345211108859064, 32'sd0.04807670734108325, 32'sd0.08502791376959903, 32'sd0.06457869410620275, 32'sd0.03505125354635993, 32'sd-0.10637807649813404, 32'sd-0.09244859060724586, 32'sd-0.0916370519250398, 32'sd-0.07604632722282537, 32'sd-0.045385870931301815, 32'sd-0.06352086337828776, 32'sd-0.03189010922468693, 32'sd1.2677136761453926e-122, 32'sd-0.052109674891829966, 32'sd0.05193962629880848, 32'sd0.08519082790538096, 32'sd0.09407705308200962, 32'sd-0.02073910955485332, 32'sd-0.0339092964016057, 32'sd-0.048587168985313775, 32'sd0.044442110484565325, 32'sd0.006828163959159184, 32'sd0.04640677334154882, 32'sd-0.16563351909361387, 32'sd-0.18770521564246742, 32'sd-0.03247217532449396, 32'sd-0.0012781241699545325, 32'sd0.07607551295365647, 32'sd-0.05369204401759212, 32'sd-0.0961521722395746, 32'sd-0.025636157151803566, 32'sd0.12153121289256466, 32'sd0.0796847873091086, 32'sd-0.025818106847131102, 32'sd0.11174385704731657, 32'sd0.17847104222795943, 32'sd-0.06870626072638841, 32'sd-0.1362576290305391, 32'sd0.016112503784284686, 32'sd0.02276877660660233, 32'sd-9.72512499030956e-116, 32'sd0.007721873972637195, 32'sd0.04090093555828735, 32'sd0.010438907393399578, 32'sd0.037345176223123486, 32'sd0.028855780330386972, 32'sd0.09331556578425117, 32'sd0.0872143114321919, 32'sd0.028996903349205256, 32'sd0.0717692473415891, 32'sd-0.003154947640284619, 32'sd-0.07360349032565715, 32'sd-0.030626678366460165, 32'sd0.0274917705272677, 32'sd0.05331672305664033, 32'sd-0.05666426077192909, 32'sd-0.060870677001776105, 32'sd-0.12627320668208938, 32'sd-0.04828406228587273, 32'sd-0.09319480020871265, 32'sd0.002775785346323522, 32'sd-0.053725440908285446, 32'sd0.10307737980274505, 32'sd0.14088130685548492, 32'sd-0.00499893790652617, 32'sd0.07568425466142285, 32'sd0.01606003556588265, 32'sd-0.09812420908137058, 32'sd-0.01039713793093785, 32'sd-0.021984921948475615, 32'sd-0.1593173949060306, 32'sd-0.05736344013769908, 32'sd0.06475773848893328, 32'sd0.09417546763222043, 32'sd0.19806562493692764, 32'sd0.14476251094089584, 32'sd0.01637086282041448, 32'sd-0.13998831179260693, 32'sd-0.02645495083618095, 32'sd0.031998375357511676, 32'sd0.05710163080978846, 32'sd-0.014324567592572337, 32'sd-0.030545711387656604, 32'sd-0.025843087355718802, 32'sd-0.06431672690540877, 32'sd-0.029066969460393777, 32'sd-0.0941957118155171, 32'sd-0.02146238208787834, 32'sd-0.051286900386335245, 32'sd0.02559571753684572, 32'sd0.026617923078395906, 32'sd2.489644023407656e-05, 32'sd0.016569649113898643, 32'sd-0.035351151189523033, 32'sd0.11946106307999144, 32'sd0.0015590606648214075, 32'sd-0.01442427097005955, 32'sd-0.01923070596428472, 32'sd-0.05211174837857072, 32'sd-0.16262961550514396, 32'sd-0.04787805679918918, 32'sd0.06463917251484184, 32'sd-0.05258388388626802, 32'sd-0.18982921111803927, 32'sd-0.13298036045285083, 32'sd-0.3222594711104183, 32'sd-0.08030724160605736, 32'sd0.0063890335176915985, 32'sd-0.062379397643625725, 32'sd-0.14440872797074245, 32'sd-0.06903795115528705, 32'sd-0.0730047578390955, 32'sd-0.008456950313958343, 32'sd0.03631022955784138, 32'sd0.09957451371599985, 32'sd0.059905889524177164, 32'sd0.018283109325889963, 32'sd0.06009071034798402, 32'sd0.026731470723876213, 32'sd0.06122671609754394, 32'sd-0.061666389313245, 32'sd0.050907802140422495, 32'sd0.11132387726160473, 32'sd-0.0829227420134132, 32'sd0.00437583032389586, 32'sd-0.09265464831716762, 32'sd0.043103735051362176, 32'sd0.05997601950086449, 32'sd-0.024166738369047393, 32'sd0.010235120767965416, 32'sd-0.20269222601409745, 32'sd-0.38047515576266816, 32'sd-0.25277677852868646, 32'sd-0.2541422805470284, 32'sd-0.14495804470289103, 32'sd0.012808637011773845, 32'sd0.024611359731920225, 32'sd-0.06019467133788619, 32'sd-0.10116424884330906, 32'sd-0.09401195998029424, 32'sd0.034273061783279414, 32'sd0.04883508912888814, 32'sd0.16596928925070029, 32'sd0.12203247736843754, 32'sd0.03664333223013194, 32'sd-0.016797482679026577, 32'sd-0.011797462937099356, 32'sd-0.020671067425970756, 32'sd0.01707737572832115, 32'sd-0.11230583224417429, 32'sd0.07743136840451409, 32'sd0.022039780786824805, 32'sd-0.010730492558548438, 32'sd-0.009225823299491835, 32'sd0.018630382198928888, 32'sd0.11658745169993902, 32'sd-0.07430717621400804, 32'sd-0.15141102901365605, 32'sd-0.10762379166256907, 32'sd-0.18840864460157208, 32'sd-0.19862397828378753, 32'sd0.0012736711569690435, 32'sd-0.03343402168315842, 32'sd-0.06264528276944817, 32'sd0.06863337797814373, 32'sd0.07647627808518541, 32'sd-0.12994403097098153, 32'sd-0.041343814249006273, 32'sd0.12137866745498659, 32'sd0.019476472608601997, 32'sd0.09930694806698032, 32'sd0.1441369730308138, 32'sd0.04073108747670337, 32'sd0.09589591323076045, 32'sd-0.05780098472538151, 32'sd0.03249575315668153, 32'sd0.01624503000841288, 32'sd-0.09217385521396614, 32'sd0.10189423515700852, 32'sd-0.02193775078884478, 32'sd-0.08438432356111769, 32'sd-0.05450341224424162, 32'sd-0.018880813984648862, 32'sd-0.08670818733733403, 32'sd0.1080655941423277, 32'sd-0.07269971502040454, 32'sd0.04646765513936568, 32'sd-0.03311266450216869, 32'sd-0.05830513588284302, 32'sd-0.031721114555875854, 32'sd-0.018875993191678295, 32'sd-0.004269084551311903, 32'sd0.10942445495652171, 32'sd0.026823526598192864, 32'sd-0.036623738621598415, 32'sd0.03578047044551034, 32'sd0.022510048733082287, 32'sd0.05778339428786853, 32'sd0.022175141048711638, 32'sd0.06181082400764083, 32'sd-0.03418392383967695, 32'sd-0.07819661711777516, 32'sd-0.11430279667425623, 32'sd-0.04226169643445264, 32'sd-0.09207837104364122, 32'sd-0.11678709503790702, 32'sd-0.10190965878016708, 32'sd-0.009004613048480261, 32'sd0.029010213758270578, 32'sd-0.006056238338821194, 32'sd-0.07050497038671617, 32'sd-0.02030772120923269, 32'sd0.046902806914772104, 32'sd0.034434592314342836, 32'sd0.010347395632978476, 32'sd0.015171473250452327, 32'sd-0.009540698295489246, 32'sd-0.11782092797883133, 32'sd-0.0776421589962282, 32'sd-0.033580402191834516, 32'sd0.03334780811008348, 32'sd-0.16006333067572956, 32'sd-0.04962519956192608, 32'sd-0.013744381275103143, 32'sd0.04484782881640349, 32'sd-0.005695727510126101, 32'sd0.039408673304631874, 32'sd0.029176594695917855, 32'sd-0.10525922583560648, 32'sd-0.17633272301584438, 32'sd-0.043006565940069824, 32'sd-0.06172162797285699, 32'sd-0.1397452977013714, 32'sd-0.03305025523948027, 32'sd-0.1232497455997751, 32'sd0.08156950413139927, 32'sd0.0367886923294282, 32'sd-0.028047171223547794, 32'sd0.06363449238938067, 32'sd0.11381400488876534, 32'sd0.019269175982458857, 32'sd0.0042333816315721605, 32'sd0.007163955358882567, 32'sd0.006393330017390375, 32'sd-0.041166363054645265, 32'sd0.06353755712997747, 32'sd-0.001994290593115773, 32'sd-0.09466299390597926, 32'sd-0.11019495691626818, 32'sd-0.09013315350289854, 32'sd0.09518588121047099, 32'sd-0.07035577086034647, 32'sd0.10474736972836145, 32'sd0.082419980562887, 32'sd-0.016852665245758864, 32'sd0.05127377468221722, 32'sd0.020251691069054747, 32'sd0.027935867976287523, 32'sd-0.08549881204990568, 32'sd-0.0029952367526955197, 32'sd-0.054913238618824765, 32'sd-0.029874775948342244, 32'sd-0.05208023431607416, 32'sd-0.01170198925069019, 32'sd0.01303397688639869, 32'sd-0.02037303430954721, 32'sd-0.006630338006390426, 32'sd-0.01007140945134376, 32'sd-0.0025050325130047445, 32'sd0.002918744989181536, 32'sd-0.010146552917323592, 32'sd-0.11756162051853322, 32'sd-0.12189878787655899, 32'sd-0.06570936801166997, 32'sd-0.040166233328171354, 32'sd-0.1319697962528201, 32'sd-0.15952416188578653, 32'sd0.02941953085851522, 32'sd0.0563993858586529, 32'sd0.014031428667669554, 32'sd0.04530039086357195, 32'sd-0.022614169063641967, 32'sd0.044808018576560846, 32'sd0.06839945658450575, 32'sd-0.013871024153409055, 32'sd0.06457525477148268, 32'sd-0.11558747315877699, 32'sd0.03549099441456339, 32'sd-0.0883299425107817, 32'sd-0.05103322108620443, 32'sd-0.06787818049611977, 32'sd0.04994896562805603, 32'sd-0.07124942381608355, 32'sd-0.000568535724809227, 32'sd-0.014327713834607061, 32'sd-0.053382815844197254, 32'sd0.0970607825017403, 32'sd-0.03547526818897682, 32'sd-0.049770918983870815, 32'sd-0.16965990574930925, 32'sd-0.07140694127868037, 32'sd-0.22053800804988355, 32'sd-0.11395794724057759, 32'sd-0.13702848199735526, 32'sd0.04775006874376327, 32'sd0.015318716801233045, 32'sd0.061735369390932764, 32'sd0.09916512908251847, 32'sd0.018851347150160656, 32'sd-0.09565566225928726, 32'sd-0.04572671925043229, 32'sd0.07930030622278349, 32'sd0.08763802485847022, 32'sd-0.0756322740847866, 32'sd0.012476574145481109, 32'sd-0.02419118230797329, 32'sd0.002867646173646813, 32'sd-0.01035784760569534, 32'sd-0.04421692084749879, 32'sd0.024148719623482907, 32'sd0.044196236928855305, 32'sd-0.07353718461092719, 32'sd0.08995434789391249, 32'sd-0.00973964532311819, 32'sd0.10273319178107673, 32'sd0.07850584770011369, 32'sd0.014421204133352145, 32'sd-0.034541232394765135, 32'sd-0.068212225908762, 32'sd-0.08601275565751608, 32'sd-0.0850166816986733, 32'sd-0.12196163727176224, 32'sd0.0607119877377119, 32'sd0.09138963009541055, 32'sd0.13595860067650897, 32'sd0.07059068768046758, 32'sd0.021439408232252613, 32'sd-0.10347247661770906, 32'sd0.009662589933341905, 32'sd-0.013190927482030995, 32'sd0.01657518546611199, 32'sd0.06570670868575844, 32'sd0.1420598423216413, 32'sd0.1389429387345234, 32'sd0.02650901575343551, 32'sd-0.07368975219386187, 32'sd0.07762337723642784, 32'sd0.05557455699413748, 32'sd-6.473848544666097e-125, 32'sd0.03899468386777834, 32'sd0.03019020574698921, 32'sd-0.024820544255754928, 32'sd0.07295537473531616, 32'sd0.10745268210987424, 32'sd0.03956063792868838, 32'sd0.038279201091908806, 32'sd0.06293371226154632, 32'sd-0.05915374694942174, 32'sd0.08214239199007414, 32'sd0.012245913951029612, 32'sd0.009609104954432839, 32'sd0.14463830463107868, 32'sd0.18535773229945815, 32'sd-0.0009988860980408654, 32'sd-0.1577687236723455, 32'sd-0.11049841957870594, 32'sd-0.032388303659732526, 32'sd0.09291468153323174, 32'sd0.04704997538065293, 32'sd0.06049809123386848, 32'sd0.02478428165041089, 32'sd0.0833166214932309, 32'sd0.1273736533164638, 32'sd0.09879208429430872, 32'sd-0.005396171640890255, 32'sd-0.00042407219715931107, 32'sd-0.03137789222734357, 32'sd0.022031359272198025, 32'sd0.12649749667655397, 32'sd0.006967714106023203, 32'sd0.004456231649344304, 32'sd0.04337255730824322, 32'sd0.05943713900992499, 32'sd0.011601150943465319, 32'sd-0.0018920356526857382, 32'sd0.1330367680058491, 32'sd0.1821047085397179, 32'sd0.1568076441705863, 32'sd-0.00837387938479496, 32'sd0.024081239604926672, 32'sd0.0471125590488902, 32'sd-0.07210767425586814, 32'sd-0.008965232083344677, 32'sd-0.07354262189638851, 32'sd-0.07349604574788682, 32'sd0.05547877114403137, 32'sd-0.02495227334564866, 32'sd-0.06423604361894064, 32'sd0.026062766029871908, 32'sd-0.0004740929748384164, 32'sd0.07628036514465, 32'sd0.08618831949980572, 32'sd0.06647798919138544, 32'sd0.047143753187660994, 32'sd0.045554831908764803, 32'sd0.01773731150035239, 32'sd-0.040655190341734294, 32'sd0.09696845115279158, 32'sd-0.07825325192904165, 32'sd-0.011876066135560375, 32'sd0.14502307917290486, 32'sd0.1208395554030816, 32'sd0.1158861847183215, 32'sd0.15194078733196545, 32'sd0.19793838855750528, 32'sd0.19878299795524154, 32'sd0.10809025018513993, 32'sd0.13788660276605563, 32'sd0.06725167522022263, 32'sd-0.03295852527893785, 32'sd-0.0597685661855136, 32'sd-0.0609263458931156, 32'sd-0.05547497543242478, 32'sd-0.02570379567183762, 32'sd-0.019310074099918098, 32'sd-0.004547607057224295, 32'sd0.040059828541252424, 32'sd0.03383793546814648, 32'sd0.03512302196358, 32'sd-0.02905581261715049, 32'sd0.015604064964365713, 32'sd0.01794736000484915, 32'sd-3.979143639725808e-127, 32'sd0.03852455226873404, 32'sd-0.10725865222950419, 32'sd0.0029633058295817027, 32'sd-0.025836443849525183, 32'sd0.06722977273240381, 32'sd0.1474969219114412, 32'sd0.12266536544654282, 32'sd0.2074375414390905, 32'sd0.18730437677836428, 32'sd0.0722454795379884, 32'sd0.0216417213503161, 32'sd-0.003226116683366995, 32'sd0.10304088389701167, 32'sd0.20496167143575836, 32'sd-0.03303291239879706, 32'sd-0.004204828460381552, 32'sd-0.02232750318657035, 32'sd-0.0938872410895441, 32'sd-0.10679825500903904, 32'sd-0.01358993131161125, 32'sd-0.014850819810757039, 32'sd-0.14588488211035922, 32'sd0.053184724439496095, 32'sd0.09888135859533269, 32'sd0.010366377529435157, 32'sd0.03707362212624845, 32'sd-0.006878851794494885, 32'sd0.007180665750181103, 32'sd0.10148158623831308, 32'sd-0.02865747091497435, 32'sd-0.0729632232040865, 32'sd0.014781220139154155, 32'sd9.432581351107989e-05, 32'sd-0.03057468650710075, 32'sd0.008331911493019933, 32'sd0.054480049274678845, 32'sd0.07287044225671115, 32'sd-0.010501068404700725, 32'sd0.04117001750625828, 32'sd0.0034742611103384994, 32'sd0.09296451837814972, 32'sd-0.024825310130077823, 32'sd-0.09767437322562661, 32'sd-0.02198438170275982, 32'sd-0.011874704197817058, 32'sd0.15097887310569993, 32'sd0.12334999434919756, 32'sd-0.02052992220251184, 32'sd-0.04170210092634506, 32'sd0.023249170921927628, 32'sd-0.08793542083068151, 32'sd-0.03291675955102371, 32'sd0.12062792768391717, 32'sd0.028407535318801202, 32'sd0.0580495974600841, 32'sd-0.02203482878431593, 32'sd-0.020189210200384923, 32'sd0.062111896283514635, 32'sd-0.11211217578052012, 32'sd-0.01646140813543513, 32'sd-0.025721175669159376, 32'sd-0.027790810734600102, 32'sd-0.04332241443411979, 32'sd0.07001561303653683, 32'sd0.07939740198423452, 32'sd0.0810887080250338, 32'sd0.07235850928452325, 32'sd-0.0727963264335165, 32'sd-0.076572819037173, 32'sd-0.05199647296030992, 32'sd0.06234104091170911, 32'sd0.0547329513548188, 32'sd0.060004019061737066, 32'sd0.17548910338585133, 32'sd0.04315762709916641, 32'sd-0.05687094872568706, 32'sd-0.060818838262101105, 32'sd-0.07704443744558118, 32'sd-0.04243984429366963, 32'sd-0.07732457694656233, 32'sd-0.06938509426945774, 32'sd0.037552143382038154, 32'sd0.029377844933398765, 32'sd3.141929155246688e-125, 32'sd0.059619430467662105, 32'sd-0.017829367771830692, 32'sd0.06097800051804104, 32'sd-0.012967158117176546, 32'sd-0.0029744963827620825, 32'sd-0.03870497283188611, 32'sd-0.14203928561631232, 32'sd-0.10959428272078661, 32'sd0.02379978218232008, 32'sd0.06596017514696707, 32'sd0.03400756906037386, 32'sd-0.09807677354945218, 32'sd0.005910521250332019, 32'sd0.11554592917321954, 32'sd0.1233340885492033, 32'sd0.12650329849353167, 32'sd0.1622948443709107, 32'sd0.1459557351994237, 32'sd0.004959325695021002, 32'sd-0.1492113365059894, 32'sd-0.0178152494786444, 32'sd0.04492556822195426, 32'sd-0.052879730366243605, 32'sd0.0558252628988455, 32'sd-0.06603139991548296, 32'sd-0.04714702682611105, 32'sd2.0460880077652284e-121, 32'sd-4.91552013110011e-126, 32'sd-3.5283243345874725e-116, 32'sd-0.0410371230881414, 32'sd0.022756034271074956, 32'sd0.0636515724928883, 32'sd-0.05262231578759281, 32'sd-0.16919305212883645, 32'sd-0.08027467611299859, 32'sd-0.22876612662534004, 32'sd-0.1163239614882993, 32'sd-0.15086262524517585, 32'sd-0.007686938384571192, 32'sd-0.061980628063792155, 32'sd0.009347852431294915, 32'sd0.06714293741891704, 32'sd0.18484761763794091, 32'sd0.16296174391402116, 32'sd0.16226379696260443, 32'sd0.07506271501182313, 32'sd0.026014459562851523, 32'sd-0.011203399293499845, 32'sd0.11046217618431711, 32'sd0.019307359713746076, 32'sd-0.10778924319890693, 32'sd0.05104621228189906, 32'sd0.07426417386210996, 32'sd0.0644982636259239, 32'sd1.0161707209042237e-121, 32'sd6.802555504451282e-126, 32'sd-4.5736298470034606e-126, 32'sd0.010449512733318126, 32'sd0.021666423433375343, 32'sd-0.025791861762649384, 32'sd-0.06502300358484804, 32'sd-0.1380387348219687, 32'sd-0.10373172312011278, 32'sd-0.028624082520512413, 32'sd-0.05196870342508092, 32'sd-0.16198408489832727, 32'sd-0.09858890099486314, 32'sd0.02721496042937885, 32'sd0.030383682299777455, 32'sd-0.026680021086061, 32'sd0.08415637569146812, 32'sd0.19842326002179037, 32'sd0.0993931453653257, 32'sd0.16654803070477497, 32'sd0.17940165132606178, 32'sd0.10669450040970706, 32'sd0.09370282533929132, 32'sd0.011373230478894901, 32'sd0.010772786508664691, 32'sd-0.05893451537791261, 32'sd0.04873518135732255, 32'sd0.04428210101194502, 32'sd-1.2333519996898975e-124, 32'sd-2.815872720549829e-122, 32'sd3.5621549108665116e-116, 32'sd6.813665942862477e-115, 32'sd0.02479833710627456, 32'sd-0.03709427985463684, 32'sd-0.07607243261799088, 32'sd-0.01968591572407307, 32'sd-0.03612566900875307, 32'sd-0.013163909082180038, 32'sd-0.05357764061824718, 32'sd-0.12357509031178787, 32'sd-0.07416854113297683, 32'sd-0.07436263246948634, 32'sd0.0228269632798326, 32'sd-0.13847153049806832, 32'sd-0.08000275793867478, 32'sd-0.0752747613755981, 32'sd-0.06053353613691297, 32'sd-0.01772035967237587, 32'sd0.0354939600065778, 32'sd0.07816950532171356, 32'sd0.1068147894223477, 32'sd-0.008920041787946491, 32'sd0.11772954573835828, 32'sd-0.014314575346219108, 32'sd-0.0031418450982914972, 32'sd2.3673148148942363e-126, 32'sd7.6697853385915074e-121, 32'sd-5.039383523895771e-124, 32'sd1.0802525244377279e-116, 32'sd5.393407683546833e-118, 32'sd-1.4390027643395278e-121, 32'sd0.020102684664119266, 32'sd-0.0033133864302373147, 32'sd-0.02036379803711943, 32'sd0.008059520979970172, 32'sd0.03633034098268453, 32'sd-0.0029232826438260902, 32'sd0.05173083547052472, 32'sd-0.0798515009520081, 32'sd-0.05585457321412954, 32'sd-0.07332095231935587, 32'sd0.00968972159398283, 32'sd-0.07931673463570336, 32'sd-0.08820125105480918, 32'sd-0.017896652687135736, 32'sd-0.0355411179644632, 32'sd-0.10386765553796812, 32'sd0.0014709360605390165, 32'sd-0.10965696292760786, 32'sd-0.06346564086856289, 32'sd0.03678661095302965, 32'sd-1.690223525616165e-123, 32'sd3.725346657948658e-122, 32'sd8.518982412336166e-118, 32'sd-1.011639789173814e-120},
        '{32'sd6.488737445019305e-124, 32'sd1.458349677517528e-121, 32'sd3.719897038762946e-123, 32'sd-3.383344721457995e-120, 32'sd-3.0298375367123977e-114, 32'sd1.1343363130947191e-117, 32'sd-1.0595375573771016e-119, 32'sd-8.263548228209138e-116, 32'sd2.658796345664038e-121, 32'sd-3.2415044412715635e-121, 32'sd-1.1233352331336062e-120, 32'sd1.1962375888385376e-118, 32'sd-0.010824146370772138, 32'sd0.08625260812290073, 32'sd0.06562420560839004, 32'sd0.03922469149930907, 32'sd3.2683395389359894e-121, 32'sd-6.641181428854168e-115, 32'sd5.892266617987494e-120, 32'sd-5.536640854170719e-116, 32'sd1.1481327151234182e-125, 32'sd-1.358452402462389e-115, 32'sd3.1987629970233554e-121, 32'sd3.922200092151272e-123, 32'sd2.961503608618256e-128, 32'sd-4.816182781980847e-118, 32'sd1.8013072621153346e-125, 32'sd1.5702580137045984e-125, 32'sd-1.1167689377145067e-119, 32'sd-5.866681731506033e-124, 32'sd1.5246022635340045e-125, 32'sd-1.2307115419029795e-124, 32'sd-0.021612850372440866, 32'sd0.016346524936894823, 32'sd0.038268113112574234, 32'sd0.004527037557079283, 32'sd0.020216764198342223, 32'sd0.004550853860791783, 32'sd0.06802891242470012, 32'sd0.009297588242740858, 32'sd0.02973371741930358, 32'sd-0.1114738592484057, 32'sd0.05237867830563451, 32'sd-0.03945535967714271, 32'sd0.02755933654407587, 32'sd0.03787699666824813, 32'sd-0.016182631180591357, 32'sd-0.031550506023215144, 32'sd-0.04618534943009895, 32'sd0.05358009492681087, 32'sd0.004785751012332904, 32'sd0.001135283868642724, 32'sd8.293409047754903e-117, 32'sd7.4947220061077e-115, 32'sd-3.4979152012789926e-122, 32'sd1.4657260446569417e-127, 32'sd2.7822794002595743e-122, 32'sd-4.9138026656099255e-117, 32'sd0.00971271750524911, 32'sd0.009780315651199644, 32'sd0.02060244379032086, 32'sd0.09681082101000386, 32'sd0.08195558689767693, 32'sd-0.06772907589512563, 32'sd-0.030742934658813604, 32'sd0.0297549047572506, 32'sd0.097529800187366, 32'sd-0.07395515374373343, 32'sd-0.011559937855744063, 32'sd-0.0015173864148523071, 32'sd0.10110444294387282, 32'sd-0.0778587678767048, 32'sd-0.0561273079173732, 32'sd0.03767408756097433, 32'sd0.005041040540846364, 32'sd-0.13093117691030146, 32'sd-0.1685349654940835, 32'sd-0.02240274112169517, 32'sd0.044496422468173875, 32'sd-0.03933581448796685, 32'sd0.003045875153929006, 32'sd0.10488433546292242, 32'sd9.464659514360144e-120, 32'sd-5.2662832498525955e-126, 32'sd7.888768001287095e-120, 32'sd-1.344360978434871e-125, 32'sd0.014685506669708132, 32'sd-0.006619820548718476, 32'sd-0.01635839654853042, 32'sd0.03345490839427005, 32'sd0.03734968313109454, 32'sd-0.024574870868338344, 32'sd0.03137056879391356, 32'sd0.05645657358339134, 32'sd0.11633345722578928, 32'sd0.0765808518540633, 32'sd-0.02876288506380127, 32'sd-0.09223956245547489, 32'sd-0.039392311637438907, 32'sd-0.04876114325933114, 32'sd0.011596485616075446, 32'sd-0.030703702588015885, 32'sd-0.10161325694417561, 32'sd-0.13602223449292614, 32'sd-0.14272396481162283, 32'sd-0.15248496964011798, 32'sd-0.14651242929754896, 32'sd-0.06635719099956398, 32'sd0.04667057808025894, 32'sd-0.041506244945549074, 32'sd0.05604782000920399, 32'sd-1.9831329728852147e-126, 32'sd-2.624220982259939e-120, 32'sd0.028038824724696976, 32'sd0.06367527015987964, 32'sd0.0022851559332019524, 32'sd0.0883850946006624, 32'sd0.03149722159307744, 32'sd-0.05216610718129739, 32'sd-0.05599115550912196, 32'sd-0.099906256715757, 32'sd-0.07765789957552567, 32'sd0.018852972397765573, 32'sd-0.018285406870466918, 32'sd0.01669000060645992, 32'sd0.12249667984891445, 32'sd0.07176967585281087, 32'sd0.04790686571925744, 32'sd0.019244318941714057, 32'sd-0.015886701136397615, 32'sd-0.08726122647554735, 32'sd-0.12679280228550938, 32'sd-0.038945352631401906, 32'sd0.0011809218983119998, 32'sd-0.034226167948924933, 32'sd-0.1603912902807286, 32'sd-0.14824562026279275, 32'sd-0.03688564380737896, 32'sd-0.043811778898172456, 32'sd0.018965120755759842, 32'sd9.942755126582453e-128, 32'sd0.04464911747571217, 32'sd0.009916930600598103, 32'sd-0.010126771859733897, 32'sd0.05511595965463598, 32'sd-0.06655870268424624, 32'sd-0.13976560650161035, 32'sd-0.13492570666299128, 32'sd-0.11310349560206788, 32'sd-0.17450327082081854, 32'sd-0.14139985940923977, 32'sd-0.059943192673770934, 32'sd0.00033892648647171033, 32'sd-0.04644662936885451, 32'sd0.13909699546091678, 32'sd0.12096668475384642, 32'sd0.19581685113972136, 32'sd0.21496482467505523, 32'sd0.11663879588947154, 32'sd0.1210779008378394, 32'sd-0.016140657995331292, 32'sd-0.023751834645213986, 32'sd-0.1599093508957856, 32'sd-0.23385852430643206, 32'sd-0.10994147340575101, 32'sd0.013535595786748976, 32'sd-0.05662527868899854, 32'sd0.05301921751294127, 32'sd-1.813901887801097e-126, 32'sd0.012651163195537636, 32'sd-0.03584775963137112, 32'sd0.03783332208709504, 32'sd0.06836115149860575, 32'sd-0.061912219642256926, 32'sd-0.0244602873813775, 32'sd-0.0033037793066526735, 32'sd-0.021401471034121815, 32'sd-0.030253631164929906, 32'sd0.054953433202422255, 32'sd-0.08434910283580126, 32'sd-0.05367698556688867, 32'sd-0.1586001259035085, 32'sd-0.10945928852335296, 32'sd0.1095140057801256, 32'sd0.0948803257963046, 32'sd0.14885204772615715, 32'sd0.15133314532428435, 32'sd0.07258169351463668, 32'sd0.04744934150904189, 32'sd-0.12572636653393862, 32'sd-0.11596330797517526, 32'sd-0.06804982948868046, 32'sd-0.06504282940156711, 32'sd0.07920038233587981, 32'sd-0.04139601871861383, 32'sd-0.019179122076822316, 32'sd0.07701239237287233, 32'sd-0.014647566101178261, 32'sd-0.13638919811347622, 32'sd0.15035330869271815, 32'sd0.10621107664709332, 32'sd0.004630274989444109, 32'sd0.03934437904454465, 32'sd-0.0520426002980358, 32'sd-0.016306687813085818, 32'sd0.02165474065628166, 32'sd0.07780190239119048, 32'sd-0.034055130355316404, 32'sd-0.046028974616883954, 32'sd-0.17712030730887984, 32'sd-0.16922293177032158, 32'sd-0.013341722824174361, 32'sd0.010213411092545751, 32'sd0.16813799827898415, 32'sd0.09232432081852428, 32'sd0.07125854838926922, 32'sd0.016265371002305472, 32'sd-0.12998724895763167, 32'sd0.01920829447490597, 32'sd-0.21502083477342826, 32'sd-0.010361946594450097, 32'sd0.0751808537178779, 32'sd-0.03513823542377371, 32'sd0.038539713773807244, 32'sd-0.0008329742755758185, 32'sd-0.015209271065146903, 32'sd-0.008235805475041495, 32'sd-0.03749092589801185, 32'sd-0.10402123312613962, 32'sd-0.051794216403510444, 32'sd-0.019895930057843538, 32'sd-0.06037665297529768, 32'sd-0.0924441774372546, 32'sd-0.09533591749195432, 32'sd0.03252868175752219, 32'sd-0.11356634028157273, 32'sd-0.13254810120590477, 32'sd-0.09643602278523945, 32'sd-0.01361309469384823, 32'sd-0.030967529425806477, 32'sd0.12926948197045654, 32'sd0.05110152977374827, 32'sd0.13300224062325627, 32'sd0.10156270954529992, 32'sd0.014178150396653435, 32'sd-0.023099848791975075, 32'sd-0.07589910925662068, 32'sd0.058933842211418896, 32'sd-0.07919962200123022, 32'sd-0.15418475460184292, 32'sd-0.08038387180794276, 32'sd0.03596630589779183, 32'sd0.04787831322736632, 32'sd-0.08515569572731327, 32'sd0.06022012867003786, 32'sd-0.07717791671245594, 32'sd-0.004830251839906295, 32'sd-0.15905759915837658, 32'sd-0.1316110263172778, 32'sd-0.11562387468245115, 32'sd-0.12434959294920303, 32'sd-0.08294356208189066, 32'sd-0.060622642128888744, 32'sd-0.001473894934465426, 32'sd0.0024649757716155504, 32'sd0.008692456977246943, 32'sd-0.045047757727173676, 32'sd0.13728553278529168, 32'sd0.10778880271335806, 32'sd0.04714040270865353, 32'sd0.09423008675675519, 32'sd0.07412127980938986, 32'sd-0.0022261586278734405, 32'sd-0.0794053372135446, 32'sd0.024193922717371988, 32'sd0.06403895038278773, 32'sd0.05098403682657048, 32'sd-0.08555088519743581, 32'sd-0.03258234667414466, 32'sd-0.018746668237259297, 32'sd-0.021901046078074374, 32'sd0.016489075639555047, 32'sd-0.10010704830797301, 32'sd-0.03737606702698558, 32'sd0.060661265390684796, 32'sd-0.08258469317523405, 32'sd-0.046808660104594696, 32'sd-0.032021196593126904, 32'sd-0.025101715696131864, 32'sd-0.166557293015494, 32'sd-0.08373648836356506, 32'sd-0.03100947940212345, 32'sd-0.023685067851894687, 32'sd-0.036061355635896596, 32'sd-0.06147197472853432, 32'sd0.054765878904965364, 32'sd0.15208365439037733, 32'sd0.008081173466607779, 32'sd0.080838748524671, 32'sd0.1366337889590966, 32'sd-0.04598380512299452, 32'sd-0.052337147372191736, 32'sd-0.008645025672802932, 32'sd-0.05275396394214648, 32'sd0.023886706412133855, 32'sd-0.17521935795784008, 32'sd-0.038195387295766534, 32'sd0.04255933381165289, 32'sd-0.013488563652728176, 32'sd-0.16513696328368685, 32'sd0.03457382642327417, 32'sd0.011680529091326558, 32'sd0.044750370953368, 32'sd-0.03502280384452264, 32'sd-0.09490609841956997, 32'sd-0.1772143786710417, 32'sd-0.1477360734915634, 32'sd-0.09370271492643119, 32'sd-0.02940739639035582, 32'sd-0.044138839098655354, 32'sd0.05866309525291978, 32'sd-0.0225880000648491, 32'sd0.013613817390955761, 32'sd-0.03977137398418461, 32'sd0.07401488636753172, 32'sd-0.13169974428273365, 32'sd0.03592907921010377, 32'sd0.06545586755543484, 32'sd-0.06013565559515206, 32'sd-0.07734591111057142, 32'sd-0.08537152343083168, 32'sd-0.027976569167204274, 32'sd0.0047810044576888, 32'sd-0.013480302321174595, 32'sd-0.02392190118980154, 32'sd-0.14173983584084074, 32'sd0.08142920674046653, 32'sd0.006142253116873611, 32'sd0.050741893374473546, 32'sd0.0615692655319194, 32'sd-0.023225361902892563, 32'sd-0.05848708124796418, 32'sd-0.033026051196163975, 32'sd-0.11971457925855286, 32'sd-0.07877009790054128, 32'sd-0.06543380846087483, 32'sd0.0896319902085315, 32'sd-0.08771667020941011, 32'sd-0.0003107500204751367, 32'sd0.011910912942242845, 32'sd-0.139671353132366, 32'sd-0.03310841566801187, 32'sd0.008198270464042142, 32'sd-0.03462399477338695, 32'sd-0.17999122082555274, 32'sd-0.018476918137911757, 32'sd-0.07884714038199828, 32'sd-0.15121691504164386, 32'sd-0.13625723564498915, 32'sd-0.010278197114547891, 32'sd-0.03671662997235416, 32'sd0.033822100429514036, 32'sd0.0377688214296862, 32'sd-0.030262650789828167, 32'sd0.034927515899779576, 32'sd0.00948248447224769, 32'sd0.00014787009267981636, 32'sd0.08943737929475715, 32'sd0.0558483549987014, 32'sd-0.07226907977413587, 32'sd0.025005051696676814, 32'sd-0.07204553191448781, 32'sd0.025979824547038222, 32'sd0.08981996169943603, 32'sd0.00631750187906923, 32'sd0.03751244861006963, 32'sd0.09749861990799692, 32'sd-0.0070101118491103405, 32'sd-0.12116131216397621, 32'sd-0.07633180148802073, 32'sd-0.06632404107702566, 32'sd-0.010517039492245429, 32'sd-0.022661448855694908, 32'sd-0.14497866420238856, 32'sd-0.014003816123675218, 32'sd-0.06052961292335413, 32'sd-0.02704470696839548, 32'sd-0.08315379809338758, 32'sd-0.046111995670381954, 32'sd0.06343183515598962, 32'sd0.014935654056487958, 32'sd-0.021110625532123704, 32'sd-0.010623696200989753, 32'sd-0.09952723360031576, 32'sd-0.07949153769604814, 32'sd-0.025745864357329, 32'sd-0.08695010585427887, 32'sd-0.10676407593746805, 32'sd-0.016998269705119504, 32'sd0.15262102408305478, 32'sd0.05383024446790887, 32'sd0.0250364431365715, 32'sd0.020826276577687198, 32'sd0.07423085896355477, 32'sd0.030966598705694896, 32'sd-0.009368421164532207, 32'sd-0.03184280668759022, 32'sd-0.09889992011780693, 32'sd-0.027135431777268407, 32'sd0.06126993633918713, 32'sd-0.15688541138442233, 32'sd-0.07150475860876304, 32'sd-0.04284265714347926, 32'sd0.05904702516013173, 32'sd-0.12783025829228098, 32'sd-0.03214198417101385, 32'sd0.03348402274467706, 32'sd0.0022409009170222434, 32'sd0.052421986591783196, 32'sd0.012572637894292561, 32'sd0.00270270636153084, 32'sd0.0006026911537906508, 32'sd-0.018283579198903565, 32'sd0.006148249604116284, 32'sd-0.06532727088055199, 32'sd0.10623102336147008, 32'sd0.15486723797059906, 32'sd0.21248071376337524, 32'sd0.18797449775005554, 32'sd0.1639870938026984, 32'sd0.01231170945408548, 32'sd-0.011551644143089203, 32'sd0.06878188528000752, 32'sd0.025895004105398647, 32'sd-0.016393583291450534, 32'sd0.040259729535516875, 32'sd0.029094598112490874, 32'sd-0.017266606525858683, 32'sd-0.08010054326286946, 32'sd0.033345369896460794, 32'sd-0.037718452234453206, 32'sd-0.08094363287705511, 32'sd0.0854647748621794, 32'sd0.06234653493950041, 32'sd0.05985053905425757, 32'sd0.13202445322768777, 32'sd-0.02785138912162626, 32'sd-0.07373077769002503, 32'sd0.050548824873035206, 32'sd-0.03341012109499888, 32'sd-0.09231028873645322, 32'sd0.05043686528330139, 32'sd-0.03695136186413169, 32'sd0.05706076888849761, 32'sd0.06336194683641962, 32'sd0.14156310937346803, 32'sd0.15547702238056607, 32'sd0.15151820883114972, 32'sd-0.1212480741206711, 32'sd-0.14277803168686953, 32'sd-0.07175168623960507, 32'sd-0.014860183067513938, 32'sd-0.10709838010605416, 32'sd-0.00373042685255685, 32'sd0.11749587858197129, 32'sd0.13549841702774004, 32'sd-0.09944797862996382, 32'sd-0.11348170113851717, 32'sd-0.08534502569866668, 32'sd0.06262121592014949, 32'sd0.1467722300025567, 32'sd0.0656532558061871, 32'sd-0.05912492040637775, 32'sd0.017287551306291567, 32'sd0.10748259357589114, 32'sd0.004867208757821318, 32'sd1.0554032617824073e-122, 32'sd0.058666872851064596, 32'sd0.031834487091488395, 32'sd-0.052009946394956166, 32'sd0.03896320951044682, 32'sd0.11015049480873823, 32'sd0.07604687620713, 32'sd0.07269598897316495, 32'sd0.11159590902278504, 32'sd0.07600677170635106, 32'sd0.03361501721589253, 32'sd-0.04822801780755324, 32'sd0.028770654109273545, 32'sd-0.03895894775343348, 32'sd0.022067415454427957, 32'sd0.10717769615067942, 32'sd0.06341245058082338, 32'sd-0.023089938700639693, 32'sd-0.10378013664120306, 32'sd-0.09394338629761473, 32'sd-0.06539439535951067, 32'sd-0.042703371506556786, 32'sd0.08786338572690554, 32'sd-0.03849328165585982, 32'sd-0.07211291596912059, 32'sd0.05255410780604806, 32'sd-0.08115293520681517, 32'sd0.06354798213902395, 32'sd0.03070254180109518, 32'sd0.029072616937755126, 32'sd-0.02481923574354794, 32'sd0.028593185957909748, 32'sd0.10391422391088345, 32'sd0.06554905088003486, 32'sd0.12244658920369458, 32'sd0.10789316128798655, 32'sd0.03469754643663681, 32'sd-0.008802051183385971, 32'sd0.007795813978203622, 32'sd-0.04949044020034068, 32'sd0.004461232062796354, 32'sd0.056505483743619744, 32'sd0.018302034112442554, 32'sd-0.007691249353457559, 32'sd0.08025098258605279, 32'sd0.013131716613086484, 32'sd0.06898690199286699, 32'sd0.0885713693052548, 32'sd0.1281823077159311, 32'sd-0.022257532246562375, 32'sd0.07382593507004884, 32'sd0.002274922723138097, 32'sd-0.03013456876648252, 32'sd0.05002431734088469, 32'sd0.058897344934586066, 32'sd-0.009717395063044703, 32'sd0.030054491784665068, 32'sd0.031852614603410635, 32'sd-0.03869969189961939, 32'sd0.024537383767706544, 32'sd-0.028801318807890237, 32'sd0.03066609071913644, 32'sd0.09526327874255686, 32'sd0.13253282987275758, 32'sd0.007841548038718598, 32'sd-0.0038753823274656875, 32'sd-0.028112242020370385, 32'sd-0.1231432967384996, 32'sd-0.08097814469008087, 32'sd-0.0355664455900923, 32'sd0.0193774963686335, 32'sd-0.16731868352105914, 32'sd0.13501510958663732, 32'sd0.07394402110706143, 32'sd0.07078058534851354, 32'sd0.16749966082117348, 32'sd0.020864268988444765, 32'sd-0.0014800979722036586, 32'sd0.10673438939937156, 32'sd0.013115568231917674, 32'sd-0.04516434948065086, 32'sd-0.003686466610368974, 32'sd0.039098029918042905, 32'sd0.08993391456355927, 32'sd-2.5828523240694635e-115, 32'sd0.0047483147804633355, 32'sd0.07363748669485405, 32'sd0.09363527039115407, 32'sd0.06607014424491023, 32'sd0.14222915460719207, 32'sd0.15636681886499829, 32'sd0.07124776678026325, 32'sd-0.06281144020662059, 32'sd-0.14131828901176163, 32'sd-0.19491373884797997, 32'sd-0.21209215183664734, 32'sd-0.13623795602221442, 32'sd-0.08122450688289146, 32'sd-0.2560533175077037, 32'sd-0.2157984702861768, 32'sd-0.017745198881343578, 32'sd0.1216148159528042, 32'sd0.064739710451855, 32'sd0.13290940776286775, 32'sd-0.01422989962478047, 32'sd0.07708443696890062, 32'sd0.04761072720115006, 32'sd0.08599984385721528, 32'sd-0.01319527414109102, 32'sd0.10173270093515395, 32'sd-0.022845025830809922, 32'sd0.016769674384011984, 32'sd0.03665418216887893, 32'sd-0.09280116978884673, 32'sd-0.03534380366175228, 32'sd0.012466085513566132, 32'sd0.09867209326359726, 32'sd0.09505106234561082, 32'sd0.05741722792929883, 32'sd0.07392892093501974, 32'sd0.12746825281306792, 32'sd-0.01520593760872651, 32'sd-0.011238492444580738, 32'sd-0.11895739131423734, 32'sd-0.21831758079074753, 32'sd-0.2119625354534461, 32'sd-0.15527231109510406, 32'sd-0.17139489558135723, 32'sd-0.04540612629691464, 32'sd0.05562730639027494, 32'sd0.03737075028907279, 32'sd0.1702093555163404, 32'sd0.06434691686742584, 32'sd-0.07922091637553298, 32'sd0.04495313356071531, 32'sd-0.019088258277842905, 32'sd-0.04804269540001884, 32'sd0.025914611674041996, 32'sd0.032039069370322075, 32'sd-0.033989937130419576, 32'sd0.007449261634739447, 32'sd0.0003999459179740502, 32'sd0.038409188201492625, 32'sd0.0414459042741836, 32'sd0.007453446007321881, 32'sd-0.08894407773310906, 32'sd-0.017055803921203923, 32'sd-0.0330080829093542, 32'sd0.1414783202236175, 32'sd0.024864515639674043, 32'sd0.009574006398079378, 32'sd-0.10224126489318623, 32'sd-0.18723710075406194, 32'sd-0.190366143606059, 32'sd-0.10780002974785419, 32'sd-0.1601418033086711, 32'sd0.08123214288906733, 32'sd0.06980111753762597, 32'sd0.04621904321877513, 32'sd-0.028638529413145247, 32'sd-0.06673199706757843, 32'sd-0.0708176972058034, 32'sd0.06368517264982945, 32'sd-0.1711328139995444, 32'sd-0.047461800093378935, 32'sd0.06544642942429195, 32'sd0.002703025626440456, 32'sd0.018742976972867566, 32'sd-4.2956998941443995e-125, 32'sd0.03149345580370748, 32'sd0.07226901239936072, 32'sd0.002014665777600909, 32'sd0.0362401976614838, 32'sd-0.14968637760527653, 32'sd-0.15020533506158568, 32'sd0.05648457778349163, 32'sd0.06876745283378104, 32'sd0.06606169063005668, 32'sd-0.01670238209788004, 32'sd-0.02678986619606439, 32'sd-0.11998615757796312, 32'sd0.03835915235941853, 32'sd-0.05544416353713006, 32'sd-0.0060449098149389004, 32'sd0.039275186998369224, 32'sd-0.14574931352420573, 32'sd0.04516822910903821, 32'sd-0.011507933428751376, 32'sd-0.051567900659524754, 32'sd-0.12345116440359982, 32'sd-0.03976372294571723, 32'sd-0.04438989173517708, 32'sd-0.06719084119042287, 32'sd-0.07902311388827957, 32'sd0.0071637986343139155, 32'sd-3.835964838300628e-125, 32'sd8.493348731075391e-120, 32'sd-8.12331930845402e-127, 32'sd-0.04703948969887355, 32'sd-0.1001540020431838, 32'sd-0.04222408020068281, 32'sd-0.043050261362698405, 32'sd-0.08447369552977115, 32'sd-0.13699537352632565, 32'sd-0.06435631835948727, 32'sd0.08098746082348207, 32'sd0.020913213019577465, 32'sd0.003258140924394936, 32'sd-0.08584800606127922, 32'sd-0.003202482136690183, 32'sd-0.09902203980646425, 32'sd-0.12825489709126678, 32'sd-0.030222148013793783, 32'sd0.011953594675817868, 32'sd0.09185220969494025, 32'sd-0.06201543462407154, 32'sd-0.001508139441891865, 32'sd0.04804103294956005, 32'sd-0.053777878531935976, 32'sd-0.06780282304475169, 32'sd-0.10462294037194773, 32'sd-0.01600466529286162, 32'sd0.08060320028086419, 32'sd4.4518737928424804e-123, 32'sd3.529145547256743e-115, 32'sd8.276809523818663e-117, 32'sd0.037066806206471827, 32'sd0.02087554377827074, 32'sd0.0030894377873095123, 32'sd-0.069630464730113, 32'sd-0.0021611361892188864, 32'sd-0.037729238756681806, 32'sd0.05842845681490834, 32'sd-0.03462472720061079, 32'sd-0.2477832552146968, 32'sd-0.23950868390523977, 32'sd-0.2254972436886641, 32'sd-0.16806276289183175, 32'sd-0.15958063808312228, 32'sd-0.06944793616380085, 32'sd-0.07944644567258397, 32'sd-0.134709792243926, 32'sd-0.04280355241681457, 32'sd-0.1646564278415699, 32'sd-0.11523254024276208, 32'sd0.04876107570483584, 32'sd0.007548567628670971, 32'sd0.023108810151191487, 32'sd0.021986128880657728, 32'sd0.04996859371114138, 32'sd0.004021085260411771, 32'sd-2.1803335406265126e-119, 32'sd-3.387583935093391e-122, 32'sd-1.0306110156684668e-119, 32'sd-1.836700203163775e-123, 32'sd0.0548779335118981, 32'sd-0.004430806154082339, 32'sd-0.013822068541040844, 32'sd-0.049316432055595584, 32'sd0.007716004824401696, 32'sd0.0569951782595057, 32'sd-0.01783344039199968, 32'sd-0.08115520923526372, 32'sd0.02951446738290519, 32'sd-0.02958339546890409, 32'sd0.01444774407107634, 32'sd-0.02729504992577218, 32'sd-0.07761649961656375, 32'sd-0.016166608754735065, 32'sd-0.03216750870073801, 32'sd-0.14725696351172227, 32'sd-0.018502669666659123, 32'sd0.007493485858806742, 32'sd0.008036916598366075, 32'sd0.04001351993113484, 32'sd-0.015388331911713807, 32'sd0.036951786449805187, 32'sd0.023433324167008954, 32'sd3.899531486941553e-115, 32'sd-3.537724115158896e-119, 32'sd2.8978423850396113e-123, 32'sd-7.078890333695646e-119, 32'sd-2.5650609372370785e-125, 32'sd-6.535686412005877e-126, 32'sd0.007787772224833098, 32'sd0.04160861633079057, 32'sd0.009588494902423172, 32'sd0.062134501777376526, 32'sd-0.04825492895915235, 32'sd-0.014271799879469867, 32'sd0.028644527528161216, 32'sd-0.009940987768229112, 32'sd0.019334436326901253, 32'sd-0.06755593495819917, 32'sd0.06754867253187039, 32'sd-0.07241327376618653, 32'sd-0.005406061159707221, 32'sd-0.07445859107342342, 32'sd0.04366901543309568, 32'sd0.014973763044066632, 32'sd-0.03065811982020215, 32'sd0.06330561894217097, 32'sd0.12691798037234828, 32'sd0.03222705391578405, 32'sd6.1431585172974844e-120, 32'sd1.1558296758278194e-126, 32'sd-1.1351779594855318e-121, 32'sd6.636114039275493e-124},
        '{32'sd-3.2377184263600217e-125, 32'sd7.234151714272859e-121, 32'sd-8.748865970871176e-120, 32'sd-1.0799746516428345e-122, 32'sd1.110150988043914e-119, 32'sd-9.118805200682455e-128, 32'sd3.0218314546028375e-124, 32'sd1.5138426203531437e-126, 32'sd-3.6507948527809566e-116, 32'sd8.7743584889542e-127, 32'sd-9.893984009326476e-120, 32'sd-1.6185279771667943e-115, 32'sd-0.016780402593839235, 32'sd-0.07274118136574319, 32'sd0.0459354272647276, 32'sd0.034361902631269356, 32'sd-6.765179332007796e-127, 32'sd-2.1145858568102296e-127, 32'sd3.7975244305869283e-122, 32'sd1.6176668773004322e-115, 32'sd-4.1256835710545897e-125, 32'sd5.659013716137368e-124, 32'sd-6.9607120881586265e-115, 32'sd-1.1696469795785843e-117, 32'sd1.1601946882176898e-123, 32'sd1.4672630190808062e-122, 32'sd2.223151475124627e-127, 32'sd7.191293046533079e-123, 32'sd-3.2052361553865504e-121, 32'sd-9.684660885758243e-125, 32'sd-1.709168712754086e-125, 32'sd-3.539015795567846e-125, 32'sd0.10197037048405155, 32'sd-0.019660435382768456, 32'sd0.09018726803446252, 32'sd0.08554782416046174, 32'sd0.01144736978283859, 32'sd-0.0006050654735395577, 32'sd0.02554485197782044, 32'sd0.05771257287950128, 32'sd0.02767538806699913, 32'sd-0.0025063517583002663, 32'sd0.01536672498232676, 32'sd-0.05118188181354909, 32'sd-0.0863193050926008, 32'sd-0.0062062788075899445, 32'sd0.06747966013584177, 32'sd0.06306634007220548, 32'sd0.004820930706172567, 32'sd0.07072017919775898, 32'sd-0.065751235734384, 32'sd0.057504604349349564, 32'sd-4.772975790934799e-123, 32'sd2.726635238627903e-116, 32'sd-8.678683741715888e-127, 32'sd-1.7075101016739932e-125, 32'sd3.4363917229923566e-116, 32'sd5.266138573218839e-126, 32'sd0.06398920827017493, 32'sd0.046581142274992896, 32'sd0.07348344512576997, 32'sd0.034366617641348865, 32'sd0.012595000685903843, 32'sd0.06550609124009908, 32'sd0.0817462268590503, 32'sd0.06457115664050053, 32'sd-0.02973201015115505, 32'sd0.0008127802822051268, 32'sd0.02488994235041537, 32'sd0.13864928517079786, 32'sd0.0706589730550225, 32'sd-0.03372964517207599, 32'sd-0.006154533956422983, 32'sd-0.056761577094160576, 32'sd-0.09555118093019557, 32'sd-0.003416412692662155, 32'sd0.046188009715670025, 32'sd-0.0340426406626726, 32'sd0.07658088058433069, 32'sd-0.0074660518983125914, 32'sd0.014903836666988857, 32'sd0.024485526708382246, 32'sd-4.910644855637368e-115, 32'sd2.6916962376293586e-124, 32'sd-5.4188425935003886e-118, 32'sd1.0236868976635833e-123, 32'sd0.048087778891880484, 32'sd0.0784677479197906, 32'sd-0.013177545079232406, 32'sd0.05697818003257609, 32'sd0.09569364905308742, 32'sd0.06770754875421277, 32'sd-0.035073515388751836, 32'sd0.0075424119644296305, 32'sd0.006398644087606738, 32'sd-0.0888947913380864, 32'sd-0.07812556873381221, 32'sd-0.07948594551493086, 32'sd-0.04779013119827726, 32'sd-0.1265847085351317, 32'sd-0.16282604525306912, 32'sd-0.06770401346326498, 32'sd-0.16806251492457733, 32'sd0.14969020305276967, 32'sd0.16463168112958249, 32'sd0.05923270168201771, 32'sd0.1228400150663818, 32'sd0.0030279631843063265, 32'sd0.05478622220122655, 32'sd-0.10883254212532414, 32'sd0.052062430795406865, 32'sd5.048827460225824e-118, 32'sd-2.807006381543265e-119, 32'sd0.07254949029172673, 32'sd0.048513015430660236, 32'sd-0.02304294545547821, 32'sd0.028334381465477874, 32'sd0.044361820167837636, 32'sd0.02326245496065864, 32'sd0.021626336127633105, 32'sd0.08597576870368787, 32'sd0.09636700708451452, 32'sd-0.07913198944968652, 32'sd-0.06226576686009391, 32'sd-0.08612345510200128, 32'sd0.11706005241561176, 32'sd-0.05344950643888945, 32'sd0.04860260952850767, 32'sd0.13552430617128772, 32'sd0.08423137890860322, 32'sd-0.0024242829886816208, 32'sd0.08593579494304564, 32'sd0.12480005954729317, 32'sd0.1760164751500328, 32'sd0.0607407267843062, 32'sd0.0027495253574176793, 32'sd-0.03389062531042399, 32'sd0.02756969089189966, 32'sd0.014836743526643227, 32'sd0.027945342001467262, 32'sd-3.630299513280629e-125, 32'sd0.046755629310339775, 32'sd-0.07460803442120548, 32'sd0.05784538030294469, 32'sd0.018959084092476805, 32'sd0.00679329470448079, 32'sd-0.006589380152103183, 32'sd0.018965150580330988, 32'sd0.0942102135952643, 32'sd0.19648046289306126, 32'sd0.15869255326629844, 32'sd-0.14378947038650278, 32'sd-0.16389219837503116, 32'sd-0.09112501206671143, 32'sd-0.13240555361723344, 32'sd-0.01553364941820381, 32'sd-0.03510861942053354, 32'sd0.013019066619265962, 32'sd0.003148023021797891, 32'sd0.01595583383425318, 32'sd0.08619773672334065, 32'sd-0.05726777939981787, 32'sd-0.052298841513300484, 32'sd-0.006004963560201174, 32'sd-0.014842057367616165, 32'sd0.05691147578018685, 32'sd0.06603040053055992, 32'sd0.044197318442406985, 32'sd2.448862511622722e-124, 32'sd0.024953504263029704, 32'sd-0.016729912722489887, 32'sd0.03470562200065312, 32'sd0.12584473304998572, 32'sd0.07361634620306264, 32'sd0.0881708317236148, 32'sd-0.0708949931979428, 32'sd0.04451650790022111, 32'sd-0.0005225241989142686, 32'sd-0.07494339898882371, 32'sd-0.11126249625329457, 32'sd-0.14940440660901502, 32'sd-0.10040751480216141, 32'sd-0.0868426765316142, 32'sd-0.07103290852029903, 32'sd-0.13469998354518684, 32'sd0.013756964858823289, 32'sd-0.07359005803338767, 32'sd-0.0361145168075847, 32'sd0.029990506917807285, 32'sd0.07748607944291819, 32'sd0.08330455093046725, 32'sd0.07394953470915183, 32'sd-0.017779873961256205, 32'sd-0.0033629399188820097, 32'sd-0.03666666690050619, 32'sd0.030724972839239334, 32'sd0.03338016484015873, 32'sd0.04068896328134678, 32'sd0.06881126434828093, 32'sd-0.029913555778675476, 32'sd-0.02265693946579919, 32'sd0.015058793296734605, 32'sd0.05481981783740984, 32'sd0.09599961295135863, 32'sd0.00016760554852922156, 32'sd-0.04552287455265453, 32'sd0.10121013112514385, 32'sd-0.0415230575209447, 32'sd-0.05025085620104082, 32'sd-0.15595392804504837, 32'sd-0.10683410047121852, 32'sd-0.12753425414887054, 32'sd-0.08437836677334229, 32'sd-0.08519406404203522, 32'sd-0.0361321878573114, 32'sd0.056513584192228364, 32'sd-0.019014841031318837, 32'sd0.09602646640902338, 32'sd-0.00815118425651632, 32'sd0.053209198936710875, 32'sd0.020015915427236766, 32'sd0.06857335178158355, 32'sd0.07741976171342142, 32'sd0.06846825854939703, 32'sd0.007340327570830104, 32'sd-0.03729908413127939, 32'sd0.009470439242181565, 32'sd0.07250079706270547, 32'sd-0.011092244450359846, 32'sd0.05807288700143988, 32'sd0.06387962023545901, 32'sd0.05012442736341003, 32'sd-0.03491585438575187, 32'sd0.15424257022749546, 32'sd0.044900048966698636, 32'sd0.10843372318499553, 32'sd0.008712015895201345, 32'sd-0.15701949124750056, 32'sd-0.1472645999291356, 32'sd-0.0720085174779613, 32'sd0.052486169598073326, 32'sd0.03224992617598533, 32'sd0.03615461040216213, 32'sd-0.02773803991359973, 32'sd0.06655631165490693, 32'sd0.13396254547840916, 32'sd0.017105729534284388, 32'sd0.03231381674506628, 32'sd0.11698032937826666, 32'sd0.047866120198426336, 32'sd0.09130449246003008, 32'sd-0.08196978571380656, 32'sd0.03241493211407251, 32'sd0.04662375147961639, 32'sd0.04850750014320198, 32'sd-0.057808115393563834, 32'sd0.11647372139210416, 32'sd-0.038971744424513226, 32'sd0.054595578707473266, 32'sd-0.012832664427677977, 32'sd0.1083454063257616, 32'sd0.05908057857285168, 32'sd0.06753078833890175, 32'sd0.04917628728314197, 32'sd0.037790074356760406, 32'sd-0.0880100842761273, 32'sd-0.21471929144476984, 32'sd-0.049436370374548386, 32'sd0.07297990505042863, 32'sd0.03767892323367912, 32'sd-0.07970261215000916, 32'sd-0.03190770603801374, 32'sd0.07696387531106824, 32'sd0.10920189851820486, 32'sd0.0028065146781277644, 32'sd0.07953155581430141, 32'sd0.022435891032188206, 32'sd0.057088119156236856, 32'sd-0.034816238719304934, 32'sd0.02780150068758277, 32'sd0.08563282844038238, 32'sd0.056788488847609335, 32'sd0.038476707285553594, 32'sd0.0782707282974474, 32'sd0.004106676392503571, 32'sd-0.018458867176303656, 32'sd-0.03306794862778894, 32'sd0.020877015411745806, 32'sd0.06305676809652312, 32'sd0.128837503357193, 32'sd0.07991094205621405, 32'sd0.09680133392880802, 32'sd0.006162890008462407, 32'sd-0.07263823017709743, 32'sd-0.2092100889491084, 32'sd0.026609553502909514, 32'sd-0.11378293911920478, 32'sd-0.026170698055567893, 32'sd-0.04411846686658737, 32'sd0.012177787450993441, 32'sd-0.09950309866278893, 32'sd-0.022765568086575677, 32'sd0.0211218865294149, 32'sd-0.10328780181496058, 32'sd-0.047387569361306545, 32'sd0.02787563829469798, 32'sd0.04228611638521322, 32'sd0.024859298411915358, 32'sd0.06282082441253202, 32'sd-0.012804720099103922, 32'sd0.06650351867334399, 32'sd0.028572425445835766, 32'sd-0.11459041215070745, 32'sd0.040881603066965734, 32'sd0.1277650308725058, 32'sd0.07971835736667959, 32'sd0.10312880503930154, 32'sd0.1615822137276811, 32'sd0.09507471814731377, 32'sd0.06412447341446369, 32'sd0.10207013830644507, 32'sd-0.2463468499050885, 32'sd-0.25640023475126433, 32'sd-0.01377855020844971, 32'sd-0.06430634743291833, 32'sd0.018958034322660175, 32'sd-0.06547617612606711, 32'sd-0.13134464900383064, 32'sd-0.04844745885941327, 32'sd-0.07231875209393022, 32'sd-0.06131510187094244, 32'sd-0.05975277440779656, 32'sd-0.09808185669190558, 32'sd0.05565672157800033, 32'sd-0.004949368985275987, 32'sd-0.014343133085453737, 32'sd-0.009248659407272923, 32'sd-0.0739344220919766, 32'sd0.061720002295453824, 32'sd0.013993816697626487, 32'sd0.003261456415398303, 32'sd0.04521901195350613, 32'sd0.03564121970236329, 32'sd0.10594908005896055, 32'sd0.10750469227247059, 32'sd0.025741354809715334, 32'sd0.21525853938679196, 32'sd0.17111707466062429, 32'sd-0.06847485064396895, 32'sd-0.15943055230094538, 32'sd-0.12240278924487766, 32'sd-0.10922882948017616, 32'sd0.026572488353790134, 32'sd-0.07799447839311151, 32'sd-0.02554471963555331, 32'sd-0.003931896122641675, 32'sd-0.05019780533565589, 32'sd-0.13819384905189047, 32'sd-0.018920536626805616, 32'sd-0.03363180433459938, 32'sd-0.12111379567318588, 32'sd-0.11698692201656405, 32'sd-0.1466702529089415, 32'sd-0.03640743864205428, 32'sd0.050593347789959414, 32'sd-0.08165108787088339, 32'sd-0.01820325290210727, 32'sd-0.0856812058646542, 32'sd-0.028734942767381217, 32'sd0.08282721603433583, 32'sd0.13073803687657443, 32'sd0.19431087708585293, 32'sd0.03642231300675295, 32'sd-0.011344889327547179, 32'sd0.16715060027270662, 32'sd0.005257410168625732, 32'sd-0.09238937767111925, 32'sd-0.20881065721021477, 32'sd-0.15147644195514884, 32'sd-0.03587474687202345, 32'sd0.0074011844810784955, 32'sd0.011468796720107094, 32'sd-0.05217810012244053, 32'sd0.08165121784572617, 32'sd-0.05514741920464322, 32'sd-0.007794441215525713, 32'sd-0.06402310975705573, 32'sd-0.068880175835409, 32'sd-0.08600620093183434, 32'sd0.05739665011283851, 32'sd-0.04571523098517288, 32'sd-0.010020187028003833, 32'sd0.14069737526062823, 32'sd0.010328983679043809, 32'sd0.02747237678984911, 32'sd-0.0595349537018039, 32'sd0.04359614240952897, 32'sd0.08995524457182515, 32'sd0.005749601161120194, 32'sd-0.007045694554087142, 32'sd0.03405946178930492, 32'sd0.0610977122087885, 32'sd0.14395119172496496, 32'sd0.028898642069471944, 32'sd-0.06930331790507055, 32'sd-0.14856547347127078, 32'sd-0.09957762688108199, 32'sd-0.05962556506600196, 32'sd0.04958330695788825, 32'sd0.002313200170063752, 32'sd0.03352128187832647, 32'sd0.07976852885874568, 32'sd0.016042252442197747, 32'sd-0.0239538654250906, 32'sd0.11246591312165088, 32'sd-0.022088043901723975, 32'sd-0.018980582799280356, 32'sd-0.13090202836806014, 32'sd0.014151710991603754, 32'sd0.042473870042410135, 32'sd-0.02537969388348746, 32'sd0.008362319445912272, 32'sd0.06255930216872585, 32'sd-0.040120961110642714, 32'sd0.05257761858869711, 32'sd-0.09609739467501788, 32'sd0.027384391110889333, 32'sd0.01802301259247109, 32'sd0.060608725139208806, 32'sd0.03725468033531117, 32'sd0.1319580267525676, 32'sd0.03987931979398692, 32'sd-0.10773282220425034, 32'sd-0.1547626794851599, 32'sd-0.15474407290475486, 32'sd0.09919210056082711, 32'sd0.01719362673925357, 32'sd-0.005146027373841968, 32'sd0.10296678419806826, 32'sd0.12713893167939277, 32'sd-0.02164274737044285, 32'sd-0.03610309054525187, 32'sd0.15197697218428688, 32'sd0.0006935988907379826, 32'sd-0.12888889338718004, 32'sd-0.06971190375197885, 32'sd-0.08752568420135669, 32'sd0.060417655306106675, 32'sd0.030332594280496068, 32'sd0.030801437970245735, 32'sd0.023180965233769012, 32'sd0.036886700445842385, 32'sd0.07683013806562589, 32'sd-0.019418301296923648, 32'sd0.1064854355601379, 32'sd0.048483817862505205, 32'sd0.13611454347815813, 32'sd0.0990144196816753, 32'sd0.025402777371381684, 32'sd-0.0689364722911082, 32'sd-0.018153554465027675, 32'sd-0.24596441892266152, 32'sd-0.17755982605171974, 32'sd0.04038892716991789, 32'sd-0.04333761567069619, 32'sd0.07375492775992644, 32'sd0.02898940913127976, 32'sd0.05668208400167147, 32'sd0.1246788813368823, 32'sd-0.02199039273281858, 32'sd-0.030966400759942253, 32'sd0.02917048590208996, 32'sd-0.004575376960828975, 32'sd-0.08877766093007547, 32'sd-0.15958845312910586, 32'sd-0.05205007656110162, 32'sd-1.026879866155344e-120, 32'sd0.06285040815322193, 32'sd-0.036496837221705714, 32'sd0.041896894253486076, 32'sd-0.007587543597705484, 32'sd-0.008863920836734469, 32'sd0.06935894366861753, 32'sd0.1062277145735056, 32'sd0.11609110328296328, 32'sd-0.019460645622517515, 32'sd0.08347132007085302, 32'sd-0.06908637469873094, 32'sd-0.22659021352605838, 32'sd-0.25092989209249006, 32'sd-0.08509166704461472, 32'sd0.07875575592877292, 32'sd0.11468991869333196, 32'sd0.08425612397841234, 32'sd0.1374969674068745, 32'sd-0.03922567867049611, 32'sd0.03872430942532835, 32'sd0.043204099803157876, 32'sd-0.07075412448493594, 32'sd-0.13558030574934885, 32'sd-0.02486913888572102, 32'sd0.03843573231753473, 32'sd-0.017125447662870743, 32'sd0.04351516598720108, 32'sd0.00944294877657804, 32'sd-0.06766605245500514, 32'sd0.11888009433749092, 32'sd-0.02377280885876518, 32'sd-0.016262375988713506, 32'sd-0.014149228142501599, 32'sd-0.032483203512843804, 32'sd-0.05630339685540032, 32'sd-0.19054144622056252, 32'sd-0.05963924100586332, 32'sd-0.1520041898736932, 32'sd-0.13199418109848826, 32'sd-0.16456645283596238, 32'sd-0.07654617391428259, 32'sd0.016319113140854363, 32'sd0.12829372279601622, 32'sd0.11993876044781956, 32'sd0.11440044522670771, 32'sd-0.010536141576857857, 32'sd-0.0560145113051065, 32'sd0.12586004914980956, 32'sd0.07287159405556307, 32'sd0.03810764273558824, 32'sd-0.10676591071604408, 32'sd0.08049588008696267, 32'sd-0.10775100766864704, 32'sd0.09260645776910031, 32'sd0.022810880084908683, 32'sd0.057542581424988866, 32'sd0.02211612922680536, 32'sd-0.07008980877514726, 32'sd0.09475013884128543, 32'sd-0.03335200535342119, 32'sd0.011846891960332914, 32'sd0.01446147177516448, 32'sd-0.21558762630413175, 32'sd-0.13159797780310467, 32'sd-0.07392565518738207, 32'sd-0.197502219013401, 32'sd-0.20512826122250663, 32'sd-0.2372043159036882, 32'sd-0.07197995720534203, 32'sd0.0013482959101652422, 32'sd0.15478911131395762, 32'sd0.015494272409308295, 32'sd-0.03202295552152674, 32'sd0.050157383385799406, 32'sd-0.03096761515596711, 32'sd-0.07859630902337511, 32'sd-0.08187138026210615, 32'sd-0.09515646385224856, 32'sd0.007191808888364518, 32'sd-0.04329432678018249, 32'sd-0.12567850674774925, 32'sd-0.028771254081963255, 32'sd0.035982211993436465, 32'sd-2.7694158122013576e-119, 32'sd0.00965063825709373, 32'sd0.041550435420947406, 32'sd0.04494057867725201, 32'sd-0.11295343477927612, 32'sd-0.09532247216761035, 32'sd0.04109083535154226, 32'sd-0.06727099883278867, 32'sd-0.06684423873453316, 32'sd-0.18426156553572967, 32'sd-0.143535015292284, 32'sd-0.09333019242353618, 32'sd-0.11859917995883731, 32'sd-0.04712710691211332, 32'sd-0.020558114736455933, 32'sd0.03804124552586484, 32'sd0.052994138847603976, 32'sd0.11140960926517596, 32'sd0.01841253155341606, 32'sd-0.03878595375906018, 32'sd-0.0033968523985709246, 32'sd0.033483066866951496, 32'sd0.038153135435979806, 32'sd0.08351273066069956, 32'sd-0.08618088331048579, 32'sd-0.10080902243446821, 32'sd0.07470981337233223, 32'sd0.07329959372303298, 32'sd0.08882301713004101, 32'sd0.040183755143639484, 32'sd0.04461070497917627, 32'sd0.044402447040223406, 32'sd-0.021667181973657038, 32'sd-0.10471558025315096, 32'sd-0.10904137280596084, 32'sd-0.1240996802291333, 32'sd-0.08236865010721123, 32'sd-0.10846760126937098, 32'sd-0.14695864122517546, 32'sd-0.16816844683452176, 32'sd0.027482273459048266, 32'sd0.11468338765867507, 32'sd-0.080095234832039, 32'sd0.04722933422926645, 32'sd-0.048866688785327614, 32'sd0.05614740234671968, 32'sd0.05604748614703791, 32'sd0.08857248797579724, 32'sd-0.018932589304446263, 32'sd0.010998344979721424, 32'sd0.10017212894318445, 32'sd-0.010290498752032824, 32'sd-0.027399985126686368, 32'sd0.05131854105967446, 32'sd-0.002439649859511906, 32'sd-0.05277858799016298, 32'sd0.16088911329141858, 32'sd0.04902349229470387, 32'sd-0.0018674611287494468, 32'sd-0.09850726390972864, 32'sd0.006514956905578199, 32'sd-0.08852946666357799, 32'sd0.0323439634876895, 32'sd-0.02242668702819802, 32'sd-0.0024514948413182185, 32'sd-0.06429710309539333, 32'sd-0.06865837782391947, 32'sd-0.14165912535904632, 32'sd-0.061686877209097074, 32'sd0.05064970685505374, 32'sd0.01617848775764498, 32'sd0.053560743066760265, 32'sd0.028761275795323407, 32'sd-0.00667048991040583, 32'sd0.10089815212502509, 32'sd0.12884537284548153, 32'sd-0.005520438344979145, 32'sd0.15228317732332966, 32'sd-0.0860711455288721, 32'sd0.06785002456690992, 32'sd0.009591828166118801, 32'sd0.0068365800225302685, 32'sd-0.01857597287004273, 32'sd0.0491273257889382, 32'sd-1.7957702448648026e-123, 32'sd0.10022922761614103, 32'sd0.053595639191093725, 32'sd-0.007892898673585376, 32'sd0.03553079968695975, 32'sd0.1059518584149222, 32'sd0.05838906043417286, 32'sd0.007892548083867301, 32'sd-0.004517143324210684, 32'sd-0.031211293239519804, 32'sd0.047063133449478274, 32'sd0.04992771538597303, 32'sd0.05390246242208289, 32'sd0.018080365814437994, 32'sd0.036289277629596536, 32'sd-0.050718351997607845, 32'sd0.11655337853453289, 32'sd0.031180108831011695, 32'sd0.022313555856882668, 32'sd-0.03290247279182745, 32'sd0.057788640701861724, 32'sd-0.007834288338458312, 32'sd-0.039917897321307565, 32'sd0.037488324249397915, 32'sd0.03183571804482073, 32'sd0.0025190437082714067, 32'sd0.045371580640977176, 32'sd3.633534558326567e-116, 32'sd6.408146193142333e-127, 32'sd-1.9050747004485037e-124, 32'sd-0.03707163525667157, 32'sd0.06847069243598529, 32'sd-0.01574860853079181, 32'sd0.12066193048352708, 32'sd0.07908954458901438, 32'sd0.0208309033051529, 32'sd0.027394144465068715, 32'sd-0.048355811272365316, 32'sd-0.15794992574787775, 32'sd0.07064866139126992, 32'sd0.053523400275101975, 32'sd0.03733734825034707, 32'sd0.06684999610556355, 32'sd-0.03470995967527321, 32'sd0.09318463774725894, 32'sd0.1086358003437309, 32'sd0.037177514045677464, 32'sd0.06035367322915915, 32'sd0.037953061714092066, 32'sd0.07141615104443075, 32'sd0.0354420966449362, 32'sd0.011726688172954617, 32'sd0.10870124390369977, 32'sd0.06702540261788949, 32'sd-0.024686214083873583, 32'sd2.1214722395234036e-116, 32'sd-1.0213890161891378e-120, 32'sd2.4146013208149917e-124, 32'sd0.02030433452409274, 32'sd0.03444012088170569, 32'sd-0.008263081016816588, 32'sd0.034343017677041794, 32'sd0.026636824783516, 32'sd-0.11971844319502063, 32'sd-0.04813183908559983, 32'sd0.03369040362800076, 32'sd-0.08744013897341127, 32'sd0.11480396235976871, 32'sd0.13101085388665118, 32'sd-0.019141971398785398, 32'sd0.04264605015897233, 32'sd0.030169510329091376, 32'sd0.02912758960112503, 32'sd0.02480989765768118, 32'sd0.022959144294550045, 32'sd-0.05962351969441287, 32'sd0.04527197464431951, 32'sd0.0665571129381523, 32'sd0.07208370343501526, 32'sd0.08734420635826673, 32'sd-0.00837475671597174, 32'sd-0.07090137524852874, 32'sd2.5238427862770778e-05, 32'sd1.1286894950080076e-119, 32'sd1.0689568359551586e-123, 32'sd8.51747886828493e-119, 32'sd-1.7897577979021327e-123, 32'sd0.07485834569736328, 32'sd0.04602027752337099, 32'sd0.028669735046964965, 32'sd-0.08848406954487503, 32'sd-0.07603372215874925, 32'sd-0.05276473209647276, 32'sd-0.007378452853475012, 32'sd-0.040800483580425775, 32'sd-0.043640627795155325, 32'sd-0.021414609489249527, 32'sd-0.053552039824024775, 32'sd-0.07794824607946921, 32'sd0.07110070649893531, 32'sd0.054545944771491106, 32'sd-0.010693830443784892, 32'sd-0.05102515096292146, 32'sd-0.04700692474814752, 32'sd-0.059447448139814736, 32'sd-0.0677594757594205, 32'sd0.05405990271983448, 32'sd0.04628544637781222, 32'sd-0.0158371435953482, 32'sd0.06632356669271348, 32'sd-3.3424068727229295e-120, 32'sd-1.7439989597258644e-117, 32'sd-1.4497480476509674e-125, 32'sd7.076802163537027e-126, 32'sd2.2437787180351958e-122, 32'sd-1.8555159196865518e-116, 32'sd0.08249938162269209, 32'sd0.025494410157920488, 32'sd0.0011155669224116116, 32'sd0.06047659417063877, 32'sd0.022695063884982193, 32'sd0.05426282419970601, 32'sd0.02208400026535334, 32'sd0.021210794198270193, 32'sd0.07526133335868332, 32'sd-0.08111121090826473, 32'sd-0.0488821424169209, 32'sd-0.10628633354953816, 32'sd-0.014333965481206364, 32'sd0.09395825724988789, 32'sd-0.052242283628473614, 32'sd0.02760923971674756, 32'sd-0.11110304510494455, 32'sd0.03600485488789786, 32'sd0.09856690130021066, 32'sd0.1194798933410599, 32'sd-1.6538044978985532e-118, 32'sd-1.4062500253461746e-118, 32'sd3.12087610899404e-123, 32'sd7.153138379127857e-115},
        '{32'sd-4.619365801370348e-127, 32'sd7.091415151477529e-125, 32'sd-1.3210746544126367e-124, 32'sd-4.280407693341764e-115, 32'sd2.716854661760557e-125, 32'sd-8.127155954629054e-122, 32'sd6.915976980962139e-120, 32'sd1.9878578963638877e-125, 32'sd1.3628724187831272e-125, 32'sd-1.5635661887772431e-117, 32'sd-5.3535828829963606e-120, 32'sd-1.5942499420711375e-115, 32'sd0.00943768501375486, 32'sd-0.034983535949679796, 32'sd-0.012577760771871985, 32'sd0.04008875507716247, 32'sd2.8140698382721805e-122, 32'sd-1.0277372755969544e-127, 32'sd-1.5868636306288766e-117, 32'sd-1.5634748053361934e-117, 32'sd3.606228403875614e-122, 32'sd3.6754129345387623e-116, 32'sd2.354639878938919e-116, 32'sd-4.9524338367821044e-117, 32'sd-7.160108724180991e-121, 32'sd2.6337856083811643e-124, 32'sd-2.082394431018769e-122, 32'sd2.701062297060474e-119, 32'sd-2.8513447832135685e-117, 32'sd1.2423605802740723e-118, 32'sd-4.1574852647031575e-117, 32'sd3.739940074416603e-122, 32'sd-0.015149986883861804, 32'sd-0.020179153529667333, 32'sd0.0024939380286306606, 32'sd-0.02378278977268682, 32'sd0.010925820989197409, 32'sd-0.08357520214138772, 32'sd0.015152200483527556, 32'sd0.033993579776836945, 32'sd-0.035810888844966304, 32'sd-0.04031611574904824, 32'sd-0.06393725147656494, 32'sd-0.02909754429455986, 32'sd-0.010741747695854363, 32'sd0.027596416736339877, 32'sd-0.046391211327339345, 32'sd0.030063292164268913, 32'sd0.002002816959662759, 32'sd0.03812550030329225, 32'sd-0.07237506166016978, 32'sd0.040975904104969665, 32'sd3.293663754013448e-119, 32'sd-8.300556764580774e-124, 32'sd1.3410104733489348e-122, 32'sd3.738278812999944e-125, 32'sd-3.7549847241425995e-119, 32'sd7.473644100300861e-115, 32'sd-0.0331793378071042, 32'sd0.019782951404620906, 32'sd-0.030184074241273572, 32'sd-0.009519447785382145, 32'sd0.011863922290383353, 32'sd-0.09520913770484707, 32'sd-0.03544776641733841, 32'sd-0.12975675645662257, 32'sd0.03203085993502181, 32'sd-0.014418380980909936, 32'sd-0.05538097433035306, 32'sd0.05481603626999774, 32'sd-0.08635146656202602, 32'sd0.054951606610269196, 32'sd0.02517710090881198, 32'sd0.07061165333480807, 32'sd0.1037974093700708, 32'sd-0.010834427162125838, 32'sd0.015255129159558643, 32'sd0.0671835236592091, 32'sd0.0634578118256016, 32'sd0.01655475493511173, 32'sd0.0636507886854949, 32'sd-0.012020264577941975, 32'sd-3.752949453222708e-127, 32'sd1.2314020854869987e-120, 32'sd2.0929196455965146e-122, 32'sd1.7243034427568744e-125, 32'sd0.008998881336346872, 32'sd-0.004437402049183413, 32'sd0.05922957537050492, 32'sd-0.021016058404883586, 32'sd-0.04465922480170907, 32'sd-0.0027717639424355693, 32'sd0.15656884247002797, 32'sd-0.105105695717663, 32'sd0.08941558556310633, 32'sd-0.11875105248422925, 32'sd-0.11661048514815786, 32'sd-0.03515923905511927, 32'sd-0.13044062816730492, 32'sd-0.03045625688300296, 32'sd-0.010568615475788596, 32'sd-0.10585219541193097, 32'sd-0.13611845333355937, 32'sd-0.12135210205404078, 32'sd-0.038809954126773474, 32'sd-0.031420639025199794, 32'sd0.015428501303437916, 32'sd0.005203734150229658, 32'sd0.025529259626834274, 32'sd-0.029589132714782588, 32'sd-0.010396740350366493, 32'sd-2.6856821558696036e-124, 32'sd-1.565874835667605e-122, 32'sd-0.01643819091675089, 32'sd0.03050988888299819, 32'sd-0.024975240447509692, 32'sd0.027434706160669987, 32'sd0.02653103915385714, 32'sd0.020769839919912422, 32'sd0.04402440752183321, 32'sd0.003559551011771442, 32'sd-0.019597421786120037, 32'sd0.12910004967247926, 32'sd0.06607947284966585, 32'sd0.07983872781764942, 32'sd0.0930812958134177, 32'sd-0.04702374692933276, 32'sd0.0009622276785646547, 32'sd-0.028488288051178236, 32'sd-0.014267586934855327, 32'sd0.10569627295289503, 32'sd0.04386665704043037, 32'sd-0.15497274635652714, 32'sd0.032039061017523046, 32'sd0.025079306532973578, 32'sd-0.0431223650965925, 32'sd0.10421713884025705, 32'sd-0.04477844376486167, 32'sd0.01753009079656385, 32'sd0.03441374203021823, 32'sd-1.0073906050545002e-121, 32'sd0.06387735961971779, 32'sd0.035344013742151695, 32'sd0.09435621969297084, 32'sd-0.08219611432197219, 32'sd-0.02012433080249903, 32'sd-0.031759637188985, 32'sd-0.011363345714020381, 32'sd0.04368719211749155, 32'sd0.04255252090594148, 32'sd0.06039741837170234, 32'sd0.10716341113951487, 32'sd0.022562920926351603, 32'sd0.009880140277928816, 32'sd-0.12600784056470352, 32'sd-0.0993804682227158, 32'sd-0.040710575053807305, 32'sd0.052429354112457846, 32'sd0.043134057067482, 32'sd0.07103436548943562, 32'sd0.056103259086373904, 32'sd0.06483943299199156, 32'sd-0.1141451361306901, 32'sd-0.08734231188439343, 32'sd0.04068099719379711, 32'sd0.014016244636200098, 32'sd-0.020361335255628082, 32'sd-0.011828185238499656, 32'sd2.3932096371026015e-122, 32'sd-0.011777664128254884, 32'sd0.0020459210719514748, 32'sd0.042305821643058746, 32'sd-0.0628419100331796, 32'sd0.05672888378638953, 32'sd0.02777658219025681, 32'sd-0.06201901703786801, 32'sd0.03929006048188163, 32'sd0.05587584638264494, 32'sd0.012627315998894812, 32'sd0.13891512218221694, 32'sd0.032970200598200765, 32'sd0.017195008104868577, 32'sd0.10818079390762785, 32'sd0.08374411944726615, 32'sd-0.0342712810011994, 32'sd-0.0016639188572727926, 32'sd0.06543620137422314, 32'sd-0.07935243588780296, 32'sd-0.0792533909326142, 32'sd0.05935177103313216, 32'sd-0.11113971047657498, 32'sd0.046104697295001065, 32'sd0.04812513808353086, 32'sd-0.10106351781858323, 32'sd-9.102848952093012e-05, 32'sd-0.058384095405064354, 32'sd0.006593512668638271, 32'sd-0.05151820695809784, 32'sd0.003567044059097422, 32'sd-0.03429274415352214, 32'sd-0.002817157574813972, 32'sd0.04820746049764293, 32'sd0.001492539264587271, 32'sd0.03828542942189689, 32'sd0.11394326772187226, 32'sd0.043708377732379254, 32'sd-0.03143070248926076, 32'sd0.05265860260026799, 32'sd0.056000732839864564, 32'sd0.1632874975318366, 32'sd0.032471011190661724, 32'sd0.07864230286737707, 32'sd0.09272367057115334, 32'sd-0.08550294826975818, 32'sd0.0319009951783172, 32'sd-0.07702494414848825, 32'sd0.05383244526555562, 32'sd0.07058093596661112, 32'sd-0.07124133890373402, 32'sd-0.19990908991846298, 32'sd-0.06058554396917792, 32'sd-0.06895043330907631, 32'sd-0.057600363424951825, 32'sd-0.018349157824974635, 32'sd0.04304313992781878, 32'sd-0.05112940084649799, 32'sd-0.07977807688478339, 32'sd0.02018587295451753, 32'sd-0.015510303613016155, 32'sd0.022207105074517324, 32'sd-0.038611075554399354, 32'sd0.051417976516773135, 32'sd0.15634864252815128, 32'sd0.13097766372864758, 32'sd0.06451153613609234, 32'sd-0.04599646504823444, 32'sd0.11104810938030087, 32'sd0.06454377119397428, 32'sd0.07165173202781742, 32'sd-0.06451665788208048, 32'sd-0.08334588227736651, 32'sd0.01104415511099318, 32'sd-0.05992689802672821, 32'sd-0.05639747329443693, 32'sd-0.04749461917858326, 32'sd-0.12840501140914845, 32'sd-0.12397981661888074, 32'sd0.013599612286579013, 32'sd-0.06193830209401793, 32'sd-0.05592275206281946, 32'sd0.03704269343117099, 32'sd-0.00768041010627808, 32'sd0.01941794743765349, 32'sd0.0022564305064288583, 32'sd0.07711794505768044, 32'sd-0.06720521850051549, 32'sd0.0055516642828830984, 32'sd0.06631396466627623, 32'sd0.06038756002592465, 32'sd0.023704200672227553, 32'sd0.12732674041378947, 32'sd-0.026534514322424704, 32'sd-0.09141288136021362, 32'sd-0.02111710044481535, 32'sd-0.0032159200272251706, 32'sd0.045524908560295195, 32'sd-0.026472709052738904, 32'sd0.06504595652354622, 32'sd0.06309116992887012, 32'sd-0.08458914127745364, 32'sd-0.08435477515212343, 32'sd-0.05513416455903266, 32'sd0.03297306307665123, 32'sd-0.08785842868798131, 32'sd-0.12144428992293603, 32'sd-0.01482978529176855, 32'sd0.05480448074374987, 32'sd0.0009463469412648767, 32'sd-0.07000123472096186, 32'sd0.07346304956198042, 32'sd-0.01935913817385424, 32'sd0.009029422956411615, 32'sd-0.04790088108336434, 32'sd0.11124405796460567, 32'sd0.003921174614259755, 32'sd0.13458132272937623, 32'sd0.04202433264301901, 32'sd0.1890619680714434, 32'sd0.016596842292286928, 32'sd-0.07808464661755105, 32'sd-0.13338033904034036, 32'sd-0.16194378564880468, 32'sd-0.15802858868835354, 32'sd0.01765552527402207, 32'sd0.04422462752964344, 32'sd0.0728759749832712, 32'sd-0.028432227312911933, 32'sd0.03968157110435332, 32'sd0.012847133179112322, 32'sd-0.08237688726085428, 32'sd0.06837266336656492, 32'sd0.009391956784100004, 32'sd-0.0010630913174480027, 32'sd-0.004351252413315976, 32'sd-0.1330381544475429, 32'sd0.04649226610307037, 32'sd0.0022136725524382595, 32'sd-0.03197933210648773, 32'sd0.04348150264369246, 32'sd-0.0770419301368507, 32'sd-0.07218142074897484, 32'sd0.05613476745233639, 32'sd0.030543100658184816, 32'sd0.008238165396683579, 32'sd-0.05937147717839438, 32'sd0.12423088750051478, 32'sd0.012460524448327683, 32'sd-0.17231107766821213, 32'sd-0.09374492479760364, 32'sd0.08113363404984322, 32'sd0.059021607006718546, 32'sd0.01439666144006999, 32'sd0.07463601048312615, 32'sd0.033913112397200885, 32'sd0.057006861807220394, 32'sd0.06529022494513542, 32'sd0.0805840503588192, 32'sd-0.07789488809373275, 32'sd0.008398946819880333, 32'sd-0.09732169954680314, 32'sd-0.06149689898078073, 32'sd-0.1356979412937497, 32'sd0.004569112738271979, 32'sd0.03962213817392719, 32'sd-0.017255427763847017, 32'sd0.01013413561685813, 32'sd-0.011422909335445215, 32'sd0.04060090907141205, 32'sd-0.024203169778857142, 32'sd0.0125577151957548, 32'sd-0.023296796031548717, 32'sd0.023421005082986397, 32'sd0.08244227233059966, 32'sd-0.09851046070820481, 32'sd0.015568681047486056, 32'sd0.021772394565200075, 32'sd0.011428907043202728, 32'sd0.1127684139217824, 32'sd0.005990027343194774, 32'sd0.11519672401003557, 32'sd0.19503298106807376, 32'sd0.04386535823578641, 32'sd0.04801693805176954, 32'sd0.056977901064294206, 32'sd0.04416118598781305, 32'sd-0.058013511563557774, 32'sd-0.06707122510626759, 32'sd-0.08127660123186356, 32'sd-0.1855296515905015, 32'sd-0.05460264352674514, 32'sd-0.0264638263966769, 32'sd-0.0037187051622975214, 32'sd-0.03124597717449228, 32'sd0.051038462617703124, 32'sd0.02118804224226697, 32'sd-0.031051697898214253, 32'sd-0.09591386866871542, 32'sd0.0040878058175592355, 32'sd-0.12309458282089, 32'sd-0.025131713136790985, 32'sd0.04571444871854234, 32'sd-0.04716304424855479, 32'sd0.04259413873874642, 32'sd-0.05366880501970721, 32'sd-0.03756003467048449, 32'sd0.07389784485079773, 32'sd0.10560655764899037, 32'sd0.12709302246653198, 32'sd0.10533815554055286, 32'sd-0.08875248287124969, 32'sd-0.05328616266326727, 32'sd0.07343028204398339, 32'sd0.007539217473258891, 32'sd-0.03729178330512375, 32'sd-0.05115830569177627, 32'sd-0.05897497038476154, 32'sd-0.08079420251279866, 32'sd-0.030369155696323716, 32'sd0.054824772768861864, 32'sd-0.07315869712249881, 32'sd-0.024606340005841075, 32'sd-0.028342788690219927, 32'sd0.019103458950691963, 32'sd-0.0008478578835214602, 32'sd-0.05517509103054172, 32'sd-0.10669100790724163, 32'sd-0.12593563080896839, 32'sd-0.013954145367456258, 32'sd-0.06145171554719042, 32'sd0.03723663565836399, 32'sd0.037787130161867084, 32'sd0.01409455168837901, 32'sd-0.10854345512130459, 32'sd-0.026366532462596855, 32'sd0.038225015553253625, 32'sd0.10134299655511124, 32'sd0.12703683633382865, 32'sd-0.0264597276441568, 32'sd-0.06936723969061105, 32'sd-0.043454660978341754, 32'sd0.03440419267292697, 32'sd0.003084388116148254, 32'sd-0.0028787409491208985, 32'sd-0.09687189619010815, 32'sd-0.08136652306066545, 32'sd-0.04647578518933723, 32'sd0.0012567194240371367, 32'sd-0.0677270768370864, 32'sd-0.09257326231908614, 32'sd0.04599709445867314, 32'sd-0.0020450076427333233, 32'sd-0.02523416620917999, 32'sd-0.048621499175385774, 32'sd-0.0706964792670625, 32'sd-0.06048999521324877, 32'sd-0.10259094030293717, 32'sd0.013550052654633256, 32'sd-0.08622807703548824, 32'sd0.08960310159882676, 32'sd0.02329343928793456, 32'sd-0.016821713872535723, 32'sd0.052765515033964615, 32'sd0.06459188751793234, 32'sd0.008087471384443757, 32'sd0.13104291544910301, 32'sd0.10231923774170808, 32'sd0.08557195220526292, 32'sd0.07541135900891703, 32'sd-0.045165532856393346, 32'sd0.08694194365105601, 32'sd0.02615755705203209, 32'sd-0.03753380373746963, 32'sd0.027627250662649493, 32'sd0.06389346489212627, 32'sd0.1010000100300912, 32'sd0.11427451009991771, 32'sd0.040635086993059996, 32'sd0.01945539570505338, 32'sd-0.03272366293616761, 32'sd-0.04141674358158881, 32'sd-0.07526244366281129, 32'sd-0.07275102936456208, 32'sd-0.07015473255872963, 32'sd-0.05225977010558409, 32'sd-0.011432654736689056, 32'sd0.00511090059301582, 32'sd-0.14918173188961661, 32'sd-0.10032091969638539, 32'sd-0.11159373853185765, 32'sd-0.046501880906299316, 32'sd-0.05656802276555851, 32'sd0.05510266449527916, 32'sd0.09558713900326725, 32'sd-0.05108862072520937, 32'sd0.01619240564708546, 32'sd-0.03024162372444123, 32'sd0.09786705594739682, 32'sd0.05448168336865389, 32'sd0.11084735666618505, 32'sd0.04581493973929185, 32'sd0.08635825635192311, 32'sd0.01650547729170666, 32'sd0.1281594777557537, 32'sd0.1116420577801654, 32'sd0.013996681616774679, 32'sd0.0014089404788840063, 32'sd-1.4514195777378173e-115, 32'sd-0.04113369009273035, 32'sd0.0238510398370762, 32'sd-0.05614544095935738, 32'sd-0.0334379688780179, 32'sd-0.059293902228849206, 32'sd0.004735212383182592, 32'sd0.06194199985105188, 32'sd-0.01982508046382285, 32'sd-0.1440190079309461, 32'sd-0.20088091178532624, 32'sd-0.21985888015255878, 32'sd-0.19356269006324792, 32'sd-0.11599564066294693, 32'sd-0.13585181564413015, 32'sd-0.13968176187913142, 32'sd-0.06455164895197148, 32'sd-0.07607641110594904, 32'sd0.12004954630502547, 32'sd0.2129975205902786, 32'sd0.11923090255163755, 32'sd0.06987777714203156, 32'sd0.11743741664876405, 32'sd0.07104172353367073, 32'sd0.03146708743506174, 32'sd-0.1090223160036208, 32'sd0.0426390311818124, 32'sd0.10546545140290034, 32'sd-0.014473553821480824, 32'sd0.01054510671954984, 32'sd0.039563712807022616, 32'sd0.07042048530856192, 32'sd-0.07594222435646428, 32'sd-0.018262198801816548, 32'sd-0.08169734330116317, 32'sd-0.019479197134994748, 32'sd-0.043744029016451774, 32'sd-0.09435883284356789, 32'sd-0.24860248431077184, 32'sd-0.2721840361378351, 32'sd-0.21079890439625348, 32'sd-0.1986247880477507, 32'sd-0.19559485601372742, 32'sd-0.18125196235568922, 32'sd-0.09199040623552901, 32'sd0.012484004784739463, 32'sd0.12794544955890935, 32'sd0.17713359915615692, 32'sd0.15055386255383485, 32'sd0.19218552018500373, 32'sd-0.021543102025527148, 32'sd-0.04924049703766603, 32'sd-0.10420350416619957, 32'sd-0.05938017533567267, 32'sd0.12930412164828015, 32'sd0.08761568118126384, 32'sd-0.005280869952304285, 32'sd-0.04920354168983839, 32'sd-0.040232614149290434, 32'sd0.07687809655502867, 32'sd-0.0841119442634531, 32'sd0.0495963591757925, 32'sd0.028293908267899147, 32'sd-0.03348909325236208, 32'sd-0.08843956505656532, 32'sd-0.01653092413037717, 32'sd0.027335346523183646, 32'sd-0.024058079937899508, 32'sd-0.062088437828942904, 32'sd-0.1350381462434164, 32'sd-0.1718056599383742, 32'sd-0.1792280294963202, 32'sd-0.08261479600177928, 32'sd-0.11410566383820071, 32'sd0.07342458236823349, 32'sd0.07762544283655722, 32'sd0.13906601605812563, 32'sd0.17538420778764358, 32'sd0.08830472224379743, 32'sd-0.021301711457984655, 32'sd-0.07041015869964112, 32'sd0.048868652522988415, 32'sd0.09590250263276096, 32'sd0.08009473334984428, 32'sd-7.483868186673886e-115, 32'sd0.029732269334591863, 32'sd0.00877351014213967, 32'sd0.035511990557945794, 32'sd-0.01478670939398915, 32'sd-0.05500467149041248, 32'sd-0.018461701131242576, 32'sd-0.03067129495259878, 32'sd-0.029049230594025706, 32'sd-0.026724885488134804, 32'sd0.01980037729090263, 32'sd-0.0297458954906943, 32'sd0.0044127253119420964, 32'sd-0.11876129494293049, 32'sd-0.16517742825282772, 32'sd-0.1354860398995563, 32'sd0.01507417385784231, 32'sd-0.0708102833833676, 32'sd0.10258899364791989, 32'sd0.14758988604605508, 32'sd0.12717710369501128, 32'sd0.1342709886090766, 32'sd0.12146930284696977, 32'sd0.06621591687768144, 32'sd-0.02504915256550803, 32'sd-0.057612708013602534, 32'sd0.06183966568355359, 32'sd0.0010889936041788447, 32'sd0.004200579177829992, 32'sd-0.02420435852178175, 32'sd0.11780475752980654, 32'sd-0.06166625870483514, 32'sd0.009876522020531521, 32'sd-0.03512322667865537, 32'sd-0.03381020289889837, 32'sd0.05613230969724318, 32'sd-0.03488410167912512, 32'sd-0.0016927849062076598, 32'sd0.0716265454208132, 32'sd0.049364105100858036, 32'sd0.07038815748617036, 32'sd0.064287932860484, 32'sd0.020702622252938414, 32'sd-0.00628460003002294, 32'sd0.10393398120579987, 32'sd0.010603653428195858, 32'sd-0.005954037199389498, 32'sd-0.03575438802387262, 32'sd0.07175227526346925, 32'sd0.03692349120109372, 32'sd0.05385497079604361, 32'sd-0.04190557211045563, 32'sd-0.04600060093743583, 32'sd-0.12631414569097194, 32'sd-0.028983482639365978, 32'sd-0.0005746993181098579, 32'sd-0.014733893588576932, 32'sd-0.01808464623272936, 32'sd0.008105193475805909, 32'sd0.05099558398910505, 32'sd0.03636803257466562, 32'sd0.07754434649463969, 32'sd0.03819556200744917, 32'sd-0.012898115656566279, 32'sd0.0715040881343813, 32'sd0.0260690714492402, 32'sd0.10461092159248303, 32'sd0.025136513446043424, 32'sd-0.00418155470982824, 32'sd-0.010494093607173986, 32'sd-0.05626161219322153, 32'sd0.0023987073934768318, 32'sd0.0890085658266689, 32'sd-0.0664945808521404, 32'sd0.0315436815827992, 32'sd0.026234056000292234, 32'sd0.0916485288271415, 32'sd0.006752084724701809, 32'sd0.04305740835007156, 32'sd-0.06493004899733078, 32'sd-0.08365716756394373, 32'sd-0.0023071029983880234, 32'sd0.05324329652598811, 32'sd-0.020956631123570404, 32'sd2.7126945334012194e-124, 32'sd0.01075011827572676, 32'sd-0.03281116430501619, 32'sd0.003407109128838847, 32'sd0.046291251488753266, 32'sd0.04798419534850466, 32'sd-0.025000030398104896, 32'sd0.02026622424216902, 32'sd0.055575645568413594, 32'sd0.012323541854684554, 32'sd-0.03568975298127711, 32'sd0.10078061295642789, 32'sd0.08131394351270443, 32'sd0.05644300657987133, 32'sd0.06313101786856225, 32'sd0.17463251686705183, 32'sd0.06701945672953165, 32'sd-0.018965130439159483, 32'sd-0.03235855841488996, 32'sd0.060309038993915855, 32'sd-0.06466165663458508, 32'sd-0.07381180170914238, 32'sd0.008886460730365428, 32'sd0.011450785009534047, 32'sd0.05876737820027421, 32'sd-0.038017028689017594, 32'sd0.06191264593884068, 32'sd-4.786902217529633e-123, 32'sd1.739457848768853e-125, 32'sd-6.893682854175438e-126, 32'sd0.0925671128656643, 32'sd0.09443894412547689, 32'sd0.056972483237979786, 32'sd0.03651839981133844, 32'sd0.12509102680242035, 32'sd0.07560174548830219, 32'sd-0.03543062466850683, 32'sd0.047847668963565244, 32'sd0.10782988361880953, 32'sd0.11196736171579899, 32'sd0.07895013717790107, 32'sd0.1191397540205779, 32'sd0.05010614770486704, 32'sd0.03496508250456517, 32'sd-0.13619435053739865, 32'sd0.023919755773339185, 32'sd-0.057609557672676746, 32'sd-0.03757624799911262, 32'sd-0.11311694119040176, 32'sd-0.060659594725621456, 32'sd-0.1140644744544618, 32'sd0.04608817818107888, 32'sd0.02491212060605121, 32'sd0.04168994450665587, 32'sd-0.033203725487552245, 32'sd4.819240201747712e-118, 32'sd7.769345082991517e-123, 32'sd2.681897234418458e-118, 32'sd0.0007035479678755488, 32'sd0.00599039535950207, 32'sd0.0230939832485854, 32'sd0.02554530448145316, 32'sd-0.05004318283272237, 32'sd0.025374073918117763, 32'sd0.04155812531329243, 32'sd-0.08074198547643101, 32'sd0.09749583711896455, 32'sd0.07559924852221218, 32'sd0.02990560793500037, 32'sd0.1588840468286339, 32'sd0.02762481793822994, 32'sd-0.0560309642942521, 32'sd-0.02014219234838498, 32'sd-0.044212857224204094, 32'sd-0.2101879959234879, 32'sd-0.11707955794334839, 32'sd-0.09540786106248633, 32'sd-0.19312477997213853, 32'sd-0.13037819874557585, 32'sd-0.023432632150880046, 32'sd-0.16121609638128298, 32'sd-0.0012882166707485147, 32'sd0.01437399565134191, 32'sd1.5523300996904123e-117, 32'sd6.413686845948652e-115, 32'sd-1.3667828762331375e-116, 32'sd-9.79443484210231e-122, 32'sd-0.0035861487837893407, 32'sd-0.08851796191733884, 32'sd0.0453484045653763, 32'sd-0.04428780532135173, 32'sd0.03451548157196717, 32'sd0.024723667596680085, 32'sd0.03398267303080044, 32'sd0.10778653109911068, 32'sd0.04221197296360502, 32'sd0.012073163371370158, 32'sd-0.017517313484235568, 32'sd-0.09262855636526748, 32'sd0.030062043455491242, 32'sd-0.07438760881162423, 32'sd0.1027657364389004, 32'sd0.1344753967629761, 32'sd-0.09801731955715562, 32'sd-0.11281637801077642, 32'sd-0.008949302231247064, 32'sd-0.040522218183201605, 32'sd0.005660462452936233, 32'sd0.0676637838739777, 32'sd-0.0061918284736591795, 32'sd5.729184016659291e-116, 32'sd1.5668702340678783e-115, 32'sd-3.3393337976132675e-123, 32'sd1.5772808262478806e-126, 32'sd-2.7541938817894024e-124, 32'sd1.2431546745694458e-118, 32'sd0.03314367909407499, 32'sd0.06345035412710935, 32'sd-0.04068217922090523, 32'sd-0.01607429565939037, 32'sd-0.03557034788903498, 32'sd-0.029686548474640535, 32'sd-0.0069480131376687074, 32'sd-0.08644317144325328, 32'sd-0.04252363501792293, 32'sd-0.028661962353713967, 32'sd0.04356403445013627, 32'sd-0.0923046555707174, 32'sd-0.0026416663664611934, 32'sd-0.10355080003284337, 32'sd-0.03852430587415493, 32'sd0.05056455180215961, 32'sd-0.07058381494730162, 32'sd0.030176914819339838, 32'sd-0.007870426420624415, 32'sd-0.04160322293747681, 32'sd-1.7199416037390554e-123, 32'sd-7.223451066126255e-115, 32'sd-7.033554953941985e-123, 32'sd-1.0696699835368048e-124},
        '{32'sd1.686590956156469e-125, 32'sd2.807921122874882e-119, 32'sd1.8132032527232373e-123, 32'sd2.2137205104391756e-125, 32'sd6.60827750418556e-115, 32'sd7.284123014519574e-125, 32'sd-1.0654607229484414e-125, 32'sd-2.5112393584931772e-114, 32'sd1.7316656129998587e-119, 32'sd-1.5458962324910911e-118, 32'sd6.309926182510949e-115, 32'sd1.221383327659987e-115, 32'sd0.03912280616215565, 32'sd0.029012406015599023, 32'sd0.011601143343822838, 32'sd0.08659079413937855, 32'sd-3.1851369557541063e-121, 32'sd2.3714114544848932e-122, 32'sd-2.5340384187361147e-120, 32'sd-8.803318139493705e-121, 32'sd-4.9477381573625724e-119, 32'sd-7.751262988182011e-128, 32'sd5.657535888938724e-118, 32'sd1.5077417436829587e-123, 32'sd-1.2850173290439704e-117, 32'sd1.1173906116849979e-123, 32'sd-1.183837373217598e-117, 32'sd5.624037722338918e-125, 32'sd-3.2703013267018587e-121, 32'sd7.651337895187559e-128, 32'sd-1.0427143642571877e-124, 32'sd-1.41527662139528e-121, 32'sd0.042288144353754435, 32'sd-0.02893971200798825, 32'sd-0.03452389303687848, 32'sd-0.0005078260186670739, 32'sd-0.007198984624917558, 32'sd0.021722924412197614, 32'sd-0.02036282154013245, 32'sd-0.06855269629968183, 32'sd-0.054173280768249864, 32'sd-0.04098948974340097, 32'sd0.023562287554857852, 32'sd-0.0015439773508532009, 32'sd0.04692403696430654, 32'sd0.022404615891816502, 32'sd-0.0018028090069692408, 32'sd-0.03491453204280822, 32'sd0.01742247240956252, 32'sd-0.04764372841847636, 32'sd-0.09124469865463114, 32'sd0.05741859011809815, 32'sd1.910855876953198e-127, 32'sd4.5531410041300146e-117, 32'sd3.8522951333346404e-126, 32'sd2.054085881657237e-117, 32'sd2.5256389299824348e-117, 32'sd-5.005612240552601e-118, 32'sd0.003919538914860426, 32'sd0.035631335549780874, 32'sd-0.010375278682552619, 32'sd-0.10362472405871376, 32'sd-0.06989968092123952, 32'sd0.04007932182730984, 32'sd-0.06172045844764074, 32'sd-0.007965761251355934, 32'sd-0.003629114665616872, 32'sd-0.011477225526657392, 32'sd-0.018380047496262805, 32'sd-0.14376435908920532, 32'sd-0.07052787027843141, 32'sd-0.11433958932744671, 32'sd-0.017409125523699356, 32'sd-0.021415838735250596, 32'sd-0.058628941034686834, 32'sd0.0575396204798944, 32'sd0.013843968480720387, 32'sd-0.007107114160850617, 32'sd-0.051006265628656795, 32'sd-0.04485380040304128, 32'sd0.06084672570612125, 32'sd-0.010068387559933542, 32'sd3.478146183909334e-124, 32'sd9.308149690242683e-121, 32'sd-3.991377377585201e-123, 32'sd-1.5688489094631226e-115, 32'sd0.0700147232966069, 32'sd-0.08142750175040098, 32'sd0.0769569244852811, 32'sd5.5013316977707276e-05, 32'sd0.06141291064355639, 32'sd-0.061863765049533746, 32'sd-0.035809513675194256, 32'sd-0.059853924154625204, 32'sd0.10146456782379819, 32'sd-0.058374936106418016, 32'sd0.014010843309040323, 32'sd-0.20537899954833383, 32'sd-0.014293356762753402, 32'sd-0.020062756694682618, 32'sd-0.04166269550015915, 32'sd0.0639315884221735, 32'sd0.17088144759164714, 32'sd-0.03902265925166195, 32'sd0.004592252979125528, 32'sd-0.08939034076520724, 32'sd0.01076823993898443, 32'sd0.015379159162471193, 32'sd-0.032068528785449905, 32'sd0.027094982556447777, 32'sd-0.027031949418182356, 32'sd1.791260825648937e-126, 32'sd-1.201849923209184e-123, 32'sd0.016067641228447303, 32'sd0.043510951254779884, 32'sd-0.016519033311343613, 32'sd-0.15774267666720201, 32'sd-0.08882590364857537, 32'sd0.10051089679130482, 32'sd0.005868782563620318, 32'sd0.008664754616509637, 32'sd-0.06501660851445697, 32'sd0.0068881784810923075, 32'sd-0.02883941850042301, 32'sd-0.13882712892266055, 32'sd-0.053026908502473144, 32'sd-0.1413203771583362, 32'sd0.006484900947651601, 32'sd-0.017127833689443518, 32'sd0.00962523717045751, 32'sd-0.07612021070752269, 32'sd-0.010945397840354684, 32'sd-0.06122843395392809, 32'sd-0.01015543891584995, 32'sd0.03098529543494918, 32'sd-0.05358698926985386, 32'sd-0.07324820478407738, 32'sd0.06140581794228295, 32'sd0.02638412517765473, 32'sd0.06399449869865383, 32'sd-3.1106953092812327e-118, 32'sd0.03296801185691243, 32'sd-0.03292255911069858, 32'sd0.010172976316433525, 32'sd0.022430392180978687, 32'sd-0.021750703434395845, 32'sd0.03399206083575277, 32'sd0.14427956152239116, 32'sd0.11179293513765597, 32'sd-0.02021651747440114, 32'sd0.09309028770108409, 32'sd0.004002339869123693, 32'sd0.08705277038794765, 32'sd0.045351334816259345, 32'sd0.05036288977365477, 32'sd-0.06017620917279386, 32'sd-0.05270966858761881, 32'sd-0.03355039023270475, 32'sd-0.027574297820454865, 32'sd-0.12136337194497392, 32'sd-0.10585794972613992, 32'sd-0.0888898408959809, 32'sd0.006688609094990762, 32'sd-0.04270201266015718, 32'sd0.030063479311508996, 32'sd0.06252211666958503, 32'sd0.01273993825182562, 32'sd-0.07762148899039434, 32'sd8.229971282477344e-122, 32'sd-0.005613779148119941, 32'sd-0.042061833065301056, 32'sd-0.008218859398983088, 32'sd0.03576996919362212, 32'sd0.04178035344300698, 32'sd-0.023361491322818936, 32'sd0.06659736441796191, 32'sd-0.01525834571583092, 32'sd0.15288448325894718, 32'sd0.01082293700043913, 32'sd0.003825992793955867, 32'sd-0.01530044670752228, 32'sd0.12993872994054675, 32'sd0.15457855804056375, 32'sd-0.039647145202074054, 32'sd0.061476502335309505, 32'sd0.08741456707565683, 32'sd0.01054537196226375, 32'sd0.026712845906107417, 32'sd-0.04996958676810446, 32'sd0.08969361781098881, 32'sd0.06890083356803102, 32'sd-0.0497929314617759, 32'sd0.02398897335975779, 32'sd-0.0930317551392441, 32'sd-0.06652384016206274, 32'sd-0.06861401311516024, 32'sd0.0166526501145787, 32'sd-0.02244983893227155, 32'sd0.035655584388291264, 32'sd0.01891980660197559, 32'sd0.024592874380485335, 32'sd-0.09415626648510018, 32'sd0.09214621808593854, 32'sd-0.026793715886579673, 32'sd-0.00505906247008727, 32'sd0.08039556472792143, 32'sd0.010703590019778157, 32'sd0.016209432998641585, 32'sd0.03388691313346535, 32'sd0.2369783056004197, 32'sd0.10472315415281427, 32'sd-0.1422054856647608, 32'sd0.035894706805718574, 32'sd-0.07352757144673873, 32'sd-0.10967783365427294, 32'sd-0.05107209767085662, 32'sd0.12896085464475004, 32'sd-0.026658938763199115, 32'sd-0.09395404387199166, 32'sd0.011015577669351297, 32'sd0.004033200129088612, 32'sd-0.13686481901599126, 32'sd-0.023021657256901668, 32'sd-0.045068135274299724, 32'sd-0.026090741810332403, 32'sd0.07486775374398566, 32'sd0.11918776400707447, 32'sd-0.0660031316315919, 32'sd0.02819473878812579, 32'sd0.0799953941037645, 32'sd0.02192299156947278, 32'sd0.048192474460662646, 32'sd0.07988717539516903, 32'sd0.14336311397835683, 32'sd0.044269004805463155, 32'sd0.1602782353301532, 32'sd0.07729826214684195, 32'sd-0.02150354870089848, 32'sd0.08966794424314839, 32'sd0.07568354283823513, 32'sd-0.06597806360678181, 32'sd-0.006664468701298291, 32'sd-0.0259005556885769, 32'sd-0.042153625588539766, 32'sd0.044174155688453606, 32'sd-0.05254192106138548, 32'sd-0.1141992594199644, 32'sd-0.021097617080026904, 32'sd-0.027553497681949306, 32'sd-0.017483212342490576, 32'sd-0.015949459376555647, 32'sd0.03624130845080228, 32'sd0.03948854268751627, 32'sd0.0976420202843507, 32'sd0.040313285643569945, 32'sd-0.023639254863958285, 32'sd0.05837680871291866, 32'sd0.1260737091758305, 32'sd0.11150794267706399, 32'sd-0.024093053214217636, 32'sd-0.05141019165523631, 32'sd0.025156599214177868, 32'sd0.09372714647229755, 32'sd0.08636005837246961, 32'sd0.08863831351903162, 32'sd-0.015099952395964731, 32'sd0.18541516792253068, 32'sd0.099837559167356, 32'sd0.038049109168539645, 32'sd0.07645243030267784, 32'sd0.057400115319831635, 32'sd-0.10893306796116786, 32'sd-0.01745956420246878, 32'sd-0.08363604064474212, 32'sd0.06574525902380218, 32'sd-0.11361397808185554, 32'sd-0.002960233078641879, 32'sd0.011275481235098412, 32'sd-0.07546358630970458, 32'sd0.036836086475920835, 32'sd0.046147368485056135, 32'sd0.023632458107185984, 32'sd0.07152586812074667, 32'sd-0.06619792831847066, 32'sd0.02927757594964746, 32'sd-0.006165353933152671, 32'sd0.11684285990176248, 32'sd-0.09741037039258689, 32'sd0.12545168525228767, 32'sd-0.046863248589970055, 32'sd0.023158741613892385, 32'sd-0.09185269962763865, 32'sd-0.12183225730047835, 32'sd0.016732141885008697, 32'sd0.13904714936131593, 32'sd0.1586924836050797, 32'sd0.08851173083611917, 32'sd-0.06053818159308145, 32'sd0.0619104501261368, 32'sd-0.05907414228196409, 32'sd-0.044795431459552906, 32'sd-0.11037301477666324, 32'sd0.020605329337968378, 32'sd0.04160198661982984, 32'sd0.05273415001772903, 32'sd0.12002333686486107, 32'sd0.028668202923197314, 32'sd0.011462345240377515, 32'sd0.042493183179648904, 32'sd0.03385524451491292, 32'sd0.0878673173776166, 32'sd0.09928161272092165, 32'sd0.08794381361807176, 32'sd-0.014682785749920177, 32'sd0.08176180139751635, 32'sd0.17073215604446168, 32'sd0.06845004379278635, 32'sd0.05744292008130699, 32'sd-0.031139504578562707, 32'sd0.041419847041523156, 32'sd-0.019001018622486213, 32'sd0.04732967073817793, 32'sd0.11408702949790657, 32'sd0.1322934411712588, 32'sd0.20261623290903416, 32'sd-0.026815004164131066, 32'sd-0.03622395361375255, 32'sd-0.015317319400393617, 32'sd-0.028441848550787345, 32'sd-0.10507113354508464, 32'sd-0.014811081586133264, 32'sd0.029665383295868254, 32'sd-0.011229701125061144, 32'sd0.07331647666600503, 32'sd0.03720972699074013, 32'sd-0.06265665215923027, 32'sd0.005128347461103419, 32'sd0.03743547965681142, 32'sd-0.048283427193623295, 32'sd-0.018552183230737276, 32'sd-0.14195117323234352, 32'sd-0.16599206483065057, 32'sd-0.08222860639903815, 32'sd-0.02710321109758331, 32'sd0.09829916120623985, 32'sd0.00419869151051668, 32'sd-0.03064303777332041, 32'sd-0.08552515133121323, 32'sd-0.028844604979151492, 32'sd0.07257257904205039, 32'sd0.01748818025991186, 32'sd0.225658231988268, 32'sd0.08938861015110051, 32'sd-0.005220184859878409, 32'sd0.029978659838168102, 32'sd-0.11667128726446038, 32'sd-0.1469113549467365, 32'sd-0.1222631640936398, 32'sd-0.12671665585202363, 32'sd-0.0661476569864362, 32'sd-0.08470615734443725, 32'sd0.05339662371248195, 32'sd0.02957471885455587, 32'sd-0.03362355081100162, 32'sd0.007007415916960873, 32'sd-0.070507701739478, 32'sd0.031071882154048287, 32'sd-0.03159865743503312, 32'sd-0.1955022479791065, 32'sd-0.08562937633914286, 32'sd-0.07324185874730689, 32'sd-0.0030666058548554707, 32'sd0.09054745585711686, 32'sd-0.017951569510444243, 32'sd-0.029194198948655506, 32'sd-0.10963645774007785, 32'sd-0.061214636754034095, 32'sd-0.015013545197183212, 32'sd-0.13699786983353693, 32'sd-0.022834871580207593, 32'sd0.12551925889280027, 32'sd0.017997541501126285, 32'sd-0.03408555150848799, 32'sd-0.17766659750318156, 32'sd-0.19561930194937754, 32'sd-0.0926600356839101, 32'sd-0.015531978877459201, 32'sd0.06978817360074255, 32'sd0.01547009926456963, 32'sd0.013599838372707843, 32'sd0.02082360708678503, 32'sd0.006598096997115497, 32'sd-0.021856105240088266, 32'sd-0.02564160999621825, 32'sd0.0375368714543855, 32'sd-0.09830841686606846, 32'sd-0.08820281820944262, 32'sd-0.16182695068652783, 32'sd-0.05196024265847254, 32'sd-0.0628611548039535, 32'sd-0.05692787909733715, 32'sd0.016129652124350715, 32'sd0.08552583716588838, 32'sd0.03476120987216325, 32'sd-0.01104100041065512, 32'sd-0.14721860273945905, 32'sd-0.05175801728545287, 32'sd-0.04425537492334462, 32'sd0.029400515290029634, 32'sd0.08219263876684586, 32'sd-0.03702871477887495, 32'sd-0.13983251761135582, 32'sd-0.09186939050712033, 32'sd-0.009512671552949393, 32'sd-0.05894780871998037, 32'sd-0.02208009670927555, 32'sd-0.07776687871591474, 32'sd-0.032590923774153756, 32'sd0.031137622438116328, 32'sd-0.05760843286350163, 32'sd-0.025438860709758253, 32'sd0.04733133437997303, 32'sd-0.00526816762000667, 32'sd-0.07544512931487954, 32'sd-0.040474723368223844, 32'sd-0.20201045182229171, 32'sd-0.24013761429197839, 32'sd-0.041336089073404914, 32'sd-0.06384139005239582, 32'sd0.0958305918468672, 32'sd0.16824926436071197, 32'sd0.1341199308050854, 32'sd0.019570585512477454, 32'sd-0.09685490254556499, 32'sd0.05012836636270554, 32'sd0.08387839441723413, 32'sd0.05774650042601675, 32'sd0.21016819824245303, 32'sd0.04786721696046146, 32'sd-0.13388614301047624, 32'sd0.04396181331060223, 32'sd0.03352513496402884, 32'sd0.08003892152222081, 32'sd0.015921369043165837, 32'sd0.007109248931278236, 32'sd-0.06692891636900324, 32'sd-0.027677273203096077, 32'sd-0.011461080437072653, 32'sd0.006083191707761094, 32'sd-0.04732547091788707, 32'sd0.02241230930025702, 32'sd-0.12148859512311597, 32'sd-0.03453712772018098, 32'sd-0.11191873405042177, 32'sd-0.09149930870003589, 32'sd0.07948682973978542, 32'sd0.10577123993518074, 32'sd0.115467381615079, 32'sd0.06473828261475822, 32'sd0.13949562367299098, 32'sd0.14033120166856872, 32'sd0.1342114623384948, 32'sd0.03802911171755873, 32'sd0.20281793735175968, 32'sd0.17659247057613697, 32'sd0.18251996723280872, 32'sd0.011938273464789996, 32'sd0.00558752998365181, 32'sd0.02760371877283997, 32'sd0.06271798992085913, 32'sd0.03913887831464929, 32'sd0.07977053480342798, 32'sd-0.12767028459035903, 32'sd-0.07030041984748348, 32'sd0.03888616132655312, 32'sd0.009406973237495987, 32'sd-1.5171280158531485e-117, 32'sd-0.02652941412289676, 32'sd-0.014916695926380124, 32'sd-0.06795075790912773, 32'sd-0.009519405166005798, 32'sd-0.0245616940379414, 32'sd0.0875467826603357, 32'sd0.11639764001301364, 32'sd0.07601132681578515, 32'sd0.012844375764675217, 32'sd0.027751559691291335, 32'sd0.008129956682093785, 32'sd0.04749345433159716, 32'sd-0.026187722438063207, 32'sd0.024918053891651495, 32'sd0.15019579806921962, 32'sd0.013939253892037755, 32'sd0.03527777785966089, 32'sd0.020290364852662952, 32'sd-0.09047525405587588, 32'sd0.04444619962804077, 32'sd0.12519148847442158, 32'sd0.128325058696602, 32'sd-0.03454254380055738, 32'sd0.04616773484584927, 32'sd0.007110508243377993, 32'sd0.014570647622592622, 32'sd0.008958643093259226, 32'sd-0.04050254453363865, 32'sd0.018187162547948593, 32'sd0.05390294929235075, 32'sd-0.0893078654871755, 32'sd-0.07974945625433373, 32'sd-0.05817048058755251, 32'sd-0.11390214147728314, 32'sd-0.007198061398156981, 32'sd-0.09382350491171815, 32'sd-0.05349623714493668, 32'sd-0.05605978253951183, 32'sd-0.10614750315731512, 32'sd-0.11112856329504406, 32'sd0.019079102219988583, 32'sd0.04732245687940593, 32'sd0.11946642834774154, 32'sd0.046747748149852615, 32'sd0.07610569192483624, 32'sd-0.18195233574321398, 32'sd-0.02513480484222889, 32'sd0.07267866131258686, 32'sd-0.05741128018665008, 32'sd-0.05092665127937187, 32'sd-0.03898631408616148, 32'sd-0.026128094761145863, 32'sd-0.09503094363675321, 32'sd0.10027181582354575, 32'sd-0.08390299653602995, 32'sd0.05368413198896206, 32'sd-0.005159793928213398, 32'sd-0.004630158671375467, 32'sd-0.006723812806911039, 32'sd-0.07547429814905321, 32'sd0.016517113584747924, 32'sd-0.21682282206865205, 32'sd-0.18345616228930148, 32'sd-0.20981491254334153, 32'sd-0.16167664831515535, 32'sd-0.24656532935770709, 32'sd-0.21857522915390518, 32'sd-0.08962266283002489, 32'sd-0.02003715200131747, 32'sd-0.06002088606301052, 32'sd0.024318219024356942, 32'sd-0.09933027825927801, 32'sd-0.08594351325639804, 32'sd-0.10992528196388343, 32'sd-0.05952934314530859, 32'sd-0.056285754560255315, 32'sd-0.04010998209666433, 32'sd-0.06971362010817461, 32'sd0.03532518400576711, 32'sd-0.057959425602628546, 32'sd-0.09556325241527125, 32'sd-0.07409940181824617, 32'sd-0.005171747028082073, 32'sd5.9614609857574726e-120, 32'sd0.0022399237942111135, 32'sd-0.05880623251211568, 32'sd-0.04956165897800477, 32'sd-0.06190809174371483, 32'sd-0.19812121325122325, 32'sd-0.23622549690844083, 32'sd-0.10542587501614992, 32'sd-0.17978996919997858, 32'sd-0.11740947495594725, 32'sd-0.15545122299157857, 32'sd-0.1289593999121651, 32'sd-0.02419146931240366, 32'sd0.06175120185187996, 32'sd-0.10641102805630169, 32'sd-0.14502832069285548, 32'sd-0.14582313999150667, 32'sd-0.21827202928676728, 32'sd-0.12030602481590821, 32'sd-0.18237855926300608, 32'sd-0.01774120448332438, 32'sd-0.039262558309550125, 32'sd0.021403966713618036, 32'sd-0.011400040357415046, 32'sd0.00215465261393814, 32'sd-0.04777884376785641, 32'sd-0.12091467676255595, 32'sd0.01101554712758631, 32'sd0.02241729244756406, 32'sd0.02398903248576039, 32'sd-0.07264357634400485, 32'sd0.04457377644371344, 32'sd0.11355628166891539, 32'sd-0.05726814737158075, 32'sd-0.192078293323365, 32'sd-0.11213488088779101, 32'sd-0.14246883650325975, 32'sd0.03244980075989636, 32'sd-0.07652943775270596, 32'sd-0.0329223613685489, 32'sd0.10960912961036286, 32'sd-0.04312601319263512, 32'sd-0.11876154642878446, 32'sd-0.08782472259006276, 32'sd-0.012692695139926925, 32'sd-0.09718691021894009, 32'sd-0.3073900072122863, 32'sd-0.11878681448802456, 32'sd-0.13658518674381734, 32'sd-0.06816515068716841, 32'sd0.08985356463916867, 32'sd0.03533805014384137, 32'sd-0.01186678853786698, 32'sd-0.016117692684494662, 32'sd-0.012199721042516007, 32'sd0.03483707068231454, 32'sd-0.009969963301773832, 32'sd0.03962696473410033, 32'sd0.010768210019708596, 32'sd-0.03070357801304206, 32'sd0.00463085443223918, 32'sd0.046489623345530466, 32'sd0.042745190117266164, 32'sd-0.04752575147351338, 32'sd0.014688072959241481, 32'sd-0.012748635783931551, 32'sd0.20370190708229954, 32'sd0.06618521734705753, 32'sd0.09493870427551705, 32'sd-0.12130056799172452, 32'sd-0.0742994915366572, 32'sd-0.0090961419092172, 32'sd-0.0617647714938161, 32'sd-0.08001949862240856, 32'sd-0.17632537095555353, 32'sd-0.10166613426464487, 32'sd-0.15414206336112968, 32'sd-0.1329657858314131, 32'sd0.07383465010190363, 32'sd-0.09101055543044911, 32'sd-0.020081448507050063, 32'sd0.05437485676206422, 32'sd-0.007179609452625646, 32'sd-0.04327505777080213, 32'sd2.20450394171646e-126, 32'sd0.07477323939773899, 32'sd-0.03645693603050657, 32'sd0.07892058018009841, 32'sd-0.03890662385498558, 32'sd0.0148008187303121, 32'sd0.09043534830107057, 32'sd0.06007594788831292, 32'sd0.03626632961513397, 32'sd0.07077705491684025, 32'sd0.03491663538179206, 32'sd0.047030715529305836, 32'sd0.03113566515216848, 32'sd-0.013733268315815866, 32'sd0.007746728971156467, 32'sd0.013511874500155965, 32'sd0.011210624708721919, 32'sd0.04954267453642649, 32'sd-0.07661785912767824, 32'sd-0.10790066508776058, 32'sd-0.08716081290811364, 32'sd0.007317975089790805, 32'sd-0.02604543434830363, 32'sd0.014401928145401127, 32'sd0.04568091088097445, 32'sd-0.013584305236337432, 32'sd-0.07151070513797701, 32'sd3.2227204317448834e-120, 32'sd7.459079557064881e-117, 32'sd2.515688003881953e-123, 32'sd-0.022651964318320016, 32'sd0.0246988500108019, 32'sd-0.07131958322285066, 32'sd0.06890573549130016, 32'sd0.07357086038025955, 32'sd0.0441444638883937, 32'sd0.07122781016134727, 32'sd-0.021263090556783687, 32'sd0.08638352679393657, 32'sd0.013459276021383002, 32'sd0.0183106361887169, 32'sd-0.045697443280180924, 32'sd0.002364293280636885, 32'sd-0.07776601224147062, 32'sd-0.0038250895818094815, 32'sd-0.05453254667254075, 32'sd-0.06501143702854488, 32'sd0.05401699852620303, 32'sd0.010437615884607593, 32'sd0.019782713914621972, 32'sd0.07424733469341112, 32'sd0.027666016420299186, 32'sd0.022777273978386296, 32'sd-0.005007094349080614, 32'sd0.02969032299721296, 32'sd3.126764514070771e-116, 32'sd-5.456418220633707e-123, 32'sd-2.7432337815204282e-123, 32'sd0.08526016947245209, 32'sd0.05504219370851781, 32'sd-0.026121089376055166, 32'sd0.08226993976972256, 32'sd-0.004284277178850918, 32'sd0.00877315386003827, 32'sd-0.01007353382910201, 32'sd0.016418849164451323, 32'sd0.06770278753494367, 32'sd-0.0677172362309219, 32'sd-0.02519611865313821, 32'sd-0.1106003167264104, 32'sd-0.13025899121906456, 32'sd-0.05002324536001252, 32'sd-0.05611391312190681, 32'sd0.060350896841790846, 32'sd-0.06298209696615374, 32'sd-0.02758523015811365, 32'sd-0.04533900407385617, 32'sd-0.006404910274985453, 32'sd-0.07352416137688648, 32'sd-0.01885763347497447, 32'sd0.019548772425990985, 32'sd0.048576448924277545, 32'sd-0.026426053172814767, 32'sd-9.286189833041321e-119, 32'sd-8.130706609875604e-117, 32'sd-3.287323623863847e-122, 32'sd-4.342576485654801e-126, 32'sd-0.01131171585623437, 32'sd0.005395010462922497, 32'sd-0.007053627407744264, 32'sd-0.05431623680395106, 32'sd0.01217100574322463, 32'sd0.060212599966192715, 32'sd0.03611015765998229, 32'sd0.1694705070911401, 32'sd0.05794205504479176, 32'sd0.0625312728761159, 32'sd0.030014922795825343, 32'sd0.016261281177594154, 32'sd0.02438091149392932, 32'sd-0.02479040048613641, 32'sd0.044639190962870556, 32'sd-0.0016304227117655242, 32'sd0.06481135756903039, 32'sd0.009667846422711927, 32'sd-0.023793497131103274, 32'sd0.04265039765141233, 32'sd0.06791774929615156, 32'sd0.0657148319621064, 32'sd0.051306178952258426, 32'sd-8.779782977731169e-126, 32'sd2.4044367108336174e-126, 32'sd-6.521382467793588e-119, 32'sd-9.926600726468912e-116, 32'sd8.798706490340451e-121, 32'sd-1.2006584309456081e-119, 32'sd0.061868533951340725, 32'sd-0.0022317051405861855, 32'sd-0.0011117584511992854, 32'sd0.08182290617261392, 32'sd-0.08209374028990292, 32'sd-0.025277105844884556, 32'sd0.05663970596015449, 32'sd-0.016110902891668957, 32'sd-0.06769320230183315, 32'sd0.03742860918578183, 32'sd0.12050231843752147, 32'sd0.050681551338173356, 32'sd0.13860180554423068, 32'sd0.056746776318573465, 32'sd0.047055925973398104, 32'sd0.05016902599819213, 32'sd-0.025062472833745464, 32'sd0.08682376819611652, 32'sd0.10068281676469888, 32'sd0.11877148226422639, 32'sd7.930232490862635e-119, 32'sd-7.523753387045692e-122, 32'sd1.353880688218552e-126, 32'sd4.837964699935177e-126},
        '{32'sd-4.189831296795278e-123, 32'sd7.642879618939195e-122, 32'sd2.4964448117682036e-126, 32'sd-9.610797594034445e-120, 32'sd1.21947698062975e-117, 32'sd-1.5872794110447918e-117, 32'sd2.9501272926240037e-121, 32'sd-2.570487270987345e-116, 32'sd8.343470537652296e-117, 32'sd-7.194086319366897e-125, 32'sd-7.606165772219849e-117, 32'sd-2.0911021672957146e-116, 32'sd-0.03112711634442731, 32'sd0.036826571643518664, 32'sd0.09758006668981115, 32'sd-0.013200635595462787, 32'sd1.190721739465101e-121, 32'sd-1.5910573630791697e-126, 32'sd8.073218923082579e-125, 32'sd1.9928924360260443e-121, 32'sd3.392248977798446e-118, 32'sd-2.4665376375888977e-125, 32'sd3.254791251041657e-125, 32'sd2.194183935883895e-124, 32'sd7.558289718577703e-115, 32'sd-1.69304639045973e-126, 32'sd-1.5712732252659041e-124, 32'sd-3.0909851397172705e-129, 32'sd-8.579612287884585e-120, 32'sd8.621359421883415e-117, 32'sd1.035550893411382e-122, 32'sd3.199786054901723e-124, 32'sd-0.012770057351253306, 32'sd0.06017773082797674, 32'sd-0.00623543911472592, 32'sd0.004123176365755373, 32'sd0.01011854008634903, 32'sd0.05649127416601607, 32'sd-0.08451664322977563, 32'sd0.01564317315785366, 32'sd-0.03165793184904436, 32'sd-0.004675406095266324, 32'sd0.03670215851749224, 32'sd0.053985260050311, 32'sd0.03341276672943909, 32'sd0.04463548075782956, 32'sd-0.03870809605987158, 32'sd-0.012865266801936991, 32'sd0.05485052767488876, 32'sd-0.03488743213022209, 32'sd0.024408455331081796, 32'sd0.0006726246808409341, 32'sd-1.98107329465328e-117, 32'sd1.1653990371136068e-118, 32'sd5.345001714757295e-117, 32'sd4.847447190318585e-118, 32'sd3.452697640963806e-125, 32'sd-6.164594780785119e-127, 32'sd0.056177295648971, 32'sd0.00407156548965251, 32'sd0.06318353608457637, 32'sd0.033683853728318544, 32'sd0.006388387824167213, 32'sd-0.02682732326191655, 32'sd-0.04155028324240732, 32'sd-0.046912711514470955, 32'sd0.0586763927237864, 32'sd0.03928995786512515, 32'sd-0.04500077107231011, 32'sd-0.17658081708185744, 32'sd0.051871271266026635, 32'sd0.022931458719531565, 32'sd0.13110239908984397, 32'sd0.11869900427151954, 32'sd0.019130776520665287, 32'sd0.007242274052436795, 32'sd-0.09676548478857466, 32'sd0.023305442741286174, 32'sd0.033083713557832246, 32'sd0.06755409383466399, 32'sd-0.061003179950971424, 32'sd0.05333970484137965, 32'sd1.6930350706344673e-122, 32'sd-4.868686933585126e-123, 32'sd7.1630572076687685e-115, 32'sd2.375608954718512e-122, 32'sd0.0713952138839464, 32'sd-0.03484609781886807, 32'sd-0.029507595822049336, 32'sd-0.02974723785343446, 32'sd0.08120424472119403, 32'sd0.055663280783009264, 32'sd0.009146950717270043, 32'sd0.00016284320194386742, 32'sd0.06134451090217473, 32'sd0.0123694590408937, 32'sd-0.0187438885130815, 32'sd-0.14034510419796598, 32'sd-0.10012975343281594, 32'sd-0.09391263947233267, 32'sd-0.03269628668872653, 32'sd0.056297315736789554, 32'sd0.04325792368226786, 32'sd0.03110870541741811, 32'sd0.022107214913666098, 32'sd0.11255901512696408, 32'sd-0.015963211314127864, 32'sd0.03457575642044634, 32'sd-0.07233522205069197, 32'sd-0.03024470246875811, 32'sd0.023512129383385854, 32'sd-3.0247389233018927e-122, 32'sd3.204139344183831e-116, 32'sd0.01529470573761734, 32'sd-0.015469572964084143, 32'sd0.08189879733959446, 32'sd0.03676788664382392, 32'sd-0.09672088730477282, 32'sd-0.12013055009447193, 32'sd-0.09750078170243229, 32'sd-0.07954204959150357, 32'sd-0.10225457369796653, 32'sd-0.029122489858601275, 32'sd0.10793862090638506, 32'sd0.020100448182092178, 32'sd-0.012661871112430017, 32'sd-0.12514774715109378, 32'sd-0.08251591419019155, 32'sd-0.024569112676959732, 32'sd-0.0892877678181769, 32'sd-0.07518246399997774, 32'sd-0.04591663782448556, 32'sd0.06760147781828796, 32'sd0.12066996929086658, 32'sd-0.005377466288562989, 32'sd-0.013159766049237456, 32'sd-0.052970682647020643, 32'sd-0.07396045569940196, 32'sd-0.04460598527537093, 32'sd-0.005416663206413233, 32'sd2.91280509236036e-118, 32'sd0.061116897904256694, 32'sd0.025355794327451456, 32'sd0.06861971653319188, 32'sd0.026370970913811576, 32'sd0.060738029972920486, 32'sd0.09205915978131399, 32'sd-0.01538522340006965, 32'sd0.10576857296369536, 32'sd0.016905108637830457, 32'sd-0.03238856137420652, 32'sd0.020717932784844798, 32'sd-0.13427714930941448, 32'sd-0.14343821839402973, 32'sd-0.15908057192951125, 32'sd-0.15638773985446472, 32'sd-0.04278976311351623, 32'sd-0.03585939943198209, 32'sd-0.047835845358740046, 32'sd0.0029836201306170465, 32'sd-0.009095261707256433, 32'sd0.06172437102139375, 32'sd0.014253571403457533, 32'sd-0.07481640404111146, 32'sd-0.021401713153178584, 32'sd-0.04093658209672267, 32'sd-0.03925402210804629, 32'sd0.038791960748505654, 32'sd-3.660936238778565e-119, 32'sd-0.008591824479268893, 32'sd-0.019202356346780233, 32'sd-0.04377153471192883, 32'sd0.1267060592167288, 32'sd0.111294981004959, 32'sd0.07184126112418017, 32'sd0.04829331226706584, 32'sd-0.0995450362013294, 32'sd0.05123930259864923, 32'sd0.10074254715044308, 32'sd-0.08163347164566273, 32'sd0.1261305478742276, 32'sd0.05765169296449556, 32'sd-0.06426850421862171, 32'sd-0.03674996374340258, 32'sd0.033090133538705845, 32'sd0.1294701294133429, 32'sd0.05050593583553315, 32'sd0.05645481468347615, 32'sd-0.08386173234371222, 32'sd0.11587018641199306, 32'sd0.014404602180316722, 32'sd-0.04537120944661925, 32'sd-0.08659308480744277, 32'sd-0.05099370502536352, 32'sd-0.06459872318302758, 32'sd0.040596288824208744, 32'sd0.03455429324304576, 32'sd-0.022506463287193478, 32'sd0.061827005856369334, 32'sd-0.05759675971809272, 32'sd0.04995598034061302, 32'sd-0.05548280802467932, 32'sd0.07859076026476783, 32'sd0.05374527377241951, 32'sd-0.0058371084322625414, 32'sd0.12913158593643445, 32'sd0.07820653489734851, 32'sd0.06084239349222341, 32'sd0.09793230961493943, 32'sd0.09350961262886251, 32'sd-0.044069376288998416, 32'sd-0.05393822908689797, 32'sd0.1264708857818902, 32'sd0.010055432106345855, 32'sd0.09461930400622137, 32'sd0.07085035401184955, 32'sd0.10332056837951745, 32'sd-0.00048013609217187515, 32'sd0.08707275680773365, 32'sd-0.001548427693122576, 32'sd0.04066696021820939, 32'sd0.05787994999817097, 32'sd-0.0664395441374647, 32'sd-0.09378820709182258, 32'sd-0.031088330339499, 32'sd-0.018269378758412145, 32'sd0.0662661392557167, 32'sd0.035431292916663436, 32'sd-0.048108266238136, 32'sd-0.03246946953090151, 32'sd-0.058715178361586136, 32'sd0.05766412410126574, 32'sd0.03981788921518928, 32'sd0.1951100379692418, 32'sd0.14499875842841856, 32'sd0.1259652734863033, 32'sd-0.017755817713299257, 32'sd0.05040654534452336, 32'sd-0.01693731465204071, 32'sd0.12203092935246937, 32'sd0.05135492189305425, 32'sd0.10575609452435128, 32'sd0.09235164052059429, 32'sd0.068127731746231, 32'sd-0.03439614226917827, 32'sd-0.04403199545784715, 32'sd0.10666529582893287, 32'sd-0.08033123915938904, 32'sd0.05122729521628015, 32'sd-0.044854113147611424, 32'sd-0.09992212323811633, 32'sd0.00016453540104273363, 32'sd0.05800083867365738, 32'sd0.06790366940346217, 32'sd-0.06012727611969694, 32'sd-0.042445449951643295, 32'sd-0.03772852598377006, 32'sd0.004957522880008076, 32'sd0.0839581000518137, 32'sd0.02342644275223271, 32'sd0.056665575062650866, 32'sd0.055844319724466414, 32'sd0.08778911996546934, 32'sd0.030374935309581425, 32'sd0.04574843311606891, 32'sd0.09341049571247685, 32'sd0.06763210595568364, 32'sd-0.029548642529052403, 32'sd0.010183797050277053, 32'sd0.00903525669375439, 32'sd-0.005972089715650387, 32'sd-0.10446108329481406, 32'sd-0.037555254845525986, 32'sd0.05256254187809881, 32'sd-0.015345113960637714, 32'sd-0.00974069605331107, 32'sd-0.027517120257055723, 32'sd-0.17615828897770053, 32'sd-0.005328924343701962, 32'sd-0.011503257152038171, 32'sd0.08143678101547745, 32'sd-0.055381144296498284, 32'sd0.02999040086873854, 32'sd-0.15209697164882285, 32'sd-0.03946398448739579, 32'sd0.07817957080548014, 32'sd0.028645753868868945, 32'sd0.0028048718473257604, 32'sd-0.04184627396283628, 32'sd-0.03459123147316159, 32'sd0.06367130004033543, 32'sd0.11252546447906728, 32'sd0.0019901684680980226, 32'sd0.061486261521139465, 32'sd-0.09015005190915103, 32'sd-0.10082936213393784, 32'sd-0.06628915431914294, 32'sd0.034802099795073774, 32'sd0.12874757670239123, 32'sd0.07459167293237369, 32'sd-0.01020190401587246, 32'sd0.02402024139585188, 32'sd-0.044035058989954814, 32'sd0.03906158303028179, 32'sd0.04840611076518478, 32'sd-0.12409443842798956, 32'sd-0.0006395244298451274, 32'sd0.012198914727972649, 32'sd0.0417224890936997, 32'sd-0.0031072699757051844, 32'sd-0.11404323018536518, 32'sd-0.016112060985003777, 32'sd-0.009844074052477543, 32'sd-0.00023290585506931176, 32'sd0.04502935105171151, 32'sd0.11670405538333178, 32'sd-0.021862199130188626, 32'sd0.11526157081979262, 32'sd0.03865977808759897, 32'sd0.13732847528287107, 32'sd0.0785672049162083, 32'sd-0.01595136691345179, 32'sd0.0019010978242779786, 32'sd0.007877062377013133, 32'sd-0.05144921505774521, 32'sd0.12849746619785818, 32'sd0.19964183200967675, 32'sd-0.030617701978587146, 32'sd0.05474425628086433, 32'sd-0.07715118330731725, 32'sd-0.0441171211685346, 32'sd0.031693436377247794, 32'sd0.04503173943745411, 32'sd-0.011182644894764083, 32'sd0.039537592617325305, 32'sd0.008895162371203445, 32'sd-0.0023571192312952546, 32'sd0.02065645970365958, 32'sd-0.013712264056809967, 32'sd-0.020951362748009603, 32'sd-0.1297875501381382, 32'sd-0.03590997776049656, 32'sd0.03136543604327225, 32'sd-0.05429999647550157, 32'sd0.03980732080915452, 32'sd-0.03538373029094236, 32'sd0.06131238260690509, 32'sd0.03221941990194412, 32'sd-0.07601603235537296, 32'sd-0.10713017986003391, 32'sd-0.17161862140594214, 32'sd0.09659566852726824, 32'sd0.14749988743286976, 32'sd0.08902766396859144, 32'sd0.03916426396203872, 32'sd-0.05673392271914866, 32'sd-0.04153150490143135, 32'sd0.020062894163582607, 32'sd-0.050171157528706115, 32'sd-0.13117841680053954, 32'sd0.06807696045616952, 32'sd0.06649660746335805, 32'sd-0.06337080022800007, 32'sd0.05574913389446082, 32'sd0.013518454298636132, 32'sd-0.004096967568805333, 32'sd0.052707740153384496, 32'sd-0.14469568704914096, 32'sd-0.08260055833504172, 32'sd-0.04192379950112126, 32'sd-0.012734683281629858, 32'sd0.007351111097977415, 32'sd0.061108176375603604, 32'sd-0.06707511372691544, 32'sd0.07561624444611821, 32'sd0.05717046125049122, 32'sd-0.08844480510239397, 32'sd-0.2189526714101159, 32'sd-0.1386130652792065, 32'sd0.012620958064068972, 32'sd0.1352734105584302, 32'sd-0.03562826137780327, 32'sd-0.01838252163452493, 32'sd-0.14438798531875174, 32'sd-0.09439862492618524, 32'sd0.022250940333581888, 32'sd-0.005888696898688684, 32'sd-0.03534207773795308, 32'sd-0.11037658868464786, 32'sd-0.10637969365943835, 32'sd-0.060116566355539684, 32'sd0.08552588156369585, 32'sd0.0111300307500548, 32'sd0.013782294570924327, 32'sd-0.004529820089432241, 32'sd-0.011597822943604633, 32'sd-0.02626857053769573, 32'sd-0.0829440389993447, 32'sd-0.11335290362712751, 32'sd0.015886947370546856, 32'sd0.019550416955727686, 32'sd-0.005403820233844569, 32'sd0.03607495354833992, 32'sd-0.03633418805400732, 32'sd-0.12251212702129695, 32'sd-0.11294769886587705, 32'sd-0.04417654699929127, 32'sd-0.07756525042307513, 32'sd0.07248974452755512, 32'sd0.08404792571657853, 32'sd-0.03859972561831026, 32'sd-0.04721610271048784, 32'sd0.05260205797402153, 32'sd-0.11076437949098515, 32'sd-0.11520809639154408, 32'sd-0.1897131961478991, 32'sd-0.10405908233436281, 32'sd0.07804738390351476, 32'sd-0.010564185445384415, 32'sd0.04107607000030059, 32'sd-0.031961580064126596, 32'sd0.028751691437074237, 32'sd-0.015478614920466344, 32'sd-0.05367704900455065, 32'sd-0.08374470601767638, 32'sd-0.12484444008812616, 32'sd-0.06426280972329527, 32'sd0.03346671520624051, 32'sd-0.02152771330545857, 32'sd-0.061200086596479075, 32'sd0.005289706035633775, 32'sd-0.04113958274260461, 32'sd-0.11410271162696678, 32'sd-0.14736997320417586, 32'sd-0.06902686877278691, 32'sd-0.07558099598253067, 32'sd0.07722970562667718, 32'sd0.10162895575536694, 32'sd0.06714586168364611, 32'sd-0.15353928031766065, 32'sd0.020228671963994523, 32'sd-0.050886019138397014, 32'sd-0.08474260244440628, 32'sd-0.10429059117454524, 32'sd0.028220681009087895, 32'sd0.07056684629203643, 32'sd0.0883242485898382, 32'sd-0.037033984615639996, 32'sd0.031978421469400865, 32'sd0.03514069357659768, 32'sd0.08540351613459901, 32'sd-0.03903647340571441, 32'sd0.04382943413760592, 32'sd-0.005293427938466634, 32'sd0.015650522131532434, 32'sd0.17235078439597826, 32'sd0.12541306172936387, 32'sd-0.03188946886148099, 32'sd0.11244601878028643, 32'sd-0.05135754568963192, 32'sd-0.02589433122872112, 32'sd-0.03793303523852949, 32'sd-0.0075645117063920094, 32'sd0.059864780962044936, 32'sd0.16920938126436139, 32'sd0.08300318710339308, 32'sd-0.09028935314447765, 32'sd-0.036400413553688164, 32'sd0.04198228071425097, 32'sd0.012648419476793456, 32'sd0.037381280332337695, 32'sd0.007887558909198959, 32'sd0.03228516948804903, 32'sd-0.0408535705990432, 32'sd-0.04595315094502754, 32'sd0.06617535720893773, 32'sd5.349780643159386e-115, 32'sd0.02201851909995213, 32'sd-0.024421567688788556, 32'sd-0.018993646768172955, 32'sd0.006095777920131362, 32'sd0.10202719650447177, 32'sd0.014509932766758122, 32'sd0.11373806550788967, 32'sd0.06366733991220111, 32'sd-0.03811834844262101, 32'sd0.013923615391078975, 32'sd0.018570589114514955, 32'sd-0.13390823482819728, 32'sd-0.144925915520868, 32'sd0.0010087015356322465, 32'sd0.15632680447076677, 32'sd0.0827971758515834, 32'sd0.01977909843594366, 32'sd0.04389674943264192, 32'sd-0.001255662276886219, 32'sd0.11805713129836674, 32'sd0.18154082071319935, 32'sd0.21175464683912817, 32'sd0.06257915361410826, 32'sd-0.0066652834528590525, 32'sd0.05068065838797476, 32'sd0.05823477042371322, 32'sd0.035479774596612404, 32'sd0.05329369008754483, 32'sd-0.0011937757218824538, 32'sd0.003196794048626148, 32'sd-0.11172305408896742, 32'sd0.13711257700022525, 32'sd-0.0388390324155013, 32'sd0.0011817517060290566, 32'sd-0.03286116454976358, 32'sd0.0008396338142155777, 32'sd-0.09751287047794957, 32'sd-0.11602421500573437, 32'sd-0.20859339550716044, 32'sd-0.1715621446969705, 32'sd-0.1064209116824612, 32'sd-0.01637992755103949, 32'sd0.015821621039437447, 32'sd0.10394890880029939, 32'sd0.041524218175414296, 32'sd0.02435755051361664, 32'sd-0.07066943946971736, 32'sd-0.023220904090659664, 32'sd0.052204510516776964, 32'sd0.17105866056984476, 32'sd0.0827744917971755, 32'sd0.05791412381935828, 32'sd0.10506474402374771, 32'sd0.07671418232043489, 32'sd0.05569121224893786, 32'sd0.03604728972954593, 32'sd-0.03716408721648792, 32'sd-0.08154471405283387, 32'sd0.0568864278259407, 32'sd0.08555761946036762, 32'sd0.018637269321658143, 32'sd-0.041459137691270624, 32'sd-0.02782534016251492, 32'sd-0.09420626208713825, 32'sd-0.09904349116318643, 32'sd-0.1125002068343555, 32'sd-0.15152929314302277, 32'sd-0.17789292160235318, 32'sd-0.09258622645913506, 32'sd0.050935901810069205, 32'sd-0.09441039728779385, 32'sd-0.0967521783588943, 32'sd-0.08646123778301991, 32'sd-0.09422095499768221, 32'sd0.005053300817125552, 32'sd0.05110283508421303, 32'sd0.13886739873626633, 32'sd0.16656755243170035, 32'sd0.16089349040001605, 32'sd0.016318844893298046, 32'sd0.024307672490379413, 32'sd0.04608941024556523, 32'sd0.04208596921187589, 32'sd8.519783830906445e-117, 32'sd-0.05150132097715579, 32'sd-0.05697496255886129, 32'sd0.033684766863949896, 32'sd0.13796405427292507, 32'sd0.058197480448082144, 32'sd-0.07215299202043246, 32'sd-0.017145367737629497, 32'sd-0.046141079348251936, 32'sd-0.1014893482568817, 32'sd-0.13684185537808694, 32'sd-0.06422935672960225, 32'sd-0.018795392292994987, 32'sd-0.08036076945287048, 32'sd-0.0075555973404468745, 32'sd-0.045688752728468875, 32'sd-0.06716939755498647, 32'sd-0.09362062499147533, 32'sd-0.1512484197886483, 32'sd-0.05621848031671012, 32'sd-0.06667216888861865, 32'sd0.035682247163253245, 32'sd0.10386759419428204, 32'sd0.13593806106309086, 32'sd0.16590629819983338, 32'sd0.0013412233964866513, 32'sd0.011170694478607779, 32'sd0.028125528807476086, 32'sd0.05979658369137054, 32'sd0.017850655674564734, 32'sd0.06304282187059798, 32'sd-0.0023706396388121454, 32'sd0.006716797749096336, 32'sd0.04788408424783853, 32'sd-0.0931920579878883, 32'sd-0.007099079852461797, 32'sd-0.16060293474843407, 32'sd0.011483010806777248, 32'sd-0.09276054929180542, 32'sd0.013701205084886408, 32'sd0.051673448765788034, 32'sd0.05814711464104793, 32'sd-0.0064303056366881925, 32'sd-0.1171199581968582, 32'sd-0.12725707119135132, 32'sd-0.126245789527698, 32'sd-0.20016276378333042, 32'sd-0.08736227420826355, 32'sd-0.18022829534214635, 32'sd-0.07256753953702631, 32'sd0.06340269357894819, 32'sd-0.003331161271630875, 32'sd-0.10093428068881526, 32'sd0.011884472781551332, 32'sd0.020420945862055177, 32'sd0.02973863749814953, 32'sd-0.01294438413917019, 32'sd-0.039515583598707084, 32'sd0.038711678130148135, 32'sd-0.05132963133551852, 32'sd-0.04211088432455317, 32'sd-0.09538432592643876, 32'sd-0.009357903980722204, 32'sd-0.04490267959030152, 32'sd-0.03851147458875017, 32'sd-0.07917977051913976, 32'sd0.03576953581252851, 32'sd-0.011853634468260234, 32'sd0.033816372454953086, 32'sd-0.014343643927495769, 32'sd-0.012316285444698897, 32'sd-0.1339188706193735, 32'sd-0.018213238315773924, 32'sd-0.10216469767641148, 32'sd-0.10436253763910334, 32'sd-0.14336714208781573, 32'sd-0.13082061699979833, 32'sd-0.07060811210217571, 32'sd0.02081760506243792, 32'sd-0.15392462216188918, 32'sd-0.05457530494880173, 32'sd-0.02811854911046472, 32'sd0.03779132890264762, 32'sd0.08778898708862902, 32'sd3.3528122556122387e-129, 32'sd0.011892043028122582, 32'sd-0.081810556577206, 32'sd-0.09396471415760069, 32'sd-0.061004670277123814, 32'sd0.03173503766779741, 32'sd0.0729209624940656, 32'sd-0.0396477442260864, 32'sd-0.05412014786806013, 32'sd-0.027379537566159136, 32'sd-0.04266778578367127, 32'sd0.011762941408155715, 32'sd0.04933315259299627, 32'sd-0.05202634531140956, 32'sd-0.0740649642886104, 32'sd0.024678760943207884, 32'sd-0.03544604624403528, 32'sd-0.06183123690193871, 32'sd-0.053746871263831285, 32'sd-0.10840355792887643, 32'sd-0.132872920191484, 32'sd-0.05470419432154152, 32'sd-0.04363291351331266, 32'sd0.01766329421197553, 32'sd0.019261582229684333, 32'sd-0.01791755000539231, 32'sd-0.04788929528207302, 32'sd6.525156391018233e-115, 32'sd-7.550170981223993e-123, 32'sd-4.873551949050259e-123, 32'sd-0.05680723253350123, 32'sd-0.09347496253561997, 32'sd0.11263739064473755, 32'sd0.06405019946035159, 32'sd-0.05072853596573981, 32'sd-0.01413397391098314, 32'sd-0.02785533743184885, 32'sd-0.029386729624572765, 32'sd0.08053559578543502, 32'sd0.02574589663859384, 32'sd0.03555249044379616, 32'sd-0.03287979296506686, 32'sd-0.03429709270669938, 32'sd-0.07174606479307055, 32'sd-0.002238211539389952, 32'sd0.02813778685237877, 32'sd-0.11558933243837728, 32'sd0.05227675221117472, 32'sd-0.038550368695768805, 32'sd0.05132449732025656, 32'sd-0.0325515113703493, 32'sd-0.044368695094963356, 32'sd-0.05789131876276469, 32'sd-0.045571874864751526, 32'sd0.056101359242868874, 32'sd2.1400698752327e-116, 32'sd-3.842299914274088e-125, 32'sd2.9432307199543074e-116, 32'sd0.014102486529195738, 32'sd0.004386544018348789, 32'sd0.047401110788579316, 32'sd0.09689632081581431, 32'sd-0.10590302552842007, 32'sd0.010158721620007933, 32'sd0.06878459523134467, 32'sd-0.06615561046311491, 32'sd0.013229936709919888, 32'sd0.13582589918743623, 32'sd0.03246462103562655, 32'sd-0.04629845471096244, 32'sd0.033169135518680816, 32'sd-0.07680142220846364, 32'sd-0.04198434755777319, 32'sd0.040329544642031485, 32'sd-0.04922757121175254, 32'sd0.03219321708782974, 32'sd-0.016046250539053623, 32'sd0.04744689586359145, 32'sd-0.03287958013921076, 32'sd-0.02740727278710286, 32'sd-0.009905023514628181, 32'sd-0.00112864051186789, 32'sd0.059394404366786495, 32'sd4.975699824272694e-115, 32'sd-1.9667316506222258e-117, 32'sd1.016987722821266e-126, 32'sd1.656030228728429e-116, 32'sd0.06884865431815429, 32'sd-0.13357105471892525, 32'sd0.03623618097167866, 32'sd-0.03645516559844538, 32'sd0.06314368036230529, 32'sd-0.0029920523294361986, 32'sd0.014454744376247426, 32'sd0.03008695563236263, 32'sd0.04725400613377517, 32'sd0.11132579646373145, 32'sd0.15055167358219715, 32'sd0.14106573845385034, 32'sd0.00037112117106005964, 32'sd0.05948979173569741, 32'sd-0.06137551877005534, 32'sd0.021114922308941277, 32'sd0.03727925676464582, 32'sd0.001965535355484108, 32'sd0.060512062926035254, 32'sd0.05728399440558008, 32'sd0.08634236590607415, 32'sd0.02343108874092118, 32'sd0.036685150322087114, 32'sd3.3411939697840625e-120, 32'sd-6.7902777307924885e-115, 32'sd-1.3504998623122147e-118, 32'sd6.558534810426332e-116, 32'sd-8.749251377271655e-127, 32'sd-1.7120862208530838e-118, 32'sd0.01625858922869315, 32'sd0.03886873809845558, 32'sd0.04944347720774978, 32'sd-0.02053092950009815, 32'sd0.02344367358631338, 32'sd-0.04118221569198734, 32'sd0.07133528293690418, 32'sd0.07742181737321052, 32'sd0.012171627296308943, 32'sd0.06777513235444567, 32'sd0.11890389774298914, 32'sd0.03584371883798606, 32'sd0.08438685384262559, 32'sd0.015648876955552993, 32'sd-0.031165879858230997, 32'sd-0.06784178618063952, 32'sd0.010610885645600124, 32'sd0.007836208034578412, 32'sd0.08602420036975707, 32'sd-0.003235559245141027, 32'sd-1.341754647651212e-122, 32'sd-8.709610531722081e-127, 32'sd-1.2037423103992335e-125, 32'sd1.0071039402106017e-115},
        '{32'sd2.831326109852331e-120, 32'sd1.3711240419368467e-126, 32'sd1.0677903430049302e-124, 32'sd1.011679900624634e-124, 32'sd3.3193666654511107e-125, 32'sd-1.7907954465701804e-122, 32'sd-2.0183278745719105e-125, 32'sd-1.7978030320122663e-127, 32'sd-6.989089940111824e-127, 32'sd2.127753259028347e-121, 32'sd6.954025714463573e-124, 32'sd2.227640283293756e-114, 32'sd-0.06011838155600882, 32'sd-0.02860763429676564, 32'sd0.016825568434004172, 32'sd-0.03907475100383915, 32'sd1.5274236142392982e-115, 32'sd-2.3329068867026425e-124, 32'sd1.2813991276309713e-118, 32'sd2.130659220282437e-126, 32'sd2.5505274095350398e-123, 32'sd5.907390403532725e-122, 32'sd-1.322096402364468e-117, 32'sd-5.2623242961569675e-124, 32'sd9.874431397005552e-120, 32'sd-6.329157590579293e-120, 32'sd6.750234157731336e-126, 32'sd3.424279052827572e-116, 32'sd3.975076644659039e-126, 32'sd3.0336299154031413e-116, 32'sd3.153655376364386e-124, 32'sd-3.3343165764742414e-120, 32'sd-0.026782862078243222, 32'sd-0.03665255507799492, 32'sd-0.06109505589173375, 32'sd-0.06528543361120963, 32'sd-0.013636120626769485, 32'sd0.11086925797303432, 32'sd0.05989801595359259, 32'sd-0.08676489296492022, 32'sd-0.1401661449737565, 32'sd-0.006145110397649029, 32'sd0.020520714093981495, 32'sd0.010200145205578834, 32'sd-0.1221047394251272, 32'sd-0.007676809054412019, 32'sd-0.007438104842537911, 32'sd0.008627145254828515, 32'sd-0.09506150389930228, 32'sd0.037927757482621595, 32'sd-0.04220276187709903, 32'sd-0.00011636360385712087, 32'sd-2.112655887628752e-117, 32'sd3.3654267052973623e-116, 32'sd-1.1458891511901066e-115, 32'sd-1.3746875722986686e-127, 32'sd5.347006162166963e-118, 32'sd-2.022379307927554e-117, 32'sd-0.0148434943737197, 32'sd0.006308646905111025, 32'sd-0.0707146584835595, 32'sd0.07876762412096217, 32'sd0.07729052778018362, 32'sd-0.037900456740271794, 32'sd-0.04602440096811942, 32'sd0.004484823449982106, 32'sd-0.008241679863359932, 32'sd0.035031922688913926, 32'sd0.049962025451741825, 32'sd-0.02223165950264322, 32'sd0.11646739335904127, 32'sd0.07012169606888141, 32'sd-0.004510367516713963, 32'sd0.007929274068028782, 32'sd-0.027121145625716957, 32'sd0.02323498472930782, 32'sd-0.02436508969831003, 32'sd-0.05338193814670457, 32'sd-0.07340109606290526, 32'sd-0.0029104013953629537, 32'sd-0.025733953962676387, 32'sd-0.034479339154491376, 32'sd6.680449927487603e-127, 32'sd-3.5050169579879267e-115, 32'sd-2.384057621035742e-125, 32'sd4.762717467799967e-122, 32'sd-0.0139947996246132, 32'sd0.06336449816037013, 32'sd0.028453457489501444, 32'sd-0.081628088532523, 32'sd-0.06706209308134528, 32'sd-0.0245432118637983, 32'sd-0.04710889238408195, 32'sd0.01774929715645498, 32'sd-0.03925843221416887, 32'sd-0.04487806911302715, 32'sd-0.013187590300841517, 32'sd-0.026195272560560222, 32'sd-0.09399549837086464, 32'sd0.033310130016695125, 32'sd0.022413400454536866, 32'sd-0.06765307807465236, 32'sd-0.06887682629697238, 32'sd0.0361470611362069, 32'sd0.05171491081069039, 32'sd0.02355381339908956, 32'sd-0.053741600379979375, 32'sd-0.033068206698222344, 32'sd-0.03663407107694673, 32'sd-0.04121088459800545, 32'sd-0.09394787220455621, 32'sd-2.0140396098833406e-121, 32'sd-1.468659154351676e-124, 32'sd0.01591238286478093, 32'sd0.041670230948256386, 32'sd-0.012952188683844944, 32'sd0.0028952438073390936, 32'sd-0.02594971303461877, 32'sd0.0107723456388564, 32'sd0.034018516009488756, 32'sd-0.01337881966712236, 32'sd-0.11093777597763939, 32'sd-0.09597008565460895, 32'sd-0.05730259885954997, 32'sd-0.0943419961011359, 32'sd-0.01849625217193773, 32'sd-0.11129385005090316, 32'sd-0.09427780317182546, 32'sd-0.12326316305697889, 32'sd-0.08519931604055583, 32'sd-0.01796068394719272, 32'sd-0.12310152695749776, 32'sd-0.015085353327408194, 32'sd0.0010397094046165022, 32'sd-0.033387790780386714, 32'sd-0.1444662428178415, 32'sd0.07271789775660227, 32'sd0.06561355910202032, 32'sd0.08762678319500523, 32'sd-0.018170592840744553, 32'sd-1.1213263445172075e-121, 32'sd-0.03968198120492697, 32'sd-0.04450468563683231, 32'sd-0.03524363858598093, 32'sd0.056255113946874186, 32'sd-0.07830446869426243, 32'sd-0.07044210447947383, 32'sd-0.09206888806976457, 32'sd-0.08931243061230157, 32'sd-0.1328038640798875, 32'sd0.061359339473700904, 32'sd-0.03179448740796569, 32'sd-0.009289479398343745, 32'sd-0.01906993744849366, 32'sd-0.04828107672686062, 32'sd-0.17146967880272437, 32'sd0.005615015996452482, 32'sd-0.12973633147956357, 32'sd-0.08767787097325376, 32'sd0.08186533355992887, 32'sd0.04793870898037563, 32'sd0.03246624435438114, 32'sd-0.09308487044932588, 32'sd-0.09277044774386992, 32'sd0.08984645284649787, 32'sd0.10918152740670028, 32'sd0.048621745163963996, 32'sd-0.052281974602845005, 32'sd-4.169644682351935e-125, 32'sd-0.02264560969192562, 32'sd0.015001954764366844, 32'sd-0.01880070090474437, 32'sd0.02607884084758641, 32'sd-0.10060661395525997, 32'sd-0.09570408070906558, 32'sd-0.09742947087180946, 32'sd0.007594335507934573, 32'sd-0.06586511717269354, 32'sd-0.014239873140278154, 32'sd0.09652387250754, 32'sd0.104012885582208, 32'sd0.042577010078941394, 32'sd-0.10010946531440827, 32'sd-0.03620773163955177, 32'sd0.12275173161507885, 32'sd0.09276088464315978, 32'sd0.02331855332446362, 32'sd0.10314018978577703, 32'sd-0.014408444144409192, 32'sd-0.06514118041941051, 32'sd-0.14932059765314287, 32'sd-0.08267325010055787, 32'sd-0.06893626154787008, 32'sd0.0427611475475635, 32'sd0.09010785531386167, 32'sd-0.004768805177304256, 32'sd-0.04176370668395741, 32'sd-0.010430147824769172, 32'sd-0.06067654295594309, 32'sd0.01565135583360006, 32'sd-0.015430064432053168, 32'sd-0.07806945486612475, 32'sd-0.12490057601785712, 32'sd-0.056976398198823344, 32'sd-0.12356259997508659, 32'sd-0.07317567853388675, 32'sd0.04329857038812833, 32'sd-0.05846714882755258, 32'sd0.04206885996275568, 32'sd0.03665253958216355, 32'sd0.0226959079927534, 32'sd0.01616800372907554, 32'sd-0.11059317052598319, 32'sd-0.07589695179966437, 32'sd0.0535599649365388, 32'sd0.17050247074405137, 32'sd0.021395293445896045, 32'sd-0.00670037673147747, 32'sd0.04391022370491471, 32'sd-0.16368181862564427, 32'sd-0.03766406729173093, 32'sd-0.060295425402534554, 32'sd-0.10520230236628778, 32'sd0.055291216387245636, 32'sd-0.028134285952516297, 32'sd0.02129292450796789, 32'sd-0.032983780744414756, 32'sd-0.004505203022882849, 32'sd0.04284549324118722, 32'sd-0.007006288035215076, 32'sd0.00547059361186145, 32'sd-0.07828878026074271, 32'sd-0.06191861366742352, 32'sd-0.14469404409196976, 32'sd-0.12678269632741365, 32'sd0.0022027490868087173, 32'sd-0.08747284064661594, 32'sd-0.07710704307524988, 32'sd0.0206453378238527, 32'sd-0.01355334178523251, 32'sd-0.11597547831373982, 32'sd-0.07006397026596703, 32'sd0.07494624586342839, 32'sd-0.054517570252870184, 32'sd-0.013669998223522679, 32'sd0.0865084942885448, 32'sd-0.062296937432137295, 32'sd-0.06514426238463285, 32'sd0.04488368398986366, 32'sd-0.10187928373728398, 32'sd-0.009827593933587444, 32'sd-0.06210823927208639, 32'sd0.042759203625032, 32'sd0.12441996156030442, 32'sd-0.10449796247970117, 32'sd0.03902944839491579, 32'sd0.05383705488913428, 32'sd-0.09312067869421722, 32'sd0.08589864546509544, 32'sd-0.0208536304682839, 32'sd-0.07295514332353602, 32'sd0.07113840893914707, 32'sd-0.0895087306771198, 32'sd0.0036344130442845035, 32'sd-0.11626033647782576, 32'sd0.07805235831056721, 32'sd0.07653133674666428, 32'sd0.03160449605547156, 32'sd-0.009157561165539889, 32'sd0.001768026703711024, 32'sd-0.046934295670766284, 32'sd-0.03829668607251203, 32'sd-0.08070774300509731, 32'sd0.14513506277799343, 32'sd-0.03112852689569623, 32'sd-0.11082069892692133, 32'sd-0.08922125758795547, 32'sd-0.10849048944407579, 32'sd-0.08985919402269646, 32'sd-0.07554965885435587, 32'sd0.07692660732507091, 32'sd-0.0617841756436608, 32'sd-0.11233668462409648, 32'sd0.005944801721006444, 32'sd-0.04288078506795271, 32'sd-0.03028902047461682, 32'sd0.006261008050036099, 32'sd-0.11042220452204309, 32'sd-0.01347264992759506, 32'sd-0.02100887907568232, 32'sd0.07898454383011416, 32'sd-0.0775423285333547, 32'sd-0.08383492700224852, 32'sd-0.014431952628758554, 32'sd0.10375557962631653, 32'sd-0.02332604195531156, 32'sd-0.023148597536265133, 32'sd-0.18966702054572526, 32'sd-0.011005193372679137, 32'sd0.012496328076542522, 32'sd-0.07127258368529601, 32'sd0.07229526787064652, 32'sd-0.07551150918403893, 32'sd-0.06566748031380676, 32'sd-0.014804439421082172, 32'sd-0.1415595637624114, 32'sd-0.010313728522779005, 32'sd-0.10027044410621168, 32'sd0.042096289651203704, 32'sd-0.20453510281636603, 32'sd-0.020777717818890987, 32'sd-0.03048838968001106, 32'sd-0.0008423046280886947, 32'sd0.07548959545949543, 32'sd0.055009974723538135, 32'sd0.06372541301543759, 32'sd0.09874673509913581, 32'sd0.020504419412013555, 32'sd-0.062274544687686804, 32'sd-0.19354498102662834, 32'sd-0.23781402759426956, 32'sd-0.16203304818857306, 32'sd-0.01516501853406353, 32'sd-0.019740835983139898, 32'sd-0.23142839224892414, 32'sd-0.13482783645103494, 32'sd0.040395962111016204, 32'sd-0.060237791296269265, 32'sd-0.005382997936556726, 32'sd0.014688162363217606, 32'sd0.03231587574139932, 32'sd0.03357412536332556, 32'sd-0.01674165215047189, 32'sd0.027394504399973575, 32'sd0.0752908711928228, 32'sd0.06375267163941616, 32'sd-0.06864636392342571, 32'sd-0.05466422785660402, 32'sd0.01365991170420438, 32'sd-0.004543332650041172, 32'sd0.0014702381302400353, 32'sd0.04483834239816632, 32'sd0.03582379577092617, 32'sd-0.0054069475925819736, 32'sd0.13931880983902756, 32'sd0.0899086375989252, 32'sd-0.014061308693408674, 32'sd-0.1314374995185553, 32'sd-0.2991460825994182, 32'sd-0.21813869407001973, 32'sd-0.07444119185696574, 32'sd-0.16711547066001428, 32'sd-0.149278620072181, 32'sd0.0585948789663326, 32'sd0.04632611932443404, 32'sd-0.02839102016650601, 32'sd0.08039646073890867, 32'sd0.1645953084448783, 32'sd-0.021801702101155295, 32'sd0.015327410548493734, 32'sd0.08275700749620107, 32'sd-0.05370901323026272, 32'sd-0.07196952768923491, 32'sd-0.011426064197513689, 32'sd-0.007030904733412499, 32'sd-0.013711689482318289, 32'sd-0.016590233666513705, 32'sd-0.09630356750267591, 32'sd-0.06386180385026179, 32'sd0.10968883947723321, 32'sd0.06594368109157676, 32'sd0.06464781136146534, 32'sd0.11708845490705988, 32'sd0.03694708392965777, 32'sd0.082031266580367, 32'sd-0.007338789209230385, 32'sd-0.11507070452484763, 32'sd-0.10471059436626623, 32'sd-0.0459428662609714, 32'sd0.13742931032348804, 32'sd0.07583225819121225, 32'sd0.08617711565282564, 32'sd0.08349844661268975, 32'sd0.08193702833259187, 32'sd0.041089950819259875, 32'sd0.15163257744403433, 32'sd0.09993987358605398, 32'sd0.03427013781491292, 32'sd-0.05712267665041825, 32'sd0.1176543000446209, 32'sd-0.00182790867595755, 32'sd-0.03024137769386496, 32'sd-0.028763528001370685, 32'sd-0.05909293204418531, 32'sd-0.047361359338858794, 32'sd-0.043636512728118616, 32'sd0.014976921958047494, 32'sd-0.040271823222333365, 32'sd0.13883818234324166, 32'sd0.004730888122507805, 32'sd0.007437230002727312, 32'sd0.08675706759704284, 32'sd0.26678169458402784, 32'sd0.187034348486129, 32'sd0.06048966215064734, 32'sd0.05673714193559468, 32'sd0.09281001334827757, 32'sd-0.010508340670215683, 32'sd0.07845348455507348, 32'sd0.11681516014294425, 32'sd0.04816031462786591, 32'sd0.038354815863910874, 32'sd-0.04238287428995214, 32'sd-0.02323747669758626, 32'sd-0.05917353049851251, 32'sd0.019770133362998422, 32'sd-0.02512126485966977, 32'sd0.06715918400274842, 32'sd0.031894196153294536, 32'sd-0.06361471122137331, 32'sd0.011211029201201664, 32'sd-0.03280702937741453, 32'sd-0.006105473841308589, 32'sd-0.02659956138756355, 32'sd0.01570345507043161, 32'sd0.0442994772846639, 32'sd0.12310007800546169, 32'sd0.03547976800530588, 32'sd0.09815941594728798, 32'sd0.2087183414427964, 32'sd0.23148213980927784, 32'sd0.16007851447232996, 32'sd0.23084902528904164, 32'sd0.06587066910178009, 32'sd0.08467904422879909, 32'sd0.034971331660896936, 32'sd0.024523696356863564, 32'sd0.11594570511142717, 32'sd0.15122984044244245, 32'sd0.03981158064932756, 32'sd-0.044380379748833625, 32'sd-0.05426733655999059, 32'sd0.02603054345572544, 32'sd0.051996333551214954, 32'sd0.025070872688640722, 32'sd0.12187111768416303, 32'sd0.10655051716536891, 32'sd0.04288886539183498, 32'sd-0.03666767092330205, 32'sd0.028995277509749926, 32'sd-0.1070208413476205, 32'sd-0.030152833563065255, 32'sd0.003684307962766699, 32'sd0.019097798895481976, 32'sd0.112533925869994, 32'sd0.0963409193921514, 32'sd0.057631573358992334, 32'sd0.06860947204850593, 32'sd0.015386946816102297, 32'sd0.09992709381064878, 32'sd0.16527631895504052, 32'sd0.20698767481039385, 32'sd-0.007741380272135087, 32'sd-0.09162543448117567, 32'sd0.11287423271538444, 32'sd0.08271865038262938, 32'sd0.026640949147342278, 32'sd-0.04033096524688412, 32'sd0.06876379090963212, 32'sd-0.03271013581667314, 32'sd0.02968340967810192, 32'sd0.0012820243223061168, 32'sd0.002323258916830575, 32'sd-0.04523837076551691, 32'sd-0.018178224852925556, 32'sd0.02096470264745403, 32'sd4.7510720309175724e-123, 32'sd-0.029710128214009816, 32'sd0.020324421640120303, 32'sd-0.0008672557236534331, 32'sd0.04199709819115484, 32'sd0.011410034758913399, 32'sd-0.020280447926025697, 32'sd-0.010116448333782455, 32'sd-0.01194313136673797, 32'sd-0.10359660613369982, 32'sd-0.06021181604373815, 32'sd-0.03623222566985453, 32'sd0.12703442222852884, 32'sd0.04500057701893225, 32'sd0.010763459633386985, 32'sd0.10470835967098867, 32'sd0.02369214625858602, 32'sd0.036272243245141306, 32'sd-0.07458873784932209, 32'sd-0.05603891900118145, 32'sd0.06278366972637757, 32'sd-0.012110768438303124, 32'sd-0.08444597723468195, 32'sd-0.08096671933974497, 32'sd0.03494911767819859, 32'sd0.027881320503977607, 32'sd0.005089542329531991, 32'sd0.0067302815214291085, 32'sd-0.031609013770127994, 32'sd0.046669746655382885, 32'sd-0.06350237540301217, 32'sd-0.03587552839788981, 32'sd0.03606556573910413, 32'sd0.055943981877007956, 32'sd0.16904842345375104, 32'sd0.10519167299991625, 32'sd-0.07898744508882, 32'sd-0.14043896377545662, 32'sd0.04584622263828837, 32'sd-0.035893620811393, 32'sd-0.017959593304926337, 32'sd0.14050470366751955, 32'sd0.13373281280198748, 32'sd-0.010195369342936947, 32'sd0.02603633079164971, 32'sd-0.06521778667092487, 32'sd0.047476763063441084, 32'sd-0.08939229215616444, 32'sd-0.004079509035363864, 32'sd-0.04074624091404451, 32'sd0.009438485195680036, 32'sd-0.0678152667177098, 32'sd-0.04775848315826465, 32'sd-0.10422880778708782, 32'sd-0.0031141769056486786, 32'sd-0.03931140495487746, 32'sd-0.05867981413757575, 32'sd0.0019823753844790165, 32'sd0.05161964878986942, 32'sd0.030859447296744065, 32'sd-0.0029574228126739164, 32'sd0.07076834329370223, 32'sd0.005997094947312723, 32'sd0.04871933969806645, 32'sd-0.06874492914486413, 32'sd-0.0011329069127894206, 32'sd-0.0160238711708093, 32'sd0.056057924158461225, 32'sd0.11835220959833617, 32'sd0.1695903891169003, 32'sd0.14991517816693672, 32'sd-0.044899845531926504, 32'sd-0.02227076065308773, 32'sd-0.06407442984340504, 32'sd-0.013513135990211887, 32'sd0.06522116367675214, 32'sd-0.10506723574638614, 32'sd0.08618795873847865, 32'sd-0.021585855603966267, 32'sd0.03189680763741573, 32'sd-0.1252982263127457, 32'sd0.010492052169202674, 32'sd0.03186380540858283, 32'sd-0.05141510684120433, 32'sd-1.0804901596082637e-121, 32'sd0.015192028097083301, 32'sd0.09555077093819327, 32'sd-0.11333007367200733, 32'sd-0.09768744880300352, 32'sd-0.00635715235510984, 32'sd-0.020856872170841718, 32'sd0.04129160626480839, 32'sd-0.033989066652087965, 32'sd-0.011709871001947736, 32'sd0.031185628406542237, 32'sd0.055422174913201804, 32'sd0.033563038088215036, 32'sd0.09293650111973502, 32'sd-0.049878030647168274, 32'sd-0.06317464788737429, 32'sd-0.0028214474797356626, 32'sd0.02058692226454173, 32'sd0.13135514326763117, 32'sd0.004055563416051332, 32'sd-0.032531853776415647, 32'sd-0.029989800931389973, 32'sd-0.027581082257051994, 32'sd0.030351858428321516, 32'sd0.010804555464930457, 32'sd-0.004017616602494371, 32'sd-0.039970273748044106, 32'sd-0.05563211906936136, 32'sd0.0022085456363718117, 32'sd0.02842188347637212, 32'sd0.12966427629011845, 32'sd-0.023711521325761497, 32'sd0.04094835953308192, 32'sd0.1704387077053587, 32'sd0.07285752435643411, 32'sd-0.08540558514439914, 32'sd0.0651057071439168, 32'sd-0.005340041340821822, 32'sd0.0522890624370435, 32'sd0.0326458975687581, 32'sd-0.054225385370191795, 32'sd-0.0005175201414754272, 32'sd0.0892651353496157, 32'sd-0.0015785828953821393, 32'sd-0.12651821650082606, 32'sd0.0031447295274462292, 32'sd-0.08133847715891662, 32'sd0.010574393643398778, 32'sd0.014874567011053805, 32'sd0.0012899903796552053, 32'sd-0.07278142061606527, 32'sd0.07825923451185768, 32'sd0.12048007535263065, 32'sd-0.12762958953005263, 32'sd-0.01760320311671876, 32'sd-0.009214095825811734, 32'sd-0.024460642818016295, 32'sd0.06040784247818368, 32'sd0.08113442559805524, 32'sd-0.05765387470673182, 32'sd0.09875531242031683, 32'sd-0.05337786057289149, 32'sd-0.056483192074414636, 32'sd0.010630981884547485, 32'sd-0.0036199392643196317, 32'sd-0.07238692667698343, 32'sd-0.10423568823811559, 32'sd-0.06914521152654521, 32'sd-0.02830610736286042, 32'sd-0.08488544312421957, 32'sd-0.13415393226200553, 32'sd-0.15384905661851817, 32'sd-0.02307685720951039, 32'sd-0.005393560950015647, 32'sd-0.06353223226230699, 32'sd-0.06279691471387369, 32'sd-0.03694341769236264, 32'sd-0.07189060400830022, 32'sd0.06920059133574162, 32'sd0.13505243418748702, 32'sd0.025491172104214515, 32'sd-0.019378073844016717, 32'sd-0.02438587395106745, 32'sd-0.027783177093522612, 32'sd-2.2059834885798783e-119, 32'sd-0.016630027173384087, 32'sd0.02039892014863727, 32'sd0.03414422990167774, 32'sd0.1231901657436675, 32'sd0.14698856603077576, 32'sd-0.03639537515560738, 32'sd0.01123812971358478, 32'sd-0.022602186413233426, 32'sd-0.06973917038876445, 32'sd0.019104433306203414, 32'sd-0.006997219416953105, 32'sd-0.11004120639710031, 32'sd-0.07449297841469651, 32'sd0.009670892922380091, 32'sd0.03704828084052026, 32'sd0.0705482765744245, 32'sd0.04603503834464101, 32'sd0.038331773832315515, 32'sd-0.06515532625431891, 32'sd0.1020988876791949, 32'sd0.027203147960631013, 32'sd0.0811777236500917, 32'sd0.06393791635862418, 32'sd-0.0023871711568467565, 32'sd-0.011228522536721474, 32'sd-0.04134367749244177, 32'sd-2.645678234630317e-120, 32'sd-6.798782601468386e-124, 32'sd2.293664513371458e-114, 32'sd-0.019859260068400404, 32'sd-0.017297653967440284, 32'sd0.08317829725900543, 32'sd-0.060432532728772775, 32'sd0.012134088671386942, 32'sd0.03330931316688097, 32'sd0.017482318861975578, 32'sd0.06194191543508187, 32'sd-0.05856436144190492, 32'sd-0.08864357542148034, 32'sd0.03502613598925972, 32'sd0.006263819030310345, 32'sd0.0005606529611494257, 32'sd0.06472416573874575, 32'sd-0.07439728203188845, 32'sd0.009793369516586825, 32'sd0.08327303392516808, 32'sd0.008048656546397264, 32'sd0.002878365157022946, 32'sd-0.023079727276766545, 32'sd0.10853321979920057, 32'sd-0.004043904873496794, 32'sd-0.00751407154430539, 32'sd-0.034598033550291285, 32'sd0.0862504859474501, 32'sd9.239054748904752e-122, 32'sd-6.884081737598312e-126, 32'sd-4.956737144006132e-126, 32'sd-0.049842633372429966, 32'sd0.020123754121002282, 32'sd-0.03088743021556828, 32'sd-0.09823493152090265, 32'sd0.054762258587895275, 32'sd-0.06920441737009143, 32'sd-0.03668950639260633, 32'sd0.0009619844262922599, 32'sd0.11616984499694447, 32'sd0.03798384956384854, 32'sd-0.09755248632041998, 32'sd-0.17181494017269192, 32'sd-0.023077868803396115, 32'sd-0.11595902117429596, 32'sd0.02728336148191272, 32'sd-0.06263771307241583, 32'sd0.010845479006898471, 32'sd0.010736733756496097, 32'sd0.0021322123604081552, 32'sd0.024366588970277228, 32'sd0.017629307317198084, 32'sd0.016898792047797408, 32'sd-0.020011159773735163, 32'sd0.013897775273102942, 32'sd0.08173859417512407, 32'sd3.577108537009587e-117, 32'sd7.820816970493253e-128, 32'sd-1.0269522564446904e-124, 32'sd6.618338464752915e-126, 32'sd-0.021714561740658455, 32'sd0.08797124526273904, 32'sd-0.07856675364340157, 32'sd0.016896189418998706, 32'sd-0.03948862810426668, 32'sd-0.019390078093567763, 32'sd0.02429432082924728, 32'sd-0.009170955874264024, 32'sd-0.12834512251054012, 32'sd-0.0706785897738432, 32'sd0.09724854121248931, 32'sd-0.021138292333097667, 32'sd-0.08673961871455955, 32'sd0.1496269949042983, 32'sd0.06197742323046368, 32'sd0.09161999475262096, 32'sd-0.00014276626622702, 32'sd-0.009362130730408213, 32'sd-0.07292085423319812, 32'sd0.00791022150223176, 32'sd0.046788963504561396, 32'sd-0.0129142668288079, 32'sd-0.05156238282496547, 32'sd8.182417152885286e-118, 32'sd1.529895703617429e-122, 32'sd6.89995862769717e-117, 32'sd-2.2811323880853553e-126, 32'sd2.4755900853419624e-126, 32'sd-3.1788062100925566e-129, 32'sd-0.06419862870994421, 32'sd-0.03199801964645676, 32'sd0.0683094193058643, 32'sd0.06030303648920428, 32'sd-0.01954338932269372, 32'sd-0.018551515876822147, 32'sd0.06274725981520912, 32'sd0.04982517011526963, 32'sd-0.01332525728857694, 32'sd-0.02101963920122549, 32'sd0.05777065921592257, 32'sd-0.00413079434510608, 32'sd-0.08692596412634994, 32'sd-0.039673570948438514, 32'sd0.02472838935551678, 32'sd0.03735836194889438, 32'sd-0.007231207776884375, 32'sd-0.015244736435487283, 32'sd-0.058695459221531444, 32'sd-0.046553593579326674, 32'sd4.787052125072658e-123, 32'sd1.5921486148574736e-114, 32'sd1.1119660161885922e-121, 32'sd6.887841466647209e-126},
        '{32'sd-5.2240101340404925e-118, 32'sd-2.7972202030925777e-119, 32'sd5.179881072208727e-127, 32'sd1.1845849165070432e-122, 32'sd-9.957102833261332e-116, 32'sd-1.8460779053868836e-117, 32'sd6.182054781298706e-115, 32'sd-1.8217077795767383e-115, 32'sd5.056510721461289e-118, 32'sd1.0093766262329878e-119, 32'sd1.0493942088522472e-120, 32'sd4.795975779030994e-123, 32'sd0.023195123562699566, 32'sd0.039518355270268125, 32'sd0.06843876147396755, 32'sd-0.007804869736097597, 32'sd-1.0900598247836635e-118, 32'sd1.6728849775463886e-127, 32'sd2.3523044926452077e-122, 32'sd-6.889375688378733e-124, 32'sd-8.326372348303577e-116, 32'sd3.2687963288939945e-120, 32'sd3.392953369977528e-120, 32'sd1.6982403302692692e-120, 32'sd3.7603717455087363e-123, 32'sd4.4819576381849984e-120, 32'sd3.3581738699838582e-121, 32'sd-3.557551289025599e-118, 32'sd7.447329863677491e-128, 32'sd2.0650400973089784e-120, 32'sd-8.880330167108226e-124, 32'sd-5.824690529713815e-117, 32'sd0.0731535420111072, 32'sd0.024631224586921286, 32'sd0.015880378384440366, 32'sd0.07508834721187715, 32'sd0.08677842246662727, 32'sd0.05540842274180621, 32'sd-0.07033957420324068, 32'sd0.006866379563108124, 32'sd0.02167500640577515, 32'sd0.0532446245936796, 32'sd-0.06863287223212453, 32'sd0.0720995050507153, 32'sd0.05282599815201123, 32'sd0.11161058980047585, 32'sd0.06582277858313239, 32'sd-0.01120360446601199, 32'sd-0.01832030501750538, 32'sd0.015640661620020136, 32'sd-0.004831270588398877, 32'sd0.022230093225112994, 32'sd-5.572978410292689e-119, 32'sd1.5259800355453702e-115, 32'sd6.428938973378362e-115, 32'sd-2.662495341474881e-114, 32'sd6.669742292446834e-127, 32'sd1.1068106868315582e-121, 32'sd-0.008572723157739957, 32'sd0.005352626665002929, 32'sd0.047004594945662635, 32'sd0.020418432435478806, 32'sd0.024646649415985888, 32'sd0.014703623138230884, 32'sd-0.10456334660307892, 32'sd0.08310621699503078, 32'sd-0.009821101389237953, 32'sd-0.016030591321385426, 32'sd-0.007927924372703916, 32'sd-0.024517648582636047, 32'sd0.03159517315917843, 32'sd0.14888542582431538, 32'sd0.04998350880308438, 32'sd0.06770708955255599, 32'sd-0.05487748389376685, 32'sd0.07690608080114537, 32'sd-0.02568695972548786, 32'sd0.061726127973058084, 32'sd-0.055674249175128906, 32'sd-0.04080703500424548, 32'sd0.01961064549963381, 32'sd0.0637045644450173, 32'sd-8.812046666161472e-127, 32'sd1.3205011419183228e-122, 32'sd-1.2464603721662268e-126, 32'sd-1.2687049736927757e-114, 32'sd0.024105103543772294, 32'sd-0.03647039608383825, 32'sd-0.003843190782500849, 32'sd-0.0744976649360094, 32'sd0.006482186372887864, 32'sd0.020739979144404858, 32'sd-0.08925093702515523, 32'sd-0.014471567511651592, 32'sd-0.042668109223238576, 32'sd-0.0858428351550096, 32'sd-0.01397312892099279, 32'sd-0.033317067424205, 32'sd-0.025436982413195884, 32'sd-0.043383338850528676, 32'sd0.028777776793892165, 32'sd-0.04674235994637453, 32'sd-0.08457371575757883, 32'sd0.056487678379713434, 32'sd-0.007514096057207576, 32'sd-0.0462373067589331, 32'sd-0.02534122898293021, 32'sd0.04500067342061391, 32'sd0.07545604646207646, 32'sd0.01797773149995729, 32'sd0.03918380148428797, 32'sd1.489474947745623e-119, 32'sd7.47972579438505e-122, 32'sd0.009848398722372781, 32'sd0.008724500418688049, 32'sd-0.11196516802361217, 32'sd-0.010419524249903854, 32'sd0.10464478120678362, 32'sd-0.06780807280646055, 32'sd-0.09658915794149366, 32'sd-0.08029067701329068, 32'sd-0.03099090695313539, 32'sd-0.001235727291627579, 32'sd0.07783605824070197, 32'sd-0.043274001295752075, 32'sd-0.06444366672552906, 32'sd-0.09380016478361597, 32'sd-0.08294819076999173, 32'sd0.11324782843598519, 32'sd-0.08449974044121863, 32'sd-0.09011268966833992, 32'sd-0.12264217919077215, 32'sd-0.07467576885757439, 32'sd-0.031666360643324475, 32'sd-0.01805228396034888, 32'sd0.012546875246425466, 32'sd-0.010424689600096015, 32'sd-0.04784901175769033, 32'sd-0.08496275335104238, 32'sd0.010858032674933094, 32'sd-7.366539828876783e-122, 32'sd-0.020851250724273896, 32'sd0.029759078430726848, 32'sd0.10604773913469602, 32'sd0.1176171576739803, 32'sd0.0023316228352939523, 32'sd0.0668300870591897, 32'sd0.12388271875259275, 32'sd0.05595787856947306, 32'sd0.02707311992133089, 32'sd0.05649764300198587, 32'sd-0.00394691907414679, 32'sd0.0014362361490651125, 32'sd0.08486447292745573, 32'sd0.06005355655256999, 32'sd0.1615866416898953, 32'sd0.16563594092112946, 32'sd-0.015953116839086297, 32'sd-0.08532004836072718, 32'sd-0.2280227230804295, 32'sd-0.03530244930459276, 32'sd-0.10373651315729672, 32'sd0.015623581619381061, 32'sd-0.02853680306954767, 32'sd-0.022206637904034616, 32'sd-0.06224495209403838, 32'sd0.00904016620386768, 32'sd-0.02132913880370944, 32'sd1.5473513139821692e-123, 32'sd0.06509701473805002, 32'sd-0.010001377075605737, 32'sd-0.023236953965582185, 32'sd-0.03941631180372112, 32'sd0.010151482629452107, 32'sd0.03475611617925662, 32'sd0.012982211741844147, 32'sd-0.018885134208166825, 32'sd0.09647043151180304, 32'sd0.07696421404003476, 32'sd0.01616382729232086, 32'sd0.09448762458353732, 32'sd0.046760434168468826, 32'sd0.10743805937342639, 32'sd0.16332382562029577, 32'sd0.17520032344867084, 32'sd0.0032312416311716776, 32'sd-0.029633643333741005, 32'sd-0.11594142549934659, 32'sd-0.09734219153755908, 32'sd0.05194821954253336, 32'sd-0.04478616338559288, 32'sd-0.035121883612317085, 32'sd-0.03673244583625538, 32'sd-0.0482312394103938, 32'sd0.032262411217689434, 32'sd-0.0630244248293343, 32'sd-0.005425069410454213, 32'sd-0.0032789321749196955, 32'sd0.025076566201446916, 32'sd0.030705225753835674, 32'sd-0.05578865700808305, 32'sd-0.01643851138327091, 32'sd-0.06407655262458367, 32'sd0.082324774513142, 32'sd-0.1543472894382984, 32'sd-0.08033059375034637, 32'sd0.04731820263831088, 32'sd0.03732898228613702, 32'sd0.07524862840247366, 32'sd0.11531231813959317, 32'sd0.03389870602693323, 32'sd-0.015570851415401907, 32'sd0.13708912458329855, 32'sd-0.0415903131299399, 32'sd-0.20053415677216505, 32'sd-0.12147047602168301, 32'sd-0.17599581806565942, 32'sd-0.12847062102378679, 32'sd-0.13396893939548712, 32'sd-0.12438256218381905, 32'sd-0.050654044871105156, 32'sd0.021674736441520553, 32'sd0.028918381082963754, 32'sd0.0016990805783476967, 32'sd0.026743245944431355, 32'sd-0.0647280343396262, 32'sd-0.05206491187146537, 32'sd-0.029209288615960765, 32'sd0.047450147532583566, 32'sd-0.010002603590198684, 32'sd-0.12227028877066365, 32'sd-0.028594584915600723, 32'sd-0.15512446883433303, 32'sd-0.12315994171735849, 32'sd-0.0033022654101136943, 32'sd0.034535523608415594, 32'sd-0.015107266471061385, 32'sd0.12686141604196752, 32'sd0.20533196935648643, 32'sd0.2639842336655796, 32'sd0.14788646938036296, 32'sd0.030204732852393806, 32'sd-0.19500510888266684, 32'sd-0.16828348401052107, 32'sd-0.16338748023466176, 32'sd-0.1359927972060631, 32'sd-0.18762750371079917, 32'sd-0.051123732663499746, 32'sd0.09131589118758295, 32'sd0.04028250812129768, 32'sd0.08043211975295608, 32'sd-0.05199084307850469, 32'sd0.03111167009921473, 32'sd0.10088313883835259, 32'sd-0.042057794416794615, 32'sd-0.08406831191358581, 32'sd0.07961691106470167, 32'sd-0.04150263510616839, 32'sd0.06468190566189304, 32'sd-0.11746324061690178, 32'sd-0.1202491911408423, 32'sd-0.09675511380803127, 32'sd-0.16268139308848173, 32'sd-0.18414898776982808, 32'sd0.09780058748183908, 32'sd0.06723101513096655, 32'sd0.082991046286289, 32'sd0.232961793706766, 32'sd0.16943389100596246, 32'sd-0.02962207012304943, 32'sd-0.1395403851610479, 32'sd-0.14367262767261604, 32'sd-0.1523050056837943, 32'sd-0.21191237263998722, 32'sd-0.10587910205067187, 32'sd-0.07943165908264305, 32'sd0.08322363694410045, 32'sd0.09039863639668017, 32'sd0.08424158142446117, 32'sd0.0011257065007846448, 32'sd0.023421335684240485, 32'sd0.019599980790891543, 32'sd-0.08655700460432747, 32'sd-0.13260468577970805, 32'sd-0.04758279648279304, 32'sd-0.029948957861058046, 32'sd0.006322164618565164, 32'sd-0.12970036177339334, 32'sd-0.08714276279370493, 32'sd-0.1499940138786691, 32'sd-0.06308370477116441, 32'sd-0.07409785731928467, 32'sd-0.030610777410994962, 32'sd0.0994320497392286, 32'sd0.1411492771853403, 32'sd0.2395513728843135, 32'sd0.0597458149832795, 32'sd-0.10196575301170234, 32'sd-0.1985244975704384, 32'sd-0.18274133318360147, 32'sd-0.11456611207826282, 32'sd-0.08474755337365175, 32'sd-0.08763090463630423, 32'sd-0.11732014011023562, 32'sd-0.04307565439249532, 32'sd0.1327987201001229, 32'sd0.10070849730800774, 32'sd0.050427243435133086, 32'sd0.00035680609958370173, 32'sd0.0066895123646102395, 32'sd-0.04929383433326951, 32'sd-0.08235585357675958, 32'sd-0.02887915697050711, 32'sd0.08932882367045338, 32'sd-0.014288778024915669, 32'sd-0.02820774377900938, 32'sd0.07518487465632939, 32'sd-0.03806284048545253, 32'sd-0.07887200230163352, 32'sd0.022596386784139316, 32'sd0.08742252863058182, 32'sd0.10000691242221381, 32'sd0.2118008685231793, 32'sd0.06890580101588713, 32'sd-0.020995543256246283, 32'sd-0.09972458613865275, 32'sd-0.16828261849668713, 32'sd-0.035533214569040655, 32'sd-0.050210467059647934, 32'sd-0.12197076791243125, 32'sd-0.030822362533810446, 32'sd-0.05371914501557687, 32'sd-0.09352319104425691, 32'sd-0.06237259805237992, 32'sd0.046434045657333535, 32'sd-0.0384837501996406, 32'sd0.020387536994847088, 32'sd-0.05091376765521896, 32'sd-0.08569350038755964, 32'sd-0.05173663093510389, 32'sd-0.049307329651729466, 32'sd0.05256281330916937, 32'sd-0.02582824851716708, 32'sd0.025535196260394143, 32'sd0.04119188950814517, 32'sd-0.09088640415477801, 32'sd0.033847590189754806, 32'sd-0.06736785600826163, 32'sd0.031041961197226, 32'sd0.167657715207526, 32'sd0.06153255665048593, 32'sd-0.0517490656726857, 32'sd-0.048950387070720344, 32'sd-0.14082010601505024, 32'sd-0.10350123253955529, 32'sd-0.13142863930464774, 32'sd-0.14695276463393014, 32'sd-0.10957672250794086, 32'sd0.05481580097461079, 32'sd-0.04816830946465977, 32'sd-0.02259906368884317, 32'sd0.027112746353237325, 32'sd-0.004852259713861064, 32'sd-0.00763649279203255, 32'sd-0.0036507180638370384, 32'sd-0.043916068909405026, 32'sd0.009884908815316434, 32'sd-0.09623585681676089, 32'sd-0.12966769006266388, 32'sd-0.018485482029582397, 32'sd0.03152530507626086, 32'sd-0.12753002275874575, 32'sd0.01820523248458226, 32'sd0.0149097081326442, 32'sd0.11212352262841738, 32'sd0.09920254675987793, 32'sd0.06423216605703629, 32'sd0.06179026982602176, 32'sd0.04428182736738433, 32'sd-0.08187230352045226, 32'sd-0.08472189737229815, 32'sd-0.020790868039142357, 32'sd-0.10025962711690972, 32'sd-0.002721265902003905, 32'sd-0.004293872326299041, 32'sd0.08220209981827047, 32'sd0.0005713047733506212, 32'sd0.03366139665164832, 32'sd-0.060207446339486326, 32'sd-0.03444481756752105, 32'sd0.05684306456462961, 32'sd0.04169833837041521, 32'sd-0.05098582559276378, 32'sd0.06994844232941799, 32'sd0.0615115483738589, 32'sd0.0952987306835173, 32'sd-0.14329299995712277, 32'sd0.09945501652546335, 32'sd0.028108032293090234, 32'sd0.0698026833653867, 32'sd0.014814171147003636, 32'sd-0.031800909592855926, 32'sd-0.012605331730072599, 32'sd0.10170704403002974, 32'sd0.04614317100167204, 32'sd0.07137567545624655, 32'sd0.17181294174073122, 32'sd-0.02892223424709915, 32'sd0.07894249081165704, 32'sd-0.1508913631843751, 32'sd-0.033827767608362126, 32'sd-0.04348933334372733, 32'sd-0.015273389781083242, 32'sd0.14766210338729777, 32'sd0.0551939685719052, 32'sd0.09415032326869595, 32'sd0.036015753673609804, 32'sd0.03988618088974947, 32'sd0.013414905038917064, 32'sd-0.04388547493756252, 32'sd0.019393715170522737, 32'sd0.019038196134416718, 32'sd-0.08912556874193911, 32'sd0.12605149479310768, 32'sd-0.11073895441865371, 32'sd0.00574700772788341, 32'sd0.12990645087576533, 32'sd0.13145922414801142, 32'sd0.007152414910679823, 32'sd-0.020909193213680403, 32'sd-0.04931488280914053, 32'sd0.15176738930422742, 32'sd0.006754212862955271, 32'sd0.0700388502226342, 32'sd0.11900751516062848, 32'sd0.1212786522843734, 32'sd-0.018601009784540667, 32'sd-0.14831999883677816, 32'sd-0.06324477649867485, 32'sd0.05388822564536455, 32'sd0.013103192755518417, 32'sd0.0428497515847595, 32'sd0.18001496102596776, 32'sd-0.069667358153465, 32'sd-0.05480756872265021, 32'sd-0.06109575826374057, 32'sd-0.02338997517093748, 32'sd-0.020079573728203633, 32'sd0.05490304211256897, 32'sd-0.052265843901230034, 32'sd-0.06470747624724513, 32'sd0.013398873866179838, 32'sd0.048971976600614246, 32'sd0.06612471889954094, 32'sd0.06987779603574676, 32'sd0.1690304320845407, 32'sd0.08919468824567744, 32'sd-0.007818868885267312, 32'sd0.014219758935723572, 32'sd0.10051825064410526, 32'sd0.11087442991418779, 32'sd0.032442423321863936, 32'sd0.1379921220299337, 32'sd0.14556415122779898, 32'sd0.14944482134909923, 32'sd-0.0654407600321147, 32'sd-0.02162495627537016, 32'sd0.025816720857201533, 32'sd-0.010323834675805495, 32'sd0.025283839609051204, 32'sd0.05399717870174714, 32'sd-0.016216865456038426, 32'sd-0.011808102572275613, 32'sd-0.2771545776568999, 32'sd0.022430919176628202, 32'sd-0.006268174937176653, 32'sd1.0285599034628197e-121, 32'sd-0.0034540221070124347, 32'sd-0.046156262716311285, 32'sd-0.09059746520514692, 32'sd-0.04970848254948598, 32'sd-0.022431998489370667, 32'sd0.01015924761367918, 32'sd0.04189804531797617, 32'sd-0.026513713120645307, 32'sd-0.002910707631887586, 32'sd-0.09468833276138315, 32'sd-0.11207822605478542, 32'sd0.0023420615590794766, 32'sd0.1823552156849123, 32'sd0.18683276628258538, 32'sd0.0852306011241166, 32'sd0.1373265155811292, 32'sd-0.03692620578369532, 32'sd-0.07615442799300787, 32'sd-0.06320971456377668, 32'sd0.10466194116763272, 32'sd0.10749243881304163, 32'sd0.061487796574556955, 32'sd0.031212407097412333, 32'sd-0.013518366693692638, 32'sd-0.05636347439826637, 32'sd0.029701965072598303, 32'sd-0.004960070936730702, 32'sd-0.03659400682994207, 32'sd-0.05937752731679588, 32'sd0.05085340801263176, 32'sd-0.02252893595989649, 32'sd0.07450287116173497, 32'sd-0.07192222991507352, 32'sd-0.1118687824781098, 32'sd-0.04460424476847168, 32'sd-0.021402789784997503, 32'sd-0.06618377292477999, 32'sd-0.04249937619596701, 32'sd-0.04184560335623085, 32'sd0.06233932799660811, 32'sd0.1957114445633278, 32'sd0.019305979887610406, 32'sd-0.07443734666211374, 32'sd-0.04446636608741356, 32'sd-0.05703094249109917, 32'sd0.043376416063720495, 32'sd-0.1166320877675149, 32'sd0.09324320658179146, 32'sd0.106958426494475, 32'sd-0.005926143469283112, 32'sd-0.05083617841016818, 32'sd-0.0802685215177227, 32'sd-0.11628028671063083, 32'sd-0.04549411347952426, 32'sd-0.08039154413078385, 32'sd0.01352950840207017, 32'sd0.059982371849388004, 32'sd-0.05809769582643284, 32'sd0.04118284732280835, 32'sd0.08070412063655212, 32'sd-0.12030853839234959, 32'sd0.01791412230894292, 32'sd0.005429536497668188, 32'sd-0.10584589740684236, 32'sd0.03578769423449487, 32'sd-0.08909841273558629, 32'sd0.08277786111709161, 32'sd0.04229604511585986, 32'sd0.06810830785901782, 32'sd-0.0421748018854318, 32'sd-0.03169491449706669, 32'sd0.022217282978352338, 32'sd-0.009431918847162305, 32'sd0.027673006365834942, 32'sd-0.05020927625706961, 32'sd0.04156499798527987, 32'sd-0.0022450486041208847, 32'sd0.11729656468589504, 32'sd-0.015068577128983001, 32'sd-0.10572700456380785, 32'sd-0.015879987896991833, 32'sd0.034223699001492816, 32'sd0.010068531457027801, 32'sd5.696161856799976e-125, 32'sd0.039758687381227904, 32'sd-0.038076112454789125, 32'sd-0.029358022962390592, 32'sd-0.029327254298422586, 32'sd-0.034029574018469094, 32'sd-0.010776879456897731, 32'sd-0.04270616827501988, 32'sd-0.05031647073545708, 32'sd-0.030712461428864156, 32'sd-0.07846901795942159, 32'sd0.061675012688598756, 32'sd-0.002865524307943089, 32'sd0.10992527564423388, 32'sd0.06953633763693329, 32'sd-0.046074484493152164, 32'sd0.022196601991634462, 32'sd0.01664732740045206, 32'sd0.07026433151062667, 32'sd0.038026809739852986, 32'sd-0.04955955106127373, 32'sd0.010428784197155485, 32'sd0.048295998334655116, 32'sd-0.07192077270062792, 32'sd-0.04237671394165172, 32'sd-0.05274680784991379, 32'sd0.037817222131726745, 32'sd-0.021748529562861, 32'sd0.021063096191903344, 32'sd-0.08754511048990439, 32'sd-0.015245517586501174, 32'sd0.02577600404209846, 32'sd-0.049706226394989575, 32'sd0.032904839099362614, 32'sd-0.04121553326358029, 32'sd-0.0700180391839791, 32'sd-0.04082323539248676, 32'sd0.0046504758268477815, 32'sd0.07154794896576178, 32'sd-0.05217375010396391, 32'sd-0.010353057031685868, 32'sd-0.037687252497379024, 32'sd0.1285164809396347, 32'sd-0.05451043018852416, 32'sd-0.012279715074955634, 32'sd0.007553905681999045, 32'sd-0.02576538406186785, 32'sd-0.047191722434421164, 32'sd-0.043773561093799915, 32'sd0.011320053724105543, 32'sd0.045657748251656194, 32'sd0.03803389230946219, 32'sd-0.05951811918919387, 32'sd-0.014064253779868278, 32'sd0.056362513982465993, 32'sd-0.009321493880659828, 32'sd-0.06514680015032641, 32'sd-0.018917477731813726, 32'sd-0.03240156620916565, 32'sd0.05674734911421235, 32'sd0.02493858589164401, 32'sd0.06262004463150342, 32'sd-0.07873162986922731, 32'sd-0.0798033476707356, 32'sd0.0481957274331425, 32'sd-0.07321407279289241, 32'sd0.027141312649304868, 32'sd-0.10279471837017767, 32'sd0.018210914495056924, 32'sd-0.00037817461295594756, 32'sd-0.03434138880241771, 32'sd0.0099329823972103, 32'sd-0.06027041028348383, 32'sd-0.03571936455141734, 32'sd0.08773644965469979, 32'sd-0.06118380126786906, 32'sd0.03373445660840265, 32'sd-0.07102153081624776, 32'sd0.10169709759600076, 32'sd-0.07539529812257063, 32'sd0.03197393518557943, 32'sd-0.020097568957520594, 32'sd-0.015745865803207814, 32'sd0.00041156264351051373, 32'sd-1.6469077499154087e-125, 32'sd0.024184632355428063, 32'sd0.024091855693139094, 32'sd0.13466977465218524, 32'sd0.006595668726852535, 32'sd-0.05278706074305672, 32'sd-0.045855871235971096, 32'sd0.000974815352484912, 32'sd-0.04094134597558885, 32'sd0.0351056307983432, 32'sd0.11870285938619632, 32'sd-0.04332404802761271, 32'sd-0.08570128845687017, 32'sd0.09022954760097869, 32'sd0.05359485687308124, 32'sd0.0042578331176544035, 32'sd-0.14481823645403766, 32'sd-0.09957416283355583, 32'sd-0.024259140197670316, 32'sd0.040628096285589416, 32'sd-0.09509237059684841, 32'sd-0.1201504555429973, 32'sd-0.09655363873831485, 32'sd0.02149853625371348, 32'sd-0.09977452577574152, 32'sd-0.04261253334240924, 32'sd0.08637274895983904, 32'sd-4.578687287439892e-127, 32'sd8.790335210950298e-122, 32'sd-1.3091305315731472e-118, 32'sd0.08015395989472757, 32'sd-0.011747632270812254, 32'sd0.07188803344382388, 32'sd-0.16383605239798882, 32'sd0.03517535338500673, 32'sd0.013242487485942705, 32'sd0.014969432039049189, 32'sd0.07819859135671443, 32'sd0.15858341262194214, 32'sd0.09714200198552288, 32'sd-0.03146680969198326, 32'sd-0.039041858833476564, 32'sd-0.03389564583020014, 32'sd0.004858733904347035, 32'sd-0.0556143806304909, 32'sd-0.05721672898209715, 32'sd-0.05978782843680459, 32'sd0.011671458955410946, 32'sd-0.09916903865458084, 32'sd0.05241806232088563, 32'sd0.07665335761316137, 32'sd-0.04266459010565457, 32'sd0.06758569781989855, 32'sd-0.028751535139010166, 32'sd0.014313848911291033, 32'sd1.6321844158548605e-115, 32'sd1.898317398913079e-115, 32'sd-1.1131229832301632e-122, 32'sd0.011082272142956947, 32'sd0.02339974032063824, 32'sd-0.09898253737797855, 32'sd-0.010789823977807821, 32'sd0.015702083513808602, 32'sd0.1418411489098301, 32'sd0.15673394575448546, 32'sd0.06679821861156365, 32'sd0.10005225966351486, 32'sd0.02274720421505338, 32'sd0.08241110567939963, 32'sd0.030860410931039015, 32'sd-0.11628541416683229, 32'sd-0.06801892077304995, 32'sd-0.009782550794275998, 32'sd-0.023629613694299927, 32'sd-0.014590315047491796, 32'sd-0.1016925052147245, 32'sd-0.16060907652722556, 32'sd-0.08479683947730939, 32'sd-0.04033324353472562, 32'sd0.1045375813282515, 32'sd-0.04297517567728186, 32'sd-0.04170922236340387, 32'sd0.00400633089555955, 32'sd1.6327561627176686e-115, 32'sd-3.101104597714936e-120, 32'sd-1.8147908889095266e-123, 32'sd-4.327735419898538e-118, 32'sd0.010281494428543357, 32'sd-0.030956147643621028, 32'sd0.02383979269681942, 32'sd0.015833216310981814, 32'sd-0.08058211058407214, 32'sd-0.041592332656299795, 32'sd0.006982020214029135, 32'sd0.019591098748826533, 32'sd-0.006765404427769608, 32'sd-0.026700976240097447, 32'sd0.03950411543978073, 32'sd-0.010766269895924753, 32'sd-0.11429016065244661, 32'sd-0.04288643704204652, 32'sd-0.016848378128824993, 32'sd-0.010397574444064112, 32'sd-0.051540760631927994, 32'sd-0.10391958704180061, 32'sd-0.012455511099933453, 32'sd-0.0026405702739379228, 32'sd-0.045330292560700876, 32'sd0.003876075691389484, 32'sd0.03808539547434374, 32'sd1.6326989856482265e-123, 32'sd-7.499763566834906e-115, 32'sd-8.001580285212484e-116, 32'sd9.807204949724801e-122, 32'sd-2.6148835288386578e-126, 32'sd2.4241306176602217e-127, 32'sd0.006230807492825501, 32'sd0.012976126381937944, 32'sd-0.008486509323368167, 32'sd0.06125935178653376, 32'sd0.04760874246780555, 32'sd0.06507393631101026, 32'sd-0.09418061297945496, 32'sd-0.010060779010124704, 32'sd-0.07506444987966232, 32'sd-0.08036417644037684, 32'sd-0.13883019176803177, 32'sd0.024591230109741468, 32'sd0.024102730157711246, 32'sd-0.02316862044306833, 32'sd-0.039821341015616726, 32'sd-0.08468670771959408, 32'sd0.010028353045379535, 32'sd0.003377094137685695, 32'sd0.004849209982399971, 32'sd0.10395236878216159, 32'sd-9.421608171440139e-116, 32'sd2.5971025864341656e-118, 32'sd-5.921449011382963e-127, 32'sd1.6051423511205485e-115},
        '{32'sd-4.437543529858713e-115, 32'sd-3.2558733319443777e-116, 32'sd-4.244403054632222e-125, 32'sd-1.7651587291619054e-127, 32'sd1.6721528522988766e-117, 32'sd2.2614245320258196e-115, 32'sd1.1377173792937832e-123, 32'sd1.2939584173503119e-126, 32'sd4.539673189257243e-121, 32'sd4.3292529509010127e-125, 32'sd-2.5586630458722978e-126, 32'sd-5.411835001633417e-117, 32'sd0.08575117210194999, 32'sd0.1065622833852017, 32'sd-0.06737922699074943, 32'sd0.06780818351652251, 32'sd9.516694262025198e-119, 32'sd-5.17337818784904e-120, 32'sd6.400864068063665e-125, 32'sd7.064620544082441e-121, 32'sd1.8166739580484716e-120, 32'sd-2.9013569397809034e-125, 32'sd-1.0938738453855398e-125, 32'sd8.62975442872328e-117, 32'sd-1.2856695285777947e-125, 32'sd3.428886419069733e-116, 32'sd-3.5447689468493914e-119, 32'sd-1.352493985099412e-119, 32'sd3.6406869514690196e-116, 32'sd-2.712422879660753e-124, 32'sd3.114593812940831e-120, 32'sd-2.114387586917288e-127, 32'sd0.047532333812404695, 32'sd0.03333957695615232, 32'sd0.0016227557441907054, 32'sd-0.11584168946268808, 32'sd-0.06726803018827754, 32'sd-0.08232310213488046, 32'sd-0.0005211478130568259, 32'sd-0.05219776431840679, 32'sd0.08920810772095882, 32'sd0.046839921093789316, 32'sd-0.012044226883301926, 32'sd0.02015903162157322, 32'sd-0.03156650605139294, 32'sd0.06043814542254752, 32'sd0.03362586229893696, 32'sd0.05404348071078259, 32'sd0.01774518693821996, 32'sd0.1044588988730558, 32'sd0.05904694392836909, 32'sd0.0070584676185305615, 32'sd2.718044693250886e-128, 32'sd-8.263736636656962e-126, 32'sd3.9501209682427386e-119, 32'sd9.61957453024479e-128, 32'sd3.955887268313633e-119, 32'sd4.378695685738467e-121, 32'sd0.08793903447092209, 32'sd-0.04107269317214375, 32'sd0.0820260291956841, 32'sd0.02131166688313016, 32'sd-0.11028479883701728, 32'sd-0.056786646118441024, 32'sd-0.04151498424776613, 32'sd0.046813406422931234, 32'sd-0.07119899783955792, 32'sd0.0778038119007951, 32'sd0.10230453651153018, 32'sd0.0864075803483067, 32'sd0.01640016937861611, 32'sd0.1840729729903146, 32'sd0.14945946984780026, 32'sd0.040023170793662945, 32'sd0.05942486818685603, 32'sd-0.02452559528120526, 32'sd-0.017207861422364946, 32'sd0.017275004944395617, 32'sd-0.015975906213595802, 32'sd-0.026207157699786855, 32'sd0.13629464730550586, 32'sd0.06449382606636295, 32'sd-9.829830623898489e-124, 32'sd-3.9192850291237155e-123, 32'sd3.2201748130561273e-128, 32'sd1.6388549385812836e-124, 32'sd-0.030875344592512326, 32'sd0.09372717834784347, 32'sd-0.01400373073027289, 32'sd-0.0014737856245693518, 32'sd-0.07838026814329907, 32'sd-0.06977345094431522, 32'sd0.03914072217526083, 32'sd-0.03258305258929128, 32'sd0.04638316052288613, 32'sd0.0323529389371228, 32'sd-0.017075375597839813, 32'sd0.07609978603586627, 32'sd0.046924173051834266, 32'sd0.09128598443200815, 32'sd0.09415368301652893, 32'sd0.1471722498333153, 32'sd0.06906563012084976, 32'sd0.2051853748089016, 32'sd-0.006224571967358662, 32'sd-0.040795279672157944, 32'sd-0.06915721911576, 32'sd-0.023084873893463594, 32'sd0.0007404842513437219, 32'sd-0.02074349791918986, 32'sd0.04244711924096166, 32'sd-3.2782683473821034e-116, 32'sd-1.24658595409523e-118, 32'sd0.06198368714927454, 32'sd0.07409411496978532, 32'sd-0.0233239874345014, 32'sd0.06501598976467671, 32'sd-0.003554338295449791, 32'sd-0.16148978922598628, 32'sd-0.043673528844798984, 32'sd0.0014140918700564194, 32'sd-0.022307553077959556, 32'sd-0.01611586562796273, 32'sd-0.058450752580436, 32'sd0.07124589964348482, 32'sd0.034703122886034374, 32'sd0.07564618570218572, 32'sd-0.029310720444487633, 32'sd-0.0723476014487638, 32'sd-0.020740338445968915, 32'sd0.09789516247212149, 32'sd-0.014986925427446519, 32'sd-0.04942658267012434, 32'sd0.09736176904532222, 32'sd0.04657125467642357, 32'sd0.01956329793692664, 32'sd0.041785709459177055, 32'sd-0.06878254263087938, 32'sd-0.06339458547743415, 32'sd-0.05203129045047554, 32'sd1.5038657503062285e-124, 32'sd0.08014398142920527, 32'sd-0.024175562352553664, 32'sd-0.03398336748566694, 32'sd0.024001603263086584, 32'sd0.00568437401131823, 32'sd-0.08630669225628274, 32'sd-0.002069146805129799, 32'sd0.017511562737064397, 32'sd0.014375117269763961, 32'sd0.01410250986932588, 32'sd0.010848847368314417, 32'sd-0.07273132598524203, 32'sd0.051157921175401515, 32'sd0.10540831787702142, 32'sd0.06869629410446654, 32'sd0.09478576275536026, 32'sd-0.011572923972416055, 32'sd0.05865929085324801, 32'sd-0.04697521921339476, 32'sd-0.036008157040454646, 32'sd-0.027876689449136592, 32'sd-0.08007360800686557, 32'sd0.034341815380795705, 32'sd-0.01046845226686587, 32'sd0.029731201972363567, 32'sd0.04451993134889433, 32'sd0.07394853035333024, 32'sd1.2369449659236253e-123, 32'sd0.06621307872168064, 32'sd-0.010386870764598984, 32'sd-0.07263374649065067, 32'sd0.017315696683475698, 32'sd0.00044584241857879283, 32'sd-0.10881453180097508, 32'sd-0.1410285767050505, 32'sd-0.22133276138239458, 32'sd-0.04103260890491394, 32'sd-0.09630068882032568, 32'sd0.01075445684299972, 32'sd0.05310296853873524, 32'sd0.04878953417012709, 32'sd0.02345123240217805, 32'sd0.004059096823987864, 32'sd-0.0482588650556846, 32'sd-0.051030558544928176, 32'sd0.08559955288762036, 32'sd0.00457490895009454, 32'sd0.01202116995304704, 32'sd0.06268766357332621, 32'sd-0.08458712964066088, 32'sd-0.01260903734688571, 32'sd-0.039823290284823544, 32'sd-0.006597756395001554, 32'sd0.10344725999472437, 32'sd-0.016986935858313356, 32'sd0.04056210071850352, 32'sd-0.043067841702831525, 32'sd0.06678943335289042, 32'sd-0.012750244540399904, 32'sd-0.03845504637204318, 32'sd-0.09931118641321235, 32'sd-0.09220023447128135, 32'sd-0.007534195492569743, 32'sd-0.1631484451118228, 32'sd-0.03717834703687816, 32'sd-0.0218616601098546, 32'sd-0.0580171058181488, 32'sd0.034320739021019314, 32'sd-0.00878811665274987, 32'sd0.08050420060112447, 32'sd-0.13222029182658382, 32'sd-0.03389761048447598, 32'sd-0.0023606700096701905, 32'sd-0.07702905707105735, 32'sd-0.04384801721779918, 32'sd-0.015989153723940972, 32'sd0.03419850103095896, 32'sd0.01749377983663714, 32'sd-0.040730803922719605, 32'sd-0.10351787554382318, 32'sd-0.06850310083734314, 32'sd0.10722785831169367, 32'sd0.0029595362356050494, 32'sd0.06346882574841745, 32'sd-0.00704275757484986, 32'sd-0.07810055545664907, 32'sd0.06140009999138834, 32'sd0.031350723447516826, 32'sd-0.03428494378786125, 32'sd0.006008516419461783, 32'sd0.028814858106251208, 32'sd-0.10198459694593416, 32'sd-0.05082464644886267, 32'sd-0.11753093653984613, 32'sd-0.1650552046116974, 32'sd-0.060128235523937194, 32'sd-0.025315187042827432, 32'sd0.067574289850384, 32'sd-0.04980718211192651, 32'sd-0.13255894893020803, 32'sd0.046860807161318505, 32'sd-0.1652482923303478, 32'sd-0.04183655174547321, 32'sd-0.09454970056668094, 32'sd-0.1192335674108213, 32'sd-0.11766016981992865, 32'sd-0.030434656710677122, 32'sd-0.05665614183326734, 32'sd-0.1172702054428584, 32'sd0.10125759696851959, 32'sd-0.02137168582484497, 32'sd0.10975278657541403, 32'sd-0.010515939902433689, 32'sd-0.028535329226314157, 32'sd-0.02389306890525429, 32'sd0.10495927277648492, 32'sd0.014493894764539213, 32'sd0.05072293481770349, 32'sd0.08239588184638183, 32'sd-0.036593153691170305, 32'sd-0.15220230309218447, 32'sd-0.25842161691271104, 32'sd-0.1666585188860931, 32'sd0.030077553534193044, 32'sd0.07928950675586309, 32'sd0.08420973565874845, 32'sd0.0552908699584154, 32'sd0.042919842659819116, 32'sd-0.06299105656692434, 32'sd-0.13654050969862497, 32'sd-0.07342102401939558, 32'sd-0.09520005068048516, 32'sd-0.15616926624395971, 32'sd-0.1215186965037824, 32'sd-0.08278193658504274, 32'sd-0.038615766787813297, 32'sd-0.07364958103107618, 32'sd0.09140580528135435, 32'sd0.03591320612242501, 32'sd0.00863211938705501, 32'sd0.1140379859167465, 32'sd-0.10372272742068256, 32'sd-0.06764662394156663, 32'sd0.018350790255589153, 32'sd-0.01183329302999957, 32'sd0.11010663433095597, 32'sd-0.011889699423793665, 32'sd-0.08146714319460804, 32'sd-0.07107111919821389, 32'sd-0.1276348047390007, 32'sd-0.09676213566570593, 32'sd0.03436517320954388, 32'sd0.17100220472470515, 32'sd0.17403986580776562, 32'sd0.13485792165485266, 32'sd0.06196467570817175, 32'sd-0.0013073983367392322, 32'sd-0.03391163653080303, 32'sd-0.11538418514968808, 32'sd-0.11053984064962696, 32'sd-0.04997741631441704, 32'sd-0.0883772906393006, 32'sd-0.17201161233221476, 32'sd-0.014536339187612752, 32'sd-0.09536373032510877, 32'sd0.08210226511317252, 32'sd-0.015832578574850438, 32'sd0.01126275390907708, 32'sd0.0026244444467676494, 32'sd-0.18222052009610815, 32'sd-0.09617058632548774, 32'sd0.056565393884258, 32'sd0.013080232008803275, 32'sd-0.00819842385000375, 32'sd0.03375210023639083, 32'sd-0.10463937876310381, 32'sd-0.16589180234374018, 32'sd-0.15244293275490153, 32'sd-0.002200766281882942, 32'sd0.1380497016994123, 32'sd0.12656857296848922, 32'sd0.15575536192071596, 32'sd0.13142974916548558, 32'sd-0.10854942321661011, 32'sd-0.12958615791150488, 32'sd-0.08488560474652788, 32'sd0.04463731014115427, 32'sd-0.06355032156787889, 32'sd-0.06989572120796088, 32'sd-0.08236275249731898, 32'sd-0.12087886000419164, 32'sd-0.18960468590436114, 32'sd0.012350326894412574, 32'sd0.07248118895030664, 32'sd-0.02205042391694274, 32'sd0.027322202568141607, 32'sd-0.08646390315272189, 32'sd0.04203016814295714, 32'sd0.025930820262395977, 32'sd0.07004899686205904, 32'sd0.015298061966650785, 32'sd-0.09233962920826491, 32'sd-0.14727068576175448, 32'sd-0.20712471028106, 32'sd-0.05685787884748027, 32'sd0.10204434540295744, 32'sd0.047785656660352435, 32'sd0.1765977853758489, 32'sd0.14234388585719207, 32'sd0.07662387549010624, 32'sd0.14189341602638914, 32'sd-0.06264815910602853, 32'sd-0.033680425487371705, 32'sd0.018919296951540175, 32'sd0.07881784966674961, 32'sd-0.04329849555441478, 32'sd0.053635406910324215, 32'sd-0.08650885666729305, 32'sd0.0803961740941489, 32'sd-0.01718205913799916, 32'sd-0.09159400144467587, 32'sd-0.08339796423104122, 32'sd-0.10494380865913865, 32'sd0.014498013577437416, 32'sd-0.0027064287434550214, 32'sd-0.0161922581405879, 32'sd0.06498742782366765, 32'sd0.0040990524488189305, 32'sd0.10168360508628405, 32'sd0.012221214503873767, 32'sd0.00414763436188949, 32'sd-0.04983305335300482, 32'sd0.04538047779722873, 32'sd0.1596838468010156, 32'sd0.06053333955828012, 32'sd-0.02199920916382837, 32'sd-0.03181726106966144, 32'sd0.02832907631060284, 32'sd0.07535434111168987, 32'sd0.009656857511820105, 32'sd0.052383515598196054, 32'sd0.02093979288051314, 32'sd0.1213855079101391, 32'sd0.11577265529572657, 32'sd0.09497391029808122, 32'sd-0.00771353932944967, 32'sd0.1267286886593869, 32'sd0.007495467555705471, 32'sd-0.10336759092047892, 32'sd-0.037441771656405214, 32'sd0.004749189357602659, 32'sd0.11499220175499622, 32'sd-0.01122175011835404, 32'sd0.014406227403551524, 32'sd0.048389210409218904, 32'sd-0.021089092684946152, 32'sd-0.012143922667162152, 32'sd0.0537491747657098, 32'sd-0.11606209088074373, 32'sd-0.04286077498899437, 32'sd-0.02083187131296445, 32'sd0.16718390917116277, 32'sd0.07749129320878462, 32'sd0.053924970203834736, 32'sd0.0399526584719878, 32'sd0.060420702722137794, 32'sd-0.08194647456554903, 32'sd0.04076250190509616, 32'sd-0.004896852868882634, 32'sd0.06942349545102526, 32'sd0.18393836396315982, 32'sd0.03557651966156944, 32'sd0.1620024000163422, 32'sd0.09224743922313386, 32'sd0.13627569108066756, 32'sd-0.006130804285720795, 32'sd-0.04340839465383473, 32'sd-0.14018138787631662, 32'sd0.015857103415154776, 32'sd0.09345894912434571, 32'sd-0.06710349950033481, 32'sd-0.02782398108263261, 32'sd-0.04137151483858111, 32'sd-0.03190815766388177, 32'sd0.0010199237575940724, 32'sd0.10633417041726223, 32'sd0.09298456096555255, 32'sd-0.004719608551025081, 32'sd0.012108111957050737, 32'sd0.11062247315722203, 32'sd0.04329040094189429, 32'sd0.005799220383364995, 32'sd-0.023874666603640928, 32'sd0.01646056011493708, 32'sd-0.04416661806246755, 32'sd-0.03487822104712312, 32'sd0.06498173087043192, 32'sd0.1562139856633706, 32'sd0.17399687884085183, 32'sd0.08878997851182752, 32'sd0.06412240083702625, 32'sd0.1060870621946182, 32'sd0.17010885648742388, 32'sd0.04536815536501983, 32'sd-0.03686347578888971, 32'sd-0.012818318901113835, 32'sd0.013138492122995959, 32'sd-0.022133320151785683, 32'sd0.006869314968328177, 32'sd0.035991192253046284, 32'sd-0.03931518168978359, 32'sd-0.03756165487903661, 32'sd-0.08547157910073788, 32'sd0.034579930029707884, 32'sd0.15549395566748608, 32'sd0.08942754919241752, 32'sd0.057431493469120465, 32'sd0.09501406114454812, 32'sd0.07917434352083236, 32'sd0.04569863806590583, 32'sd0.05060777533986875, 32'sd-0.014555955873378257, 32'sd-0.042647669331823845, 32'sd0.040345659053191256, 32'sd-0.05503798033775504, 32'sd0.1220003912063561, 32'sd0.10673358369584356, 32'sd0.007660669739560361, 32'sd0.15314954942626266, 32'sd0.006875936033502677, 32'sd0.04299681095247933, 32'sd0.07344536197749292, 32'sd-0.17421076820399664, 32'sd0.048447247408766984, 32'sd0.049183100246652796, 32'sd1.742681320303349e-125, 32'sd0.045259335931102214, 32'sd-0.019466600273882327, 32'sd0.007559178127802824, 32'sd0.1657377238493002, 32'sd0.041161623153326506, 32'sd0.007574693113675878, 32'sd0.08887364846234569, 32'sd-0.01007339264631237, 32'sd-0.06374775053103215, 32'sd0.048799274641631064, 32'sd-0.06536851549910644, 32'sd-0.05954008208291167, 32'sd0.015239777492834191, 32'sd0.041040663746945434, 32'sd-0.12183681954776676, 32'sd0.10926504121518012, 32'sd0.01671637827029966, 32'sd-0.04530227739019646, 32'sd-0.0006305499691026954, 32'sd0.05310583606467463, 32'sd0.10875781320570736, 32'sd0.01808202035801339, 32'sd0.05979876824456472, 32'sd0.035372598065781705, 32'sd-0.06216445520446194, 32'sd0.08267607308358256, 32'sd-0.09874417962656275, 32'sd-0.039157383566968774, 32'sd0.03388960665085615, 32'sd-0.07682491381594213, 32'sd0.06913807735678272, 32'sd0.071014800074612, 32'sd-0.00883376090857932, 32'sd0.00034618296155003306, 32'sd0.05440048547135551, 32'sd-0.09119441833535206, 32'sd-0.00943425799474693, 32'sd-0.04294063194562684, 32'sd-0.09666111408523484, 32'sd-0.10200625369586815, 32'sd0.16541721364804401, 32'sd0.039109846348599576, 32'sd0.010596265439573092, 32'sd-0.04287739726189563, 32'sd-0.03071844313636728, 32'sd-0.011906034008847897, 32'sd0.01936945346547157, 32'sd-0.0582462062323059, 32'sd-0.012208241082769794, 32'sd0.03469724468331806, 32'sd-0.1179799954817582, 32'sd-0.03586970303980669, 32'sd-0.02957423986855246, 32'sd0.08460827458806973, 32'sd-0.01201938238053485, 32'sd0.022172153754593214, 32'sd0.02506920367876053, 32'sd-0.045492523794788506, 32'sd-0.018200947342438257, 32'sd0.016070118008829067, 32'sd0.016088551566068032, 32'sd0.007497171233313918, 32'sd-0.05055162181360676, 32'sd-0.1378593231875074, 32'sd0.12492286835529365, 32'sd-0.10117342903953852, 32'sd-0.058541544408927455, 32'sd0.13598326852253992, 32'sd0.05390770318587008, 32'sd-0.015587324220465127, 32'sd0.03593165410247246, 32'sd-0.025522640683715053, 32'sd-0.036684226047758686, 32'sd0.04874537947832786, 32'sd0.005214675453846664, 32'sd-0.08989917681840572, 32'sd-0.06527121436186953, 32'sd-0.12609744302565387, 32'sd-0.0900066135860673, 32'sd-0.08989541642674378, 32'sd-0.13227323948343991, 32'sd-0.039090196854559375, 32'sd-0.028099020906707656, 32'sd-1.9905235074006132e-122, 32'sd-0.0429172063410837, 32'sd0.012304217989269303, 32'sd-0.022134945023146144, 32'sd-0.002478578962223205, 32'sd-0.0016809310811578345, 32'sd-0.025234906566412207, 32'sd-0.0062645271588115895, 32'sd-0.10306272479170756, 32'sd-0.05250937709727794, 32'sd-0.012371136089011043, 32'sd0.04233184150158807, 32'sd0.01040400684793132, 32'sd0.1588067673342434, 32'sd0.09945651896603237, 32'sd0.09279234813605904, 32'sd0.1307582808785914, 32'sd-0.12762186064248054, 32'sd0.05441954857271771, 32'sd-0.12877857683569127, 32'sd-0.009490514568031214, 32'sd-0.0761868786567945, 32'sd-0.08124198744495971, 32'sd-0.14697896727267035, 32'sd-0.08283054863809276, 32'sd-0.11547954566988845, 32'sd0.06457257286911965, 32'sd-0.021625188383725617, 32'sd0.07730057089631334, 32'sd0.06917510641957927, 32'sd0.053456688716231555, 32'sd-0.11022899020057557, 32'sd-0.09733391317560537, 32'sd-0.10391573925802579, 32'sd-0.047710573025289964, 32'sd-0.06983204399898701, 32'sd-0.03807597725844324, 32'sd-0.07416473174004243, 32'sd-0.015758095538732402, 32'sd-0.0016532406057666379, 32'sd0.03475631257169453, 32'sd0.011909153779230979, 32'sd0.0965294336355672, 32'sd0.09301296169195467, 32'sd0.11572346658695018, 32'sd0.013910861419709184, 32'sd0.07902946183705253, 32'sd-0.01442860335369392, 32'sd-0.09676501085103367, 32'sd-0.16851925805176832, 32'sd-0.09400959633700921, 32'sd-0.0641770651672579, 32'sd0.0154152669638936, 32'sd0.007739953212163087, 32'sd0.059658170698083685, 32'sd0.007385233759701466, 32'sd-0.0013634830062224125, 32'sd0.09033858536710974, 32'sd0.06839953434264094, 32'sd-0.03301775975823738, 32'sd-0.07687726789559714, 32'sd0.05030499192554051, 32'sd-0.09716399465612914, 32'sd-0.11386449571224735, 32'sd-0.07706409404525669, 32'sd-0.12638105045844872, 32'sd-0.001881283041987939, 32'sd0.007625865301164559, 32'sd0.02003904354444908, 32'sd0.005698693734718884, 32'sd-0.04704004786415476, 32'sd0.00435441452470046, 32'sd0.04238905932526317, 32'sd-0.06140466270142148, 32'sd-0.056688212698435006, 32'sd-0.05419207542505063, 32'sd-0.020730705308166474, 32'sd-0.06425930622892008, 32'sd0.05379575947479837, 32'sd-0.07267488265537346, 32'sd-0.10278386839441231, 32'sd-0.04306393989962402, 32'sd0.04815713015070464, 32'sd0.026633529024945594, 32'sd-3.117406216858371e-119, 32'sd0.08415358953412366, 32'sd0.009248109258695101, 32'sd0.08403364393063906, 32'sd0.08926945935847252, 32'sd0.05251084902021182, 32'sd0.026109814149465945, 32'sd0.03867400849871633, 32'sd0.0355223810840993, 32'sd0.07013732429591345, 32'sd0.07639378795923688, 32'sd0.14740258930673078, 32'sd0.05095710995062696, 32'sd0.0030174704151725573, 32'sd0.04379459559820684, 32'sd0.10082375216397696, 32'sd-0.07456643026530824, 32'sd-0.07482011052493995, 32'sd-0.09007100994809192, 32'sd0.02722276758713526, 32'sd-0.011469935815048677, 32'sd0.027819905312755074, 32'sd0.04224131629867278, 32'sd-0.04807999159470952, 32'sd-0.05692601606709492, 32'sd0.055968165156326403, 32'sd-0.06933126175629782, 32'sd-1.8168649295427094e-118, 32'sd-1.5426080310381822e-117, 32'sd9.582542308249074e-119, 32'sd-0.007560722069865412, 32'sd-0.0712461291080626, 32'sd-0.04335595868065368, 32'sd-0.03683939592076056, 32'sd-0.07763053812472068, 32'sd0.047764601671090784, 32'sd-0.08606209759673125, 32'sd0.12331689123453599, 32'sd-0.0017931403440280347, 32'sd0.0002452832423649679, 32'sd-0.04224012164550107, 32'sd-0.039215646265996586, 32'sd0.08651669113987899, 32'sd-0.0240160228854134, 32'sd-0.05091525839845884, 32'sd-0.06791092212430846, 32'sd-0.03790386044703106, 32'sd0.01787649177242615, 32'sd0.03706634289179638, 32'sd-0.09746612424371474, 32'sd-0.08360951033462616, 32'sd0.04818267209038439, 32'sd0.06671963053035128, 32'sd0.026247558426937757, 32'sd0.03449134999461185, 32'sd5.403931945340856e-118, 32'sd2.0477915650691097e-116, 32'sd-1.7856710534411967e-127, 32'sd0.008745550285686451, 32'sd0.028168473429295696, 32'sd0.10055946187496063, 32'sd0.061167108071018404, 32'sd0.08834098746006652, 32'sd0.07122081338444665, 32'sd-0.022479781428026663, 32'sd0.048192213590763415, 32'sd0.031583347749906766, 32'sd0.06879342491826772, 32'sd0.02754799156888008, 32'sd0.059845736094268735, 32'sd-0.11112938296043971, 32'sd0.00484046319763351, 32'sd0.0746274464470057, 32'sd-0.1197614550489032, 32'sd-0.023668382462639102, 32'sd-0.09577676048793175, 32'sd-0.09262423486915576, 32'sd-0.16080188802798856, 32'sd-0.11553516315428468, 32'sd0.017805135288466115, 32'sd0.030620464680078528, 32'sd0.025741737340471343, 32'sd0.07391726029997822, 32'sd-3.32558786538926e-119, 32'sd5.5265169492491644e-117, 32'sd-3.789032072368278e-122, 32'sd7.22805869668252e-121, 32'sd0.01841471477087464, 32'sd-0.12135768581067455, 32'sd-0.09988431624746259, 32'sd-0.021983196384663548, 32'sd-0.09612135681633438, 32'sd-0.18602714240786877, 32'sd-0.09475060335233977, 32'sd-0.007489820963477828, 32'sd0.01955878927318176, 32'sd-0.031120188187916578, 32'sd0.09602452498055986, 32'sd0.04684095728798938, 32'sd0.08985711658217005, 32'sd0.04811285119460857, 32'sd-0.045847946770936704, 32'sd-0.004959560057981941, 32'sd-0.022748475347677398, 32'sd-0.06172124802932529, 32'sd-0.08906946202970403, 32'sd-0.02008392136117461, 32'sd-0.03488241720998061, 32'sd0.027848399742621894, 32'sd0.06778642770442861, 32'sd3.6380073163598807e-127, 32'sd-2.2825981912440398e-114, 32'sd-1.8513258449223745e-126, 32'sd6.378767103167953e-126, 32'sd3.2744047851330604e-115, 32'sd-3.722116125764244e-125, 32'sd0.10201032512021073, 32'sd0.05855737785217699, 32'sd0.0016463503335921806, 32'sd0.058176293239903074, 32'sd-0.04722431661710732, 32'sd0.070693625475384, 32'sd-0.049520364428275974, 32'sd0.017258236178965804, 32'sd0.027533271161304766, 32'sd-0.027259727012996917, 32'sd0.09474177145217398, 32'sd-0.02152826149982896, 32'sd0.0065289075632612974, 32'sd0.00366379868861249, 32'sd-0.013471596365475501, 32'sd-0.09235126589641279, 32'sd0.0519716191653563, 32'sd-0.051032224385737734, 32'sd0.0250211537958253, 32'sd0.0023435269810829157, 32'sd1.7289628414606428e-125, 32'sd-3.631544093190946e-125, 32'sd-1.430338100957574e-123, 32'sd-3.407341775780303e-118},
        '{32'sd1.818644835710224e-123, 32'sd5.057569273165777e-118, 32'sd2.8773003188338535e-123, 32'sd-1.1596744686935125e-126, 32'sd-3.334065129054431e-116, 32'sd-6.893846140464742e-120, 32'sd6.3894227662575475e-115, 32'sd-1.104421364462367e-119, 32'sd-2.8590165901550036e-119, 32'sd-4.85139410630674e-123, 32'sd1.0911442932960038e-119, 32'sd-1.3404190765707564e-122, 32'sd0.030028427915950395, 32'sd-0.014598599421583017, 32'sd0.03264548369268323, 32'sd0.03844120743789293, 32'sd-2.070921212551198e-117, 32'sd-4.212553239259526e-126, 32'sd-2.215218662762347e-125, 32'sd3.1202801483966147e-119, 32'sd7.359022203807725e-122, 32'sd1.5428680843589896e-126, 32'sd-5.16416508921138e-122, 32'sd1.3333398506374e-123, 32'sd9.220011876999935e-125, 32'sd2.738883173390372e-125, 32'sd-2.2052323711579534e-121, 32'sd4.654375986673318e-115, 32'sd3.629636285951361e-114, 32'sd-1.7842169539410823e-123, 32'sd-1.5218708676212822e-125, 32'sd-2.2959533502775275e-126, 32'sd0.014310123619379061, 32'sd-0.03589846069407556, 32'sd-0.0557584398251688, 32'sd0.016355512985286858, 32'sd0.004026849549422332, 32'sd-0.056557943683382086, 32'sd0.047791364538919294, 32'sd0.03143713988436121, 32'sd-0.10193709777107231, 32'sd-0.05188828900086117, 32'sd-0.036467639973030916, 32'sd-0.05900289317485072, 32'sd0.06480618446967183, 32'sd-0.019264865982834205, 32'sd-0.019763595835658402, 32'sd0.0634510514152318, 32'sd-0.04036811335113243, 32'sd0.015140394829250212, 32'sd0.021774680546928195, 32'sd0.031170502440028065, 32'sd-5.835619853553475e-125, 32'sd-1.7237021675132928e-119, 32'sd1.7397291845570418e-125, 32'sd-3.9601771614640344e-119, 32'sd-2.53318596942371e-119, 32'sd3.0387440234830424e-127, 32'sd0.015907988503928674, 32'sd0.04567632826672663, 32'sd-0.004725831068877376, 32'sd0.008077427650985257, 32'sd0.07066746905196239, 32'sd-0.040544954728515714, 32'sd0.019506182104788748, 32'sd-0.003947646166217987, 32'sd0.013608656912021193, 32'sd0.07451051420954205, 32'sd-0.011858263873451588, 32'sd-0.05213123628672022, 32'sd-0.06579121724535869, 32'sd0.007718718254385378, 32'sd0.06771742243013881, 32'sd0.029076260019207066, 32'sd0.11442884768019358, 32'sd0.026600827255037852, 32'sd0.01535598409471233, 32'sd-0.015645441036157528, 32'sd0.07612389734865081, 32'sd0.011632530694573255, 32'sd0.013890944106731442, 32'sd0.03977560716892123, 32'sd4.8761633388785495e-120, 32'sd3.649889789635093e-122, 32'sd-5.863142101289702e-119, 32'sd6.137638468517629e-126, 32'sd0.06384537375958586, 32'sd0.034423837648647114, 32'sd0.024428076158564477, 32'sd0.032107459998130104, 32'sd0.06700143919254385, 32'sd0.05825233227835191, 32'sd0.06952635320996828, 32'sd0.038854458503048195, 32'sd0.10172509722109532, 32'sd0.06690305132198411, 32'sd0.18980559335315128, 32'sd0.12625817993550514, 32'sd0.08320272840026563, 32'sd0.08691329341595323, 32'sd0.14093809377906025, 32'sd-0.005647551367814473, 32'sd-0.06022254084899439, 32'sd0.01687121093850721, 32'sd0.0013029197409574324, 32'sd-0.08013787782134758, 32'sd0.019513074117835847, 32'sd0.06659359108147288, 32'sd-0.02592655223659149, 32'sd0.007630694309191869, 32'sd-0.0063522092962136146, 32'sd-7.594526078912348e-124, 32'sd-5.1172280137462e-127, 32'sd0.04076071524630105, 32'sd-0.07900165262767751, 32'sd0.0017307124844933616, 32'sd-0.09008950313575945, 32'sd-0.03719237895178475, 32'sd0.02300286778711069, 32'sd0.0511372801441904, 32'sd0.059002244121504524, 32'sd0.007047918741351944, 32'sd-0.0861967725832561, 32'sd0.02034025912673724, 32'sd0.05493382877537751, 32'sd0.15173961171489248, 32'sd0.10099860193159235, 32'sd0.17218926514677818, 32'sd0.06818733267600141, 32'sd0.004348576912334254, 32'sd-0.0696019767369623, 32'sd0.09137906905666378, 32'sd0.11115597793554931, 32'sd-0.0025559914530394992, 32'sd0.039403996898304434, 32'sd0.080712598605916, 32'sd-0.0035785667336038153, 32'sd0.05009061810207615, 32'sd0.06028711023720025, 32'sd-0.03911688710375345, 32'sd2.4464753038594175e-121, 32'sd0.037117515062904574, 32'sd0.04976430569430227, 32'sd-0.1045055660391159, 32'sd0.014356093147273919, 32'sd-0.04330990611114722, 32'sd-0.055505839827067194, 32'sd-0.07913775874037085, 32'sd-0.034261530833971834, 32'sd-0.012935233085006303, 32'sd-0.06333290016009184, 32'sd0.16972332913492758, 32'sd0.11289072403881412, 32'sd0.03590112874531271, 32'sd0.013440332344949322, 32'sd0.046955621250501185, 32'sd0.08371819603326372, 32'sd0.02908495652704854, 32'sd0.039779010630040364, 32'sd0.0670710346276962, 32'sd0.01996692641040569, 32'sd-0.0030109065936772847, 32'sd-0.047109197748608354, 32'sd0.05137987032848997, 32'sd-0.031468972649170056, 32'sd-0.05932951433555823, 32'sd0.06869220191974072, 32'sd0.09268386034251253, 32'sd-2.8522318648447412e-129, 32'sd0.07806360253089967, 32'sd-0.004407956614522393, 32'sd0.06429060878731999, 32'sd0.04101217493189997, 32'sd-0.06662469906603138, 32'sd0.03158508442076809, 32'sd-0.08193798414719596, 32'sd-0.028480158285876533, 32'sd0.15206061620938713, 32'sd-0.022852920116525493, 32'sd0.043221407436337726, 32'sd-0.0028613602282526332, 32'sd0.07978983942436421, 32'sd0.0032177899669541773, 32'sd-0.004693340741405857, 32'sd0.07095183303054559, 32'sd0.028643540573076387, 32'sd0.06848689149792224, 32'sd-0.0663570396990781, 32'sd-0.1498810135861009, 32'sd0.008772092598881651, 32'sd-0.10160158270140132, 32'sd0.008273034593539806, 32'sd0.09336860730024558, 32'sd0.0780460843196497, 32'sd0.06787926975084202, 32'sd0.006147238718012805, 32'sd0.015259774183944313, 32'sd-0.022565622111118264, 32'sd0.054868824420264146, 32'sd-0.032381716719837465, 32'sd0.06571521050557953, 32'sd0.008540770915103267, 32'sd0.021009230823087664, 32'sd-0.031044997504518945, 32'sd0.028913974114844258, 32'sd0.03347181106223635, 32'sd0.0491325365048943, 32'sd0.25759498138286774, 32'sd0.09758390845189399, 32'sd0.07955491162295313, 32'sd-0.003139778076468519, 32'sd0.08743116129739995, 32'sd0.10260866296742564, 32'sd-0.004261532084247997, 32'sd0.008431411742941028, 32'sd-0.0007148847824134085, 32'sd-0.027607351113318607, 32'sd-0.04729804621958266, 32'sd-0.04475557297972316, 32'sd-0.07633015909855198, 32'sd0.04237011143085494, 32'sd0.1278411871393412, 32'sd-0.04521840261613839, 32'sd-0.047599006807166645, 32'sd0.03214319068705765, 32'sd0.03823422648535828, 32'sd-0.11077414943622349, 32'sd-0.0420258895844223, 32'sd-0.0026101687046366923, 32'sd-0.0314646214358136, 32'sd-0.04751402530278033, 32'sd0.07680700107038099, 32'sd0.221455195817558, 32'sd0.07308912718404785, 32'sd0.008962173244367419, 32'sd0.09266531488930657, 32'sd0.01910014950019964, 32'sd0.01131599906688935, 32'sd-0.036228091059051136, 32'sd-0.13008430655232672, 32'sd-0.16823460936939016, 32'sd-0.12105796548316543, 32'sd-0.0736016883739348, 32'sd0.03338909427129972, 32'sd-0.030247544576388764, 32'sd0.005081979040848314, 32'sd-0.06418952110894355, 32'sd-0.0011208424577225846, 32'sd-0.09294973734038722, 32'sd0.07283285210093374, 32'sd0.053603179370595964, 32'sd0.05166310347119388, 32'sd-0.052785991850326654, 32'sd-0.0377665485102192, 32'sd0.006546659646323582, 32'sd-0.07505535341286912, 32'sd0.00713165838084698, 32'sd0.09056884459801445, 32'sd0.06032047396813847, 32'sd0.06160448087114202, 32'sd0.12442910343894076, 32'sd0.09817336807666384, 32'sd0.03637549700532295, 32'sd0.0338999244700925, 32'sd0.006965950030936743, 32'sd-0.027522847522080014, 32'sd-0.0779722773232355, 32'sd-0.011420791438177622, 32'sd-0.02611000837147941, 32'sd-0.08311435783419324, 32'sd-0.03687759881859852, 32'sd-0.07651037914263875, 32'sd-0.06140357297680889, 32'sd-0.03613790323699389, 32'sd0.04380180051414473, 32'sd-0.023137554981100785, 32'sd-0.12284251690837501, 32'sd-0.07984652674081696, 32'sd0.020244570947571643, 32'sd-0.08972337382144445, 32'sd0.0068571860495756495, 32'sd-0.1370906131341425, 32'sd-0.029393906004238073, 32'sd0.06434576971712687, 32'sd0.08277767815425045, 32'sd0.017718400599682403, 32'sd0.05034073437783459, 32'sd0.010807770714683097, 32'sd-0.12383463847726453, 32'sd-0.005912719433188222, 32'sd0.048080533913933715, 32'sd-0.07436003359366739, 32'sd0.04650358015910282, 32'sd0.056676955538674696, 32'sd0.06386074298277705, 32'sd-0.016874826030107128, 32'sd0.05920550117419924, 32'sd0.021349402258017135, 32'sd-0.03875117630919607, 32'sd0.02772555600062444, 32'sd-0.08345943173253934, 32'sd-0.06746693861337227, 32'sd-0.056035068078309706, 32'sd-0.060261906277657776, 32'sd0.050031545880760704, 32'sd0.004203129822981597, 32'sd-0.04374006166777731, 32'sd0.05635307186641696, 32'sd-0.023512716470782045, 32'sd0.040129992299737446, 32'sd-0.009437112497169055, 32'sd0.020490618325590612, 32'sd0.02849401461471376, 32'sd0.011607793769222113, 32'sd0.004114674491420226, 32'sd-0.016495269049398905, 32'sd-0.14930754100889107, 32'sd-0.18637816064537485, 32'sd0.08186547872900214, 32'sd0.13280583523705827, 32'sd0.08220260776382207, 32'sd0.07508651706295089, 32'sd0.11389626401235778, 32'sd-0.002611022535875481, 32'sd0.1268696949924514, 32'sd-0.01424068474191001, 32'sd-0.10036102214420974, 32'sd-0.127749493597833, 32'sd-0.1696394662913736, 32'sd-0.06752556436019803, 32'sd-0.09298291264510423, 32'sd-0.048962286393900725, 32'sd-0.010379381562142676, 32'sd-0.026559608581983883, 32'sd-0.03715188930073431, 32'sd0.10235344172612139, 32'sd0.03914677191373905, 32'sd-0.07217677290684239, 32'sd-0.019989768986069013, 32'sd-0.05775021660914916, 32'sd0.06259841160885346, 32'sd-0.029289566117404044, 32'sd-0.13996460424255908, 32'sd-0.07418986749401889, 32'sd-0.06354850487951201, 32'sd-0.02058054447291199, 32'sd0.024064251922045272, 32'sd-0.017964645430388487, 32'sd0.034093598373231435, 32'sd0.06336105585477331, 32'sd0.04276024862215511, 32'sd0.02311174132835116, 32'sd-0.00503442887434822, 32'sd0.01436242937804574, 32'sd-0.01014222164980825, 32'sd-0.01073114363339604, 32'sd0.09782844597613982, 32'sd0.06796643727590021, 32'sd-0.08052531287055498, 32'sd-0.01604685068298843, 32'sd-0.059663976101803906, 32'sd-0.03682123243164616, 32'sd-0.047732006354765544, 32'sd0.0001361005391331325, 32'sd0.039187069232700295, 32'sd0.05180724930018722, 32'sd-0.00538037598746715, 32'sd-0.021200492026036726, 32'sd0.00024176618611579883, 32'sd0.04216845631434299, 32'sd-0.1355920443493365, 32'sd-0.07923656249102294, 32'sd-0.13759446333062753, 32'sd-0.0604803472085062, 32'sd-0.06785427683515387, 32'sd0.014161154583099463, 32'sd0.02834696391801157, 32'sd-0.01140980706017449, 32'sd-0.05349865598573467, 32'sd-0.1990089547531047, 32'sd-0.08307959313703737, 32'sd0.012302325508260378, 32'sd0.08987513228072398, 32'sd0.11796723342370831, 32'sd0.15493401522715794, 32'sd0.18579295100617788, 32'sd-0.036562433075696336, 32'sd0.026572908544937743, 32'sd0.04718903694429079, 32'sd0.03965044134003205, 32'sd-0.03116211037341192, 32'sd0.06833495830007236, 32'sd0.06437560996383544, 32'sd-0.022873214181880347, 32'sd-0.07966101067447715, 32'sd0.05944636316666386, 32'sd-0.2033381656013416, 32'sd-0.08780701877928308, 32'sd-0.12368255659014551, 32'sd-0.055050848491805665, 32'sd-0.21272524494824005, 32'sd-0.17450912468043958, 32'sd-0.2738414662483489, 32'sd-0.14777915551419582, 32'sd-0.062064979143297436, 32'sd0.009117603862501659, 32'sd0.023589713774479135, 32'sd-0.044574126210707596, 32'sd0.046523146441660584, 32'sd-0.11887977608209062, 32'sd0.06755800349900065, 32'sd-0.006221550759134686, 32'sd0.0781824708385698, 32'sd0.03479942797520199, 32'sd0.01430205994926187, 32'sd0.03022243631249387, 32'sd-0.1030468391751575, 32'sd-0.026045768921469075, 32'sd-0.027614116566978302, 32'sd0.11101293483978458, 32'sd0.10470830565366762, 32'sd0.06647553629335051, 32'sd0.10341879653920814, 32'sd-0.0327680052858909, 32'sd-0.2046205193460202, 32'sd-0.17239372124513053, 32'sd-0.20356537524487792, 32'sd-0.17906147859445112, 32'sd-0.22084747182872735, 32'sd-0.34893154345384225, 32'sd-0.22624239689294146, 32'sd-0.2154026660063228, 32'sd-0.0807250599025776, 32'sd-0.05430864144146091, 32'sd0.1511086008098315, 32'sd0.11902376836051189, 32'sd0.07264481838425337, 32'sd0.03657930685272959, 32'sd-0.05959566397272405, 32'sd0.050269468047384136, 32'sd0.039417108576784585, 32'sd0.016132369568937356, 32'sd0.018864764960223226, 32'sd0.04084003846075713, 32'sd-0.070166142675649, 32'sd-0.032537531815761044, 32'sd-0.015268294138319292, 32'sd0.04150646688520955, 32'sd0.036615757058114595, 32'sd-0.07485374732946458, 32'sd0.02809456766167354, 32'sd0.04933985230130189, 32'sd-0.11317532182470082, 32'sd-0.0846349591116487, 32'sd-0.21333861021930528, 32'sd-0.24423175869779054, 32'sd-0.36260616945472685, 32'sd-0.2957239750159591, 32'sd-0.20495031925100285, 32'sd-0.3208682839689979, 32'sd-0.13735677144632014, 32'sd0.018826862905737693, 32'sd0.12229246485818328, 32'sd0.11754929076882949, 32'sd0.01521682655409186, 32'sd0.07381727391860629, 32'sd-0.031117918846992415, 32'sd0.048714676211070826, 32'sd0.007990242158172607, 32'sd0.06903405370860945, 32'sd0.09889993001472837, 32'sd-0.020912805566750223, 32'sd-0.05932228842596895, 32'sd0.10455129312494912, 32'sd0.04913808832694487, 32'sd-0.03474707058278969, 32'sd2.94087802148018e-125, 32'sd0.04452549246293342, 32'sd-0.047797891946003444, 32'sd-0.04343689741245498, 32'sd-0.15591808234007268, 32'sd-0.012058102461470245, 32'sd-0.16109927567308965, 32'sd-0.19071704616203722, 32'sd-0.11677545128265238, 32'sd-0.2510500494112236, 32'sd-0.24352910822909193, 32'sd-0.24846747800367114, 32'sd-0.2696956791523027, 32'sd-0.007683636955012435, 32'sd0.03243691431628684, 32'sd0.042310061484663736, 32'sd-0.11411953739048451, 32'sd0.00888941676510773, 32'sd0.031115579258776206, 32'sd-0.07320291132599457, 32'sd0.019767026262901603, 32'sd0.0566096746146036, 32'sd-0.07274015492284318, 32'sd-0.09508544580293843, 32'sd-0.0418374679584905, 32'sd0.14723424419550754, 32'sd0.07514493589052623, 32'sd0.05469012089505737, 32'sd-0.010356246069068844, 32'sd0.07112504263285956, 32'sd0.08663433631266691, 32'sd0.08882499757043091, 32'sd-0.0033708082488619912, 32'sd-0.010298535001717844, 32'sd-0.06976690631561612, 32'sd-0.12688579133952496, 32'sd-0.08265070664231897, 32'sd-0.12229347892501449, 32'sd-0.10690984741537363, 32'sd-0.13895967007819818, 32'sd-0.2110860908265047, 32'sd-0.03023729999332797, 32'sd-0.06034890150365711, 32'sd0.025021183023191236, 32'sd0.08594558311181713, 32'sd0.027789935228072233, 32'sd-0.03127647944836111, 32'sd0.015059337385821842, 32'sd-0.05997757310140685, 32'sd0.03863199298681399, 32'sd-0.018698714624668766, 32'sd0.044774392675534916, 32'sd-0.07808302477490352, 32'sd0.02689552165989919, 32'sd-5.6180092272353116e-05, 32'sd-0.045675105663574384, 32'sd0.0260424163663931, 32'sd-0.020335515331796207, 32'sd0.006096307212507621, 32'sd0.07559776461029094, 32'sd-0.0075614813066243475, 32'sd-0.0012945656011408356, 32'sd0.04806240526733662, 32'sd-0.013659469140698415, 32'sd0.017356133145431725, 32'sd-0.05889217374391746, 32'sd0.14132812801973998, 32'sd0.05334929703677297, 32'sd-0.08534948042916668, 32'sd-0.007614528330352364, 32'sd-0.06826988539069735, 32'sd-0.05353631840330304, 32'sd0.14399284003837318, 32'sd0.05500917780265465, 32'sd-0.05918780580760055, 32'sd-0.016200190925381906, 32'sd-0.030620755630310192, 32'sd-0.1229645761100829, 32'sd0.01098193084635888, 32'sd0.04351325048221535, 32'sd-0.04924052980541345, 32'sd-0.032675119636982226, 32'sd0.09155879343950457, 32'sd0.01660198276186365, 32'sd-6.1087935574188635e-124, 32'sd0.048920193389630336, 32'sd0.03464614232748958, 32'sd-0.0810714285680619, 32'sd0.0136331767924716, 32'sd0.04794344149960297, 32'sd0.12545961121514598, 32'sd0.047849049602433635, 32'sd0.14787529117875822, 32'sd0.0936969448552681, 32'sd0.20392690723390894, 32'sd0.19030143342872624, 32'sd0.18342440268457932, 32'sd0.1431656409709795, 32'sd-0.05521610872590768, 32'sd-0.01663730894986078, 32'sd0.16482260077380528, 32'sd0.03283414484007208, 32'sd0.00469599005621428, 32'sd-0.02480572548066717, 32'sd-0.0503008605197248, 32'sd0.026730533854401047, 32'sd0.05614937644043957, 32'sd-0.07604228391065453, 32'sd0.02865645119566393, 32'sd0.00905245513732802, 32'sd0.10579241067118164, 32'sd-0.03015696034402488, 32'sd0.09887013345017306, 32'sd-0.0077128017633491565, 32'sd0.04902032176571394, 32'sd-0.054658762693800995, 32'sd0.060241783823272874, 32'sd0.08635975926097404, 32'sd0.04856851014705233, 32'sd0.08525748236099345, 32'sd0.10720061042912372, 32'sd0.18839664818308657, 32'sd0.2688314735325629, 32'sd0.2549455833094254, 32'sd0.2318594315021431, 32'sd0.23246285748431159, 32'sd-0.007798058673438133, 32'sd-0.005939088531350739, 32'sd0.09805466938590343, 32'sd0.14664601645509068, 32'sd0.1388447000755711, 32'sd0.02323994545547362, 32'sd0.15617268876311705, 32'sd0.06503677983483297, 32'sd-0.05157789988810686, 32'sd0.09326146802836116, 32'sd0.13248520351600646, 32'sd-0.014654229260172083, 32'sd-0.02939268360183129, 32'sd0.030611865023497335, 32'sd0.05206185839792443, 32'sd0.03986234494697037, 32'sd-0.009208480871392737, 32'sd0.09094299441524774, 32'sd0.0631412449790258, 32'sd-0.08087673297024371, 32'sd0.03502900073167775, 32'sd0.13309001423776542, 32'sd0.12939243236937104, 32'sd0.11544680766597179, 32'sd0.1296358589860374, 32'sd0.09087569456565021, 32'sd0.12633752141573715, 32'sd0.1603187169551588, 32'sd0.15668298011110046, 32'sd0.1818268291293327, 32'sd0.09648279214278552, 32'sd0.045997749251074915, 32'sd0.11764917711398722, 32'sd-0.04181630532133785, 32'sd0.09634557984439106, 32'sd0.041312715007625865, 32'sd0.07279041887328981, 32'sd0.19852822688310795, 32'sd0.014953247963904157, 32'sd0.11565611531364524, 32'sd0.03172350446537159, 32'sd0.055301547928115986, 32'sd1.5541421663218633e-123, 32'sd0.079140120928213, 32'sd0.10630112839363975, 32'sd0.04739719284344979, 32'sd-0.016542984885578572, 32'sd-0.059377550793437234, 32'sd0.02892504962482459, 32'sd-0.019916664045370232, 32'sd0.15229905085382553, 32'sd0.11242840054459942, 32'sd0.11780996056180162, 32'sd0.1799524321674088, 32'sd0.13367487982665308, 32'sd0.15504114646475625, 32'sd0.1377951669044043, 32'sd0.15335420210738068, 32'sd0.13684413424274638, 32'sd-0.038416414528660174, 32'sd-0.03131176946611865, 32'sd0.05715156299510823, 32'sd-0.016937022004652746, 32'sd0.1051824981067755, 32'sd0.0817913898716215, 32'sd0.03671241819876544, 32'sd-0.03048986705127529, 32'sd-0.07944657408883922, 32'sd-0.03565491884332993, 32'sd7.885815416727625e-124, 32'sd-1.6931088420788894e-127, 32'sd2.9526915995469055e-120, 32'sd-0.025926208102561455, 32'sd-0.13534231227875865, 32'sd-0.14967173192717087, 32'sd-0.0007596983997393582, 32'sd0.09258027308679148, 32'sd0.07234775237938212, 32'sd-0.042125792823074916, 32'sd-0.07923895892334103, 32'sd-0.03657408650042241, 32'sd0.022611323011647227, 32'sd-0.03303772883348611, 32'sd-0.03129971710368749, 32'sd0.13932826334274, 32'sd-0.06590476131889593, 32'sd0.05307284968317279, 32'sd0.02389099567416532, 32'sd0.1137341719108599, 32'sd0.11845434956213734, 32'sd-0.02742689456787213, 32'sd0.055023937052918595, 32'sd0.00430296248606877, 32'sd0.04604188439163694, 32'sd0.05666486845899605, 32'sd-0.025547817835485327, 32'sd0.015925849584907312, 32'sd-5.066599297713245e-125, 32'sd7.240461017623326e-117, 32'sd1.789238068004187e-121, 32'sd-0.0008827078966026107, 32'sd0.06785782762918935, 32'sd-0.10776271529075752, 32'sd-0.10739938211481347, 32'sd0.06139818193073564, 32'sd-0.030857254427082283, 32'sd-0.058321489316591826, 32'sd-0.08153941509489385, 32'sd-0.047943799115606985, 32'sd0.021178707462142243, 32'sd0.07291799989365924, 32'sd0.11853902895522485, 32'sd0.14061744766774378, 32'sd0.04929182658224123, 32'sd-0.03293566914652963, 32'sd0.05631204904303766, 32'sd-0.0666231882782998, 32'sd0.014901242250146414, 32'sd0.009180976738801685, 32'sd-0.09526237831303833, 32'sd-0.09233048382052983, 32'sd-0.0802204363097709, 32'sd0.04659330122582516, 32'sd-0.001996789165446223, 32'sd0.07621109392847908, 32'sd-1.8348957521591966e-117, 32'sd-2.614566352386443e-119, 32'sd6.032585568879411e-115, 32'sd1.1021266208274721e-119, 32'sd0.0792731392251807, 32'sd0.029288573980595665, 32'sd-0.028039550162674644, 32'sd-0.02817346027633221, 32'sd0.06299029670777116, 32'sd0.056456364200761146, 32'sd-0.052178486327442306, 32'sd-0.04634115467742227, 32'sd0.05926990731005707, 32'sd-0.019258552455709663, 32'sd0.011924561481816446, 32'sd-0.08728706208201138, 32'sd-0.09893106971443412, 32'sd-0.05274027477513178, 32'sd0.019704686262072023, 32'sd-0.021445039745192403, 32'sd-0.09561356404723523, 32'sd-0.03599422342210741, 32'sd-0.0012039254687711497, 32'sd0.04587954599843492, 32'sd-0.011902468052421131, 32'sd0.0367017223323357, 32'sd-0.03390511259242446, 32'sd3.5164613496001497e-115, 32'sd-2.2704295036987318e-126, 32'sd-2.9069674400280614e-120, 32'sd-7.529238960072882e-115, 32'sd1.5352743816323588e-123, 32'sd3.39089099234941e-114, 32'sd0.013036659197471757, 32'sd0.043650745503186685, 32'sd0.00010404485763539762, 32'sd0.0741506496806668, 32'sd0.09265674907935492, 32'sd0.08529045495798357, 32'sd-0.020507707551870247, 32'sd-0.009810137969182215, 32'sd0.057558181925192006, 32'sd-0.03150694905223872, 32'sd0.061346547404174265, 32'sd-0.03207034628764497, 32'sd0.07642066340314395, 32'sd0.006242263516086151, 32'sd0.014588816803091993, 32'sd0.03329169035965678, 32'sd-0.05423069730458297, 32'sd0.01516831711449067, 32'sd-0.012246907573983404, 32'sd0.032077712800868484, 32'sd-7.560293869257927e-115, 32'sd8.731455091118764e-126, 32'sd-1.7737074648971658e-123, 32'sd-1.0977121011523024e-117},
        '{32'sd1.7306085827309038e-125, 32'sd1.4838386639216176e-115, 32'sd-6.051485448664465e-125, 32'sd-1.5964820172596355e-115, 32'sd2.593885736960388e-126, 32'sd-1.0175003846393201e-126, 32'sd2.6018699324143223e-124, 32'sd2.1420427527595954e-124, 32'sd1.5858207004047734e-115, 32'sd1.1757050319653796e-127, 32'sd1.9206724187186552e-127, 32'sd1.5952547507602145e-124, 32'sd-0.0015866801358493312, 32'sd-0.06761513431331757, 32'sd-0.04305936821945786, 32'sd0.02437402282311584, 32'sd-8.429949597886047e-121, 32'sd-2.5904219987288354e-115, 32'sd-1.391431505532871e-125, 32'sd7.295180388867555e-128, 32'sd-1.0878724767761663e-121, 32'sd1.1261677850600817e-119, 32'sd-6.59328157252185e-123, 32'sd-2.6169344931941395e-126, 32'sd-5.070641101565789e-120, 32'sd-9.063857655828833e-126, 32'sd-6.648392148755906e-117, 32'sd-9.364357549529916e-123, 32'sd9.613664733031365e-115, 32'sd3.662070495484468e-116, 32'sd-6.170694102014112e-119, 32'sd3.3123634477296496e-117, 32'sd0.0008137167276948383, 32'sd0.0031219336301476896, 32'sd0.010728052543404094, 32'sd-0.050587306295848324, 32'sd-0.041116773901489385, 32'sd-0.05240348604315397, 32'sd-0.09103216641611964, 32'sd-0.09423660767591377, 32'sd-0.08722630219009037, 32'sd-0.01605359742812377, 32'sd0.017286029815645455, 32'sd-0.007316781881856364, 32'sd0.014617686913038167, 32'sd-0.1047960778562697, 32'sd0.03776206702318817, 32'sd-0.06981671359747131, 32'sd0.03410522306015194, 32'sd0.06862839638991726, 32'sd-0.024959999318111162, 32'sd-0.06632028505285611, 32'sd-5.270896928691387e-116, 32'sd-3.633964606540965e-122, 32'sd-9.585567229458736e-125, 32'sd2.9609111420155894e-125, 32'sd-1.1036818033978683e-121, 32'sd-5.950344772548353e-126, 32'sd0.0026730281958323616, 32'sd-0.004992831351291879, 32'sd-0.0892306879015412, 32'sd-0.04832480237154688, 32'sd-0.022961011220293485, 32'sd-0.06802251784020048, 32'sd-0.04717980079825192, 32'sd0.029209183124617476, 32'sd0.04166344176304928, 32'sd0.01340105825469727, 32'sd0.12479218275593879, 32'sd-0.07626868037874819, 32'sd-0.033418341425172665, 32'sd0.02258824581096013, 32'sd-0.10590600689497912, 32'sd0.020780527016909935, 32'sd-0.01572362533570961, 32'sd-0.015305298056387322, 32'sd-0.047648844686743075, 32'sd0.0747327529062266, 32'sd0.06557261888564599, 32'sd-0.08914339994711239, 32'sd-0.009770905802446744, 32'sd-0.07310868583480842, 32'sd3.6777156320850704e-116, 32'sd-5.376922139148805e-118, 32'sd8.318126455374282e-121, 32'sd2.3450148418660716e-116, 32'sd0.013483232092307385, 32'sd-0.05370154053646526, 32'sd-0.08390798898930817, 32'sd-0.0782673071691814, 32'sd-0.10728818472825916, 32'sd-0.13943869814965998, 32'sd-0.045406365780838245, 32'sd0.004354839494627252, 32'sd0.026092829553057396, 32'sd0.0249609446233979, 32'sd-0.01503760826918531, 32'sd0.0534683956351805, 32'sd0.1336078838556053, 32'sd0.04245033075109304, 32'sd0.028482453793545356, 32'sd-0.05862106227527355, 32'sd-0.005791210724329413, 32'sd-0.0019740043040747273, 32'sd-0.07356332611941982, 32'sd0.11994405479388356, 32'sd-0.045731938463332594, 32'sd0.013201947693704573, 32'sd0.048558361711830415, 32'sd0.005465641799319566, 32'sd-0.01911946206574159, 32'sd-1.2940327900218089e-120, 32'sd5.113442717021331e-123, 32'sd0.01620819888444104, 32'sd-0.07749869034686209, 32'sd-0.007456623501760617, 32'sd-0.10988644964599344, 32'sd-0.018661590103516177, 32'sd-0.017701168478346723, 32'sd0.037157073706398765, 32'sd-0.0189351522110435, 32'sd0.1327365589940892, 32'sd0.019936998087024226, 32'sd-0.027707106237440163, 32'sd-0.08480414526852903, 32'sd0.04932891269573041, 32'sd0.01959023112795787, 32'sd0.08170807708897647, 32'sd0.0483298975827548, 32'sd0.13617156221727897, 32'sd0.05105455689339709, 32'sd-0.027410171340524522, 32'sd0.07940092380039769, 32'sd0.1089524225276802, 32'sd0.09460301437376942, 32'sd-0.025219441047845164, 32'sd0.09617700098697582, 32'sd-0.030774768072919005, 32'sd-0.0003353333716972471, 32'sd0.020473670016520916, 32'sd-3.24835429930648e-123, 32'sd0.03336942057232815, 32'sd-0.016762591990978414, 32'sd-0.018316407318363277, 32'sd-0.08552781654786537, 32'sd-0.04811867494925131, 32'sd0.09037503948191304, 32'sd-0.016328700304020047, 32'sd-0.027580388859232186, 32'sd-0.04190801145632618, 32'sd-0.06548246672308317, 32'sd-0.05662578709469888, 32'sd0.09250459196502064, 32'sd0.15769149329683296, 32'sd0.08040005793798838, 32'sd0.08229683525337148, 32'sd0.09250984785695525, 32'sd0.10002064944323089, 32'sd0.016837062248352585, 32'sd0.09715436435128504, 32'sd0.16129904106633292, 32'sd0.11201220969024722, 32'sd0.027947026571700354, 32'sd0.01139418629931842, 32'sd0.03564158919318981, 32'sd0.007572082903468056, 32'sd0.01292586392999006, 32'sd0.012798975452500036, 32'sd-4.0858431915988045e-125, 32'sd0.02327271767503844, 32'sd0.07369259844581928, 32'sd-0.052746489724016875, 32'sd-0.06553458034642456, 32'sd0.018459034322020586, 32'sd0.010483178910585466, 32'sd-0.08009067664326196, 32'sd0.00962622230167377, 32'sd-0.009180241238722289, 32'sd-0.015493618980183426, 32'sd0.0374882736079716, 32'sd0.0701941449180616, 32'sd0.03172889028635997, 32'sd0.0474576493539745, 32'sd-0.13043185712411096, 32'sd-0.024984595744105456, 32'sd0.0498677486365355, 32'sd-0.0072032871062039545, 32'sd0.09788511117957796, 32'sd-0.028273798818048146, 32'sd-0.007827252397929961, 32'sd0.14017334749338642, 32'sd-0.0149261485539201, 32'sd0.027785804908068427, 32'sd0.06084844860407725, 32'sd0.031151746956465567, 32'sd-0.00043772150926972705, 32'sd0.01466986945005114, 32'sd0.023908828224641958, 32'sd0.07752450352463429, 32'sd0.09278393729183425, 32'sd0.0258393924600045, 32'sd-0.10531754064348006, 32'sd-0.0025811155040092386, 32'sd0.04436410065875756, 32'sd-0.020716841737778713, 32'sd0.07966610395554986, 32'sd0.051376546629429386, 32'sd-0.06620960713527269, 32'sd0.06724213796484572, 32'sd0.056154931581165676, 32'sd-0.10772577887697904, 32'sd0.011834511440263864, 32'sd-0.12453802459889264, 32'sd-0.05460499895402863, 32'sd0.10747153513433431, 32'sd-0.0989713134078939, 32'sd-0.033495475088384324, 32'sd-0.05157640509873393, 32'sd-0.03803661074560778, 32'sd0.04270156384814578, 32'sd0.033969676987117205, 32'sd0.07582130393895731, 32'sd-0.02684388032738472, 32'sd0.058083360610134235, 32'sd0.0055311014578497564, 32'sd0.04516755298344031, 32'sd-0.028436174301077838, 32'sd-0.0666013564782998, 32'sd0.05209015680862235, 32'sd-0.03813245972332941, 32'sd0.04521028706294515, 32'sd-0.04232601471020703, 32'sd-0.07298883647403168, 32'sd0.03968788344927288, 32'sd0.004092845351108662, 32'sd-0.05371365880376011, 32'sd-0.026015953099829545, 32'sd0.09570879818222576, 32'sd-0.006508379992653506, 32'sd-0.08645442092850156, 32'sd-0.08057471796332216, 32'sd-0.0879094281065373, 32'sd0.0978519235074823, 32'sd0.05723493233313174, 32'sd0.00977886167459471, 32'sd0.03360316557986199, 32'sd0.013405236915213, 32'sd0.042218626478726894, 32'sd-0.04517664960340171, 32'sd0.027221766996220025, 32'sd0.036102252601855504, 32'sd0.016590230549285653, 32'sd-0.06073006996728456, 32'sd-0.07786025113292228, 32'sd-0.12346851742721734, 32'sd-0.03096498248227405, 32'sd0.08923680118449545, 32'sd0.06067210573095893, 32'sd-0.04190472254366608, 32'sd-0.03267831595658, 32'sd-0.011416915666008375, 32'sd0.0011534136716421094, 32'sd-0.1017878482244873, 32'sd-0.039805394799528215, 32'sd-0.039182771309789255, 32'sd0.04199673473824253, 32'sd-0.023272531212667494, 32'sd-0.14045500790380205, 32'sd-0.2466073950770088, 32'sd-0.059626229236904124, 32'sd0.06781803007485271, 32'sd0.1512740805815109, 32'sd0.09175325632204356, 32'sd0.10991682566297813, 32'sd0.09759694182314237, 32'sd0.1250919226410858, 32'sd-0.020668155042831628, 32'sd0.06431674305185825, 32'sd0.04281229177779298, 32'sd0.045756788734952605, 32'sd-0.08147920600435246, 32'sd-0.04648827777473257, 32'sd0.005146959258780318, 32'sd0.11556841773866616, 32'sd-0.07420473962377923, 32'sd0.0038961837693015536, 32'sd0.06048765609800823, 32'sd0.006548689060073952, 32'sd0.057628463208841664, 32'sd-0.07301747084582932, 32'sd-0.10942938539366007, 32'sd-0.10575081803208165, 32'sd-0.07361641257950455, 32'sd0.038910579671340755, 32'sd0.22952783549228006, 32'sd0.024190090783697514, 32'sd-0.0666218040109105, 32'sd-0.13221447802090988, 32'sd0.08211837674390687, 32'sd0.043710398825260614, 32'sd0.17150526213119396, 32'sd0.18046107715608353, 32'sd0.09552463253954818, 32'sd0.06307408053111899, 32'sd-0.2059145793765005, 32'sd-0.1597723466104224, 32'sd-0.047076885695463526, 32'sd0.025532458145038964, 32'sd-0.04303324320350804, 32'sd-0.004605994581905949, 32'sd0.09998294976024417, 32'sd0.0162089042037783, 32'sd-0.0704942843599223, 32'sd-0.026343308957968135, 32'sd0.05698253550013611, 32'sd0.08151043340856691, 32'sd-0.0011657974666842768, 32'sd-0.16847710650496447, 32'sd-0.07099122358812691, 32'sd-0.19698322149645403, 32'sd0.040595530407300184, 32'sd0.12221706149764279, 32'sd0.2530171251854844, 32'sd0.1797409225163586, 32'sd-0.010142884070166468, 32'sd-0.003236264943433327, 32'sd0.08571519979631591, 32'sd0.1829415015132049, 32'sd0.15874225851743162, 32'sd0.052027311170033286, 32'sd0.10744483090273986, 32'sd0.012497046347855648, 32'sd-0.11180118260499641, 32'sd-0.04724390153946801, 32'sd0.008420541380954586, 32'sd0.0030044671010888042, 32'sd0.04889011521283729, 32'sd0.08162200398582778, 32'sd0.03530717959833099, 32'sd-0.018326767117812857, 32'sd-0.07551768981826279, 32'sd0.07019825466819803, 32'sd0.0040694314326236445, 32'sd-0.13900986001917887, 32'sd-0.1730601408542573, 32'sd-0.18828533956508203, 32'sd-0.15058254950468164, 32'sd-0.004287602876592843, 32'sd0.07661207472477302, 32'sd0.17307680521026553, 32'sd0.2918781495351751, 32'sd0.2460998596911154, 32'sd0.06526324389365429, 32'sd0.1428257519807394, 32'sd0.05090537865645746, 32'sd0.07755387483259676, 32'sd-0.0186357583630194, 32'sd-0.026170266616315968, 32'sd-0.03535413166198512, 32'sd-0.1433231747512815, 32'sd-0.0413386334310755, 32'sd-0.08143226707252511, 32'sd-0.0011026057615437334, 32'sd-0.07615729609965993, 32'sd-0.06356131328090332, 32'sd0.045876315636481625, 32'sd0.03983593722551087, 32'sd-0.0715649131313613, 32'sd-0.12341039615117591, 32'sd-0.09219584337500303, 32'sd-0.10831653518256328, 32'sd-0.10534744996108518, 32'sd-0.029289621928726077, 32'sd-0.13358305404306486, 32'sd0.01687196433658129, 32'sd0.2212927196002224, 32'sd0.2408467607728732, 32'sd0.19451953144561684, 32'sd0.23689977695144182, 32'sd0.1056826157921672, 32'sd0.06234408007892151, 32'sd0.0766998344472911, 32'sd0.021938171863115474, 32'sd-0.10084453921809974, 32'sd-0.12417366204853002, 32'sd-0.08043407735085092, 32'sd-0.06520805788597658, 32'sd-0.16590007039806096, 32'sd-0.14774943109878702, 32'sd-0.010623752366363667, 32'sd0.044766739258148135, 32'sd0.05000476987781062, 32'sd-0.02494490796492122, 32'sd-0.054475235167129335, 32'sd-0.12113437995026106, 32'sd-0.013916616028734757, 32'sd-0.0448252525366729, 32'sd0.09003927838799126, 32'sd-0.14190482787380934, 32'sd-0.14443779635898676, 32'sd-0.14332220686870809, 32'sd-0.06918461563139759, 32'sd0.08150548931871307, 32'sd0.08949056446149371, 32'sd0.03313819019231912, 32'sd-0.00760170808363251, 32'sd0.08745247563432769, 32'sd0.058139098483259925, 32'sd0.15955128574768446, 32'sd0.1630516602531792, 32'sd-0.06400945014159562, 32'sd-0.166822903479702, 32'sd0.013669233478065024, 32'sd0.005570164783636624, 32'sd-0.02536235798520942, 32'sd-0.08759988351347119, 32'sd-0.0756128870753358, 32'sd-0.048803441138677475, 32'sd-0.11147314392221931, 32'sd-0.04950749375868496, 32'sd-0.07464931914814242, 32'sd-0.01438101277517809, 32'sd0.0035518579624177933, 32'sd-0.03596635229588577, 32'sd0.030631505342255394, 32'sd0.006693114620975648, 32'sd-0.011422376602919681, 32'sd-0.08033589198806831, 32'sd-0.03210110748999156, 32'sd0.10608111566190935, 32'sd-0.0325446212089767, 32'sd0.058012623492682824, 32'sd-0.14523454135506814, 32'sd-0.01780445405567543, 32'sd0.08295281238538699, 32'sd0.07994770636895769, 32'sd0.09515125491683164, 32'sd0.007278136039517123, 32'sd-0.05515495721191325, 32'sd-0.08646112866304115, 32'sd0.053353888080520585, 32'sd0.1103379476884151, 32'sd-0.018084446306877337, 32'sd0.14551350545331712, 32'sd0.06754627468736467, 32'sd0.08573651719697967, 32'sd-0.05862641490004648, 32'sd-0.0035707034760918306, 32'sd0.04374819430820498, 32'sd-0.06277702251241098, 32'sd0.03214663927837569, 32'sd0.09828744242930966, 32'sd-0.02082545222519595, 32'sd0.02431407083109913, 32'sd-0.034980455795958446, 32'sd0.06314824448122995, 32'sd0.11703490333289371, 32'sd0.20460863463008153, 32'sd0.05884630204702025, 32'sd0.08817688363137245, 32'sd0.0412683585157595, 32'sd0.03973813451095639, 32'sd-0.04986729472844005, 32'sd0.002505590100939266, 32'sd0.03157189504652505, 32'sd-0.031328444473761985, 32'sd-0.04105852099949466, 32'sd0.004570695124820265, 32'sd0.10216242899358365, 32'sd0.09371703770515434, 32'sd0.038017618608642334, 32'sd0.09592213199044618, 32'sd0.09104674129398248, 32'sd-0.01383995768193219, 32'sd-0.04605350715702916, 32'sd0.04943419577942328, 32'sd1.0445293464753906e-119, 32'sd0.004915309475752125, 32'sd-0.015000729827119256, 32'sd0.07598106156504422, 32'sd0.12203069890904657, 32'sd0.005173560762626141, 32'sd-0.005160867312198126, 32'sd0.09499225203155505, 32'sd0.15608322587989482, 32'sd0.15823782151995078, 32'sd0.04367581970434194, 32'sd0.03430436081657921, 32'sd-0.008008814666923648, 32'sd-0.08891297247365626, 32'sd-0.05678804181647315, 32'sd-0.08133933743862827, 32'sd-0.03290487445296649, 32'sd-0.04908140644441666, 32'sd-0.02366067428998891, 32'sd-0.022656737846229943, 32'sd0.026290270839373752, 32'sd0.12487628732870873, 32'sd-0.016838146758746727, 32'sd0.1750569002598486, 32'sd0.053112960418050234, 32'sd-0.04767852173606947, 32'sd0.04790000243426257, 32'sd-0.03675066041943222, 32'sd-0.07177964675084346, 32'sd-0.06982640507137203, 32'sd-0.06952931764864644, 32'sd0.04377840378762367, 32'sd0.026973603773349012, 32'sd0.05879945471944728, 32'sd0.07907019988015829, 32'sd0.08213288347664459, 32'sd0.03883389656290562, 32'sd0.0631943252032601, 32'sd0.07607018832717494, 32'sd-0.0001565796954974421, 32'sd-0.14026521105912979, 32'sd-0.16356463940981075, 32'sd-0.13549081469191776, 32'sd0.04656654458608574, 32'sd-0.10566419314072609, 32'sd0.0033585824306435995, 32'sd0.04790820036748923, 32'sd-0.07655509419834075, 32'sd-0.021617716625936746, 32'sd0.13348076641761503, 32'sd0.0006823085342288569, 32'sd0.059121789091432266, 32'sd-0.03634122673258959, 32'sd-0.18095998426353965, 32'sd-0.07289485759145983, 32'sd-0.07019848807835868, 32'sd-0.03911777936115062, 32'sd-0.052701299306177216, 32'sd-0.050087350541148004, 32'sd-0.00700296873790852, 32'sd0.049567195439976036, 32'sd0.10299794168519227, 32'sd0.07486554535227395, 32'sd0.017897833741532674, 32'sd0.13928983530275754, 32'sd-0.004031872259332982, 32'sd0.06597790737970627, 32'sd-0.10180665352109407, 32'sd-0.1909788594683363, 32'sd-0.1905645917758542, 32'sd-0.03382589239942226, 32'sd0.043119567419505664, 32'sd-0.037338648886787944, 32'sd0.033101168025270626, 32'sd0.0350557056987784, 32'sd0.08475533528579597, 32'sd-0.0010118900093475376, 32'sd-0.008143247611743119, 32'sd0.13235911582971102, 32'sd0.10592458637164866, 32'sd-0.05170372620140659, 32'sd-0.13873023200378282, 32'sd0.009306906834587462, 32'sd-0.06253894618730287, 32'sd-3.022933416888783e-122, 32'sd0.04743091535661127, 32'sd0.039090502529688056, 32'sd0.02427990746641824, 32'sd0.017632980488027878, 32'sd0.022121665029685208, 32'sd-0.03084568815734225, 32'sd0.06705064777694177, 32'sd0.08330164463457572, 32'sd-0.013814715036652148, 32'sd-0.030876353796177886, 32'sd-0.15310866806947152, 32'sd-0.1436891059219744, 32'sd-0.024135480331091853, 32'sd0.05723154779875615, 32'sd0.06321133518132874, 32'sd-0.04831135949802552, 32'sd-0.10899963524949394, 32'sd-0.08408396024887836, 32'sd0.047492518604578475, 32'sd-0.09561683149261674, 32'sd-0.06484448656635897, 32'sd-0.027222360484015776, 32'sd0.042885586969698256, 32'sd-0.036152902105721946, 32'sd-0.021524800602306573, 32'sd-0.0032234412791600723, 32'sd-0.05578010433993206, 32'sd-0.010574255138042372, 32'sd0.007097418967011165, 32'sd-0.02168737204044003, 32'sd-0.09908372103684622, 32'sd-0.11911224993718114, 32'sd0.026934245247552634, 32'sd0.1122967593491056, 32'sd0.12968236019373797, 32'sd0.05123628705836054, 32'sd-0.063450828169751, 32'sd0.10997423587424762, 32'sd0.07787665783035783, 32'sd-0.035097973262402646, 32'sd-0.07950921353075692, 32'sd0.010772806633272214, 32'sd0.09753664327719044, 32'sd-0.014804285608576278, 32'sd-0.034128184357731316, 32'sd-0.12310122386196286, 32'sd-0.08636832355365322, 32'sd-0.03486198533345298, 32'sd-0.013191549468564821, 32'sd0.024981751468274093, 32'sd-0.06510697336829926, 32'sd-0.007428452839637089, 32'sd-0.11472826866352429, 32'sd0.0010239392715831355, 32'sd0.009077857808984485, 32'sd-0.053815998665100076, 32'sd0.02924402284423218, 32'sd-0.0667280099262455, 32'sd-0.02139213699008055, 32'sd-0.11415978665741484, 32'sd-0.07361854869534035, 32'sd0.11123924794962747, 32'sd0.07640180669922114, 32'sd-0.11443666189896888, 32'sd0.016737384295264494, 32'sd0.05669219535071491, 32'sd0.018662383933800018, 32'sd0.12154052971159457, 32'sd0.007325320569101099, 32'sd0.00884914059724591, 32'sd0.011599037940859341, 32'sd0.05244048987518787, 32'sd0.006602710050900032, 32'sd-0.07650691526688755, 32'sd-0.039222871337944915, 32'sd0.09430571905283718, 32'sd-0.081072076821104, 32'sd0.022237730794124607, 32'sd-0.13030988753228806, 32'sd0.010357432542176026, 32'sd-0.09989410309946821, 32'sd-0.04470763026244669, 32'sd-0.04997860368286272, 32'sd-3.5809927900969033e-119, 32'sd0.026858882945209214, 32'sd0.009564605474393344, 32'sd-0.05423129513441579, 32'sd0.03991605075457584, 32'sd0.07397719009742358, 32'sd-0.09859432581528164, 32'sd-0.024814813407131403, 32'sd0.03407660142381127, 32'sd-0.07546573744939074, 32'sd0.025955695355743522, 32'sd0.10135775833940289, 32'sd0.0923642759284453, 32'sd0.15299056867922706, 32'sd0.004422916185372604, 32'sd0.02017622792267079, 32'sd-0.13180351543354, 32'sd-0.1170424592281939, 32'sd-0.03901078333035011, 32'sd0.16324344780547895, 32'sd-0.013686376112658157, 32'sd0.01846404578824537, 32'sd0.05122316342598794, 32'sd-0.02100972636837216, 32'sd0.06614994725708093, 32'sd0.07285028092298719, 32'sd0.07389244045632433, 32'sd3.964038102723716e-125, 32'sd-3.180007370038339e-122, 32'sd-2.5612200007260566e-117, 32'sd0.060155669541978304, 32'sd0.10768951662625006, 32'sd-0.09392382963911224, 32'sd-0.016358531948861953, 32'sd0.03129744947208251, 32'sd-0.05577570422347183, 32'sd-0.043803741381761685, 32'sd0.010476103602943503, 32'sd-0.05300723184123201, 32'sd-0.04837835925194537, 32'sd0.05271556975302627, 32'sd-0.01102182017162792, 32'sd-0.0015368217849543757, 32'sd-0.051542486009549936, 32'sd0.0727671203403159, 32'sd-0.013789401626050286, 32'sd0.0024008707794828965, 32'sd-0.09397920092608619, 32'sd-0.09164030508703247, 32'sd-0.0771517232705141, 32'sd-0.04350369390706083, 32'sd0.004053710542670425, 32'sd-0.06097446286714607, 32'sd0.0021247538058410237, 32'sd-0.021630511162921823, 32'sd2.763622003253297e-119, 32'sd2.4289722600888156e-124, 32'sd-2.0734523157721593e-126, 32'sd-0.015468071687329438, 32'sd-0.07323300853488326, 32'sd0.030656176411726608, 32'sd0.024852184085483616, 32'sd0.055486363139708575, 32'sd-0.03649045843348742, 32'sd-0.15228263615069285, 32'sd0.1273674336988487, 32'sd0.06469429610277572, 32'sd0.05068688226862004, 32'sd-0.0027088292258791546, 32'sd-0.06449972724111852, 32'sd0.028121066310306753, 32'sd-0.021028252485604738, 32'sd-0.0028652976769647106, 32'sd0.013137681598949121, 32'sd-0.05417462343992253, 32'sd-0.03736138398548056, 32'sd0.012301889627911875, 32'sd0.029606760626772945, 32'sd0.0935053477418475, 32'sd-0.02055791459958667, 32'sd-3.814181145666813e-05, 32'sd-0.06643174656407586, 32'sd-0.03841912216477876, 32'sd-1.0427844932968622e-124, 32'sd-2.4531602519711596e-121, 32'sd-8.155199952544796e-116, 32'sd-2.284487426237737e-125, 32'sd-0.05960993448044977, 32'sd-0.006031311858796529, 32'sd-0.007112020432885854, 32'sd0.047761852759169145, 32'sd-0.07100508019100615, 32'sd-0.08048075568558923, 32'sd0.053137108058277566, 32'sd0.06630978413679951, 32'sd-0.061829610548298095, 32'sd-0.16382158964262553, 32'sd-0.08254326723381442, 32'sd-0.13460144259675202, 32'sd-0.0639800003105325, 32'sd-0.016897946132526445, 32'sd-0.09891212124059677, 32'sd-0.08138337097465406, 32'sd0.10947251532924811, 32'sd0.022972061478736115, 32'sd0.0961606971471119, 32'sd-0.029245157276692944, 32'sd-0.06499174004471789, 32'sd-0.018735000044521933, 32'sd0.02797966222767738, 32'sd4.0168323754294548e-115, 32'sd2.966977252387812e-124, 32'sd-1.2133036284801253e-123, 32'sd7.192911646139456e-116, 32'sd-2.6107160360544517e-126, 32'sd1.7318583634347597e-127, 32'sd-0.0063155267260941615, 32'sd-0.08900484347143793, 32'sd-0.03557782603473878, 32'sd0.011530874358253757, 32'sd-0.02361790818409287, 32'sd0.015407192557061938, 32'sd-8.342267204317693e-05, 32'sd-0.10818970069579655, 32'sd-0.09911334034431883, 32'sd-0.09581578589453868, 32'sd0.17601605819953425, 32'sd0.15934324416940482, 32'sd0.05572334525559087, 32'sd-0.052086965288039154, 32'sd0.03661054892242493, 32'sd-0.1009040188469144, 32'sd-0.0248974197863719, 32'sd-0.09353880726209221, 32'sd0.03311623759015987, 32'sd-0.07414287715400304, 32'sd3.0191500260508925e-118, 32'sd-1.0606860779934843e-122, 32'sd2.5980859825138505e-126, 32'sd-2.279757218095423e-118},
        '{32'sd3.525143547644976e-126, 32'sd-1.693840128536243e-117, 32'sd-3.529745336705862e-126, 32'sd-1.925897881672167e-120, 32'sd-6.524022603593701e-126, 32'sd1.4534673329700308e-115, 32'sd-1.696432720144701e-125, 32'sd7.287059354843195e-115, 32'sd2.148957094920734e-127, 32'sd6.246361781153257e-117, 32'sd3.196442766489245e-126, 32'sd-1.2711077884399134e-115, 32'sd0.1647710104032046, 32'sd0.07292173808096107, 32'sd0.0701057641278798, 32'sd0.07698598470806055, 32'sd-8.050968473172573e-116, 32'sd6.516668346384401e-128, 32'sd6.53583122936966e-116, 32'sd9.949261775178182e-122, 32'sd1.0697884218111216e-115, 32'sd-1.6694763940913213e-122, 32'sd1.3546887783400545e-119, 32'sd-1.611132776007281e-121, 32'sd1.7107051251150124e-125, 32'sd1.0715633508995344e-118, 32'sd2.856568099059957e-127, 32'sd1.198681778607912e-117, 32'sd-5.82309881020053e-122, 32'sd-2.3078772201973304e-125, 32'sd-2.9503949068510062e-120, 32'sd3.6133682409866945e-122, 32'sd0.056293824433530947, 32'sd0.06025468106220562, 32'sd-0.05077244092634294, 32'sd0.01179271493492611, 32'sd0.0742600194900253, 32'sd-0.010178889143546385, 32'sd0.02551197015524827, 32'sd0.055804671697799915, 32'sd0.08905530083913998, 32'sd0.05608263107244354, 32'sd0.09220015075987108, 32'sd0.12203749952213774, 32'sd-0.04137013127576219, 32'sd0.0028783558583356217, 32'sd0.08654538720496309, 32'sd0.0482594140815076, 32'sd0.09557330829707841, 32'sd0.025685984358623182, 32'sd0.061274339028258365, 32'sd0.029403512234003577, 32'sd-3.6777872695861547e-116, 32'sd-3.082580846344072e-122, 32'sd5.413928093166655e-126, 32'sd1.0040436529042689e-123, 32'sd-1.6258697234947202e-127, 32'sd-2.8906026952438884e-116, 32'sd0.04406278069820454, 32'sd0.06884136629490477, 32'sd0.084339903638206, 32'sd-0.05082191583099518, 32'sd-0.06230120861058095, 32'sd-0.10328562327093116, 32'sd0.06070932544399041, 32'sd0.1378696570726533, 32'sd-0.0002854220585035392, 32'sd0.024212836661335342, 32'sd0.06225972166739005, 32'sd0.17410479114433147, 32'sd0.2464460992771179, 32'sd0.1650281135836178, 32'sd0.15968321632432536, 32'sd0.04687876596569616, 32'sd-0.08418466721397722, 32'sd-0.07920349134697673, 32'sd0.016677462687698257, 32'sd-0.00031636975794334946, 32'sd-0.046744504820714065, 32'sd-0.0821527964120717, 32'sd0.03867157857830767, 32'sd0.12376925825874509, 32'sd-1.1544179732462364e-127, 32'sd-8.364660559390657e-121, 32'sd1.0440394004569974e-121, 32'sd1.1871876335019338e-126, 32'sd0.1278503035163955, 32'sd0.014065288442264548, 32'sd-0.03469835164867679, 32'sd0.04838387957416443, 32'sd0.15565851521867413, 32'sd0.11518224778467483, 32'sd0.034061911180472214, 32'sd0.05027056229613497, 32'sd0.03160136690448599, 32'sd0.0016554394899492234, 32'sd0.01969938085969237, 32'sd0.12270033827895556, 32'sd-0.05671747086226272, 32'sd0.0025971869029168815, 32'sd0.057117009872015415, 32'sd0.09792561468072543, 32'sd0.0017707330192462695, 32'sd-0.06171255476716444, 32'sd0.03816208120407176, 32'sd-0.12719517471119215, 32'sd0.0022195230390671017, 32'sd-0.04110447797148951, 32'sd-0.0077381221721839625, 32'sd0.025052586192204126, 32'sd0.04954310335656096, 32'sd-6.863258280333358e-124, 32'sd-1.1950873118335775e-127, 32'sd0.04479774544417649, 32'sd-0.04182091084368677, 32'sd0.001031700329356238, 32'sd0.014748345604004202, 32'sd0.06708545766872662, 32'sd0.09046124925571716, 32'sd-0.04087080708565557, 32'sd0.0770032785404794, 32'sd0.06598720545612013, 32'sd0.025340734079662093, 32'sd0.17739000397199978, 32'sd0.1325107521671456, 32'sd0.20973266903622942, 32'sd0.0698631660969049, 32'sd-0.1233493115899317, 32'sd0.05200523781038393, 32'sd-0.046590078388340596, 32'sd0.12964187346508885, 32'sd0.008026190515886064, 32'sd-0.08701448072150422, 32'sd0.0019420861522586217, 32'sd0.018939267292349446, 32'sd0.12769378702728781, 32'sd-0.0345662933348689, 32'sd0.06459115429204448, 32'sd-0.014351802299427771, 32'sd0.012576476543806536, 32'sd-3.5441099965477226e-119, 32'sd0.06306843401500284, 32'sd0.05782580378658314, 32'sd0.04594282368332575, 32'sd0.052631591672881006, 32'sd0.05584762576896196, 32'sd0.01280378440259344, 32'sd0.07849796440308528, 32'sd0.1529713948556242, 32'sd0.16476602021354544, 32'sd0.09290349777641431, 32'sd0.053603144907210624, 32'sd0.002131877765009306, 32'sd0.0072714599149385035, 32'sd0.02402281316145671, 32'sd-0.11963185362768204, 32'sd-0.10611707019362607, 32'sd-0.0372712982686691, 32'sd-0.0260375549888311, 32'sd0.0537318350494511, 32'sd-0.030049997093757646, 32'sd0.001974894291763019, 32'sd-0.1166663710991535, 32'sd-0.07508369363322957, 32'sd-0.016604162372864408, 32'sd-0.01440728998343339, 32'sd0.026403608891991462, 32'sd0.05376199370555561, 32'sd-7.274217890641038e-123, 32'sd0.07546342909677951, 32'sd0.006450003768906163, 32'sd-0.08119739803915359, 32'sd0.03839174096914528, 32'sd0.008836487347635612, 32'sd0.10722851992101813, 32'sd-0.02897123122896209, 32'sd0.009840663946889514, 32'sd0.11122351999604783, 32'sd0.0024623425516323567, 32'sd-0.051878960358345154, 32'sd-0.0352859297967207, 32'sd-0.0980816670065752, 32'sd-0.08578324327713638, 32'sd-0.0466819411093409, 32'sd-0.18781531951806543, 32'sd-0.11973620957948866, 32'sd0.02526408956605703, 32'sd-0.018610966876698654, 32'sd0.08462566001794566, 32'sd-0.09625972533147334, 32'sd-0.09092279386424461, 32'sd0.010302834872842852, 32'sd-0.0011361986575932784, 32'sd-0.01418194128450222, 32'sd0.023969359026891842, 32'sd0.029333690866048298, 32'sd0.054119341784409504, 32'sd0.03839202146309214, 32'sd0.04112758867860153, 32'sd-0.09385275717750004, 32'sd-0.16208326933751618, 32'sd-0.11953582676976422, 32'sd0.06821488851178689, 32'sd-0.07161467817490644, 32'sd-0.00010031693426285109, 32'sd-0.0746181178569175, 32'sd-0.018511958636046297, 32'sd0.0164765330906072, 32'sd0.08966574579720049, 32'sd0.0059092510288103976, 32'sd0.10141769215786027, 32'sd-0.15224790780541167, 32'sd-0.14496750035274256, 32'sd-0.14883880229659607, 32'sd0.008170482907770407, 32'sd-0.07346924954526975, 32'sd-0.05411755813451896, 32'sd0.04710708606659235, 32'sd-0.10993654469723757, 32'sd0.08498242398568136, 32'sd0.10881857164172355, 32'sd-0.023494529788221297, 32'sd0.061831730890686804, 32'sd0.013010745379978187, 32'sd-0.02410204386069024, 32'sd-0.043843380940259725, 32'sd-0.030555665125834512, 32'sd-0.015882973884109666, 32'sd-0.09114947212395996, 32'sd-0.15623023094895583, 32'sd-0.07755052207688069, 32'sd-0.01465980401553383, 32'sd0.03165444863782907, 32'sd0.009744663204833645, 32'sd-0.07255041879420622, 32'sd0.08415272193819828, 32'sd0.0712069204633497, 32'sd0.12197341251471878, 32'sd-0.02210221272510033, 32'sd0.015468245747225232, 32'sd-0.20533963545770884, 32'sd-0.1585892498684123, 32'sd0.024600774930672583, 32'sd-0.1131418585543828, 32'sd0.028546965183877008, 32'sd-0.03673921535898203, 32'sd-0.008232702533442231, 32'sd0.044465922038557586, 32'sd0.05209195194912349, 32'sd0.07717683294621289, 32'sd0.04666197904478657, 32'sd-0.029497255128439218, 32'sd0.017866247789719923, 32'sd0.12230647971298904, 32'sd0.019194127694127396, 32'sd0.03970231944315231, 32'sd0.005037081941827677, 32'sd-0.09156006709578421, 32'sd-0.07844673321505992, 32'sd0.07161187183260993, 32'sd-0.08016797767487563, 32'sd-0.1706905289596723, 32'sd-0.02925385113397908, 32'sd0.08830437128645101, 32'sd0.150481012921728, 32'sd-0.0015935715408187672, 32'sd-0.02278040008914596, 32'sd-0.23404644372580446, 32'sd-0.1911849801959681, 32'sd-0.06328901983964502, 32'sd-0.0407085842354072, 32'sd0.0191170017454932, 32'sd0.14833910504271663, 32'sd0.0968457782452827, 32'sd-0.016565720894773116, 32'sd-0.058604160370825505, 32'sd-0.08002574363942055, 32'sd0.034267341447235235, 32'sd0.036572629388051656, 32'sd-0.017319949988095558, 32'sd0.0893344642621779, 32'sd0.12563669010902517, 32'sd0.11460094817228472, 32'sd0.054923977411160646, 32'sd0.05387155868315848, 32'sd-0.004634796213463324, 32'sd-0.00814527244156645, 32'sd-0.03731271278179061, 32'sd0.037452984007473086, 32'sd-0.09980214501452742, 32'sd0.08678335918588424, 32'sd0.15778408846541495, 32'sd0.14889369408374606, 32'sd0.04290242568022119, 32'sd-0.1703985572823762, 32'sd-0.2801226082017424, 32'sd-0.13219868165430035, 32'sd-0.031946231361948456, 32'sd0.02436000461310971, 32'sd0.0416334433560939, 32'sd-0.013243688373635725, 32'sd0.05404816559224517, 32'sd0.0508613632132089, 32'sd-0.08190183380278912, 32'sd0.04916990988073866, 32'sd0.09876871804222549, 32'sd-0.010279469992461498, 32'sd-0.08650328578710073, 32'sd-0.02893361390115491, 32'sd0.037331986832602776, 32'sd-0.05079120898973805, 32'sd0.07790738356936612, 32'sd0.0312007885605857, 32'sd-0.026594664871732825, 32'sd0.03264595786253391, 32'sd-0.02593009350131261, 32'sd0.05353829090314043, 32'sd0.11825920144846905, 32'sd0.04351383422545533, 32'sd0.12663449258506226, 32'sd0.010214992234194293, 32'sd-0.06411087853308758, 32'sd-0.1322568159266249, 32'sd-0.20190128515973293, 32'sd-0.1052292390689264, 32'sd0.03655963485773388, 32'sd0.04781251835641648, 32'sd0.09215531302163893, 32'sd0.1121484209887553, 32'sd0.00749202084240254, 32'sd0.05058563544984107, 32'sd0.008065178495909391, 32'sd-0.1279103446495787, 32'sd0.004267187510115875, 32'sd-0.07178174007993257, 32'sd0.044745169320356916, 32'sd0.05065660573338517, 32'sd0.025231339561845437, 32'sd0.023479403149906968, 32'sd-0.09595164436117508, 32'sd0.08909463716381932, 32'sd0.02138907761945738, 32'sd-0.11445161887778349, 32'sd0.04184320112028194, 32'sd0.08308422324948132, 32'sd0.11022866714630776, 32'sd0.11646359127155619, 32'sd0.1667542016153948, 32'sd0.11812928858945573, 32'sd-0.2063692970856047, 32'sd-0.20226502680639002, 32'sd0.009877204889204266, 32'sd0.08052666513102116, 32'sd-0.061167872853128004, 32'sd0.05386230784032315, 32'sd0.013447567763727328, 32'sd0.03843570345069346, 32'sd-0.006563034426702652, 32'sd0.0374192242318752, 32'sd-0.12800688656328713, 32'sd0.00012608152740593148, 32'sd-0.00224194732833496, 32'sd0.05013341586893186, 32'sd-0.06585385934870643, 32'sd0.07298898695197749, 32'sd-0.010378963557401411, 32'sd0.1029142986900703, 32'sd-0.0021589218231317514, 32'sd0.0545937358515657, 32'sd0.011408361622921793, 32'sd0.022262943314539842, 32'sd-0.04666050422757961, 32'sd0.08759127018517507, 32'sd0.03432071604792599, 32'sd0.04969582490155236, 32'sd0.08644318257655505, 32'sd-0.04920077658300959, 32'sd-0.21538735007961823, 32'sd-0.10602048779992788, 32'sd0.024120886290032246, 32'sd0.07870229808770046, 32'sd0.19271793437318493, 32'sd0.028845172291439628, 32'sd0.1105106612540967, 32'sd-0.067530335340273, 32'sd0.09568305821624118, 32'sd0.028809054805671412, 32'sd-0.09743599309928892, 32'sd-0.0374562900930874, 32'sd-0.04871055950903393, 32'sd-0.05219115235740828, 32'sd0.03302791355406948, 32'sd0.050636337429828995, 32'sd-0.02545427422527676, 32'sd0.026519145169297646, 32'sd0.01449471231568783, 32'sd0.057006354417552974, 32'sd-0.07304566285189422, 32'sd0.01572645647948654, 32'sd0.11907651749840685, 32'sd0.13432988789489078, 32'sd-0.0019610347947258597, 32'sd-0.1129468894243853, 32'sd-0.09302870803151995, 32'sd-0.14110644627965888, 32'sd-0.06887595414599555, 32'sd-0.03794393899850079, 32'sd0.09866689648099909, 32'sd0.0837198696608075, 32'sd0.13626265127560924, 32'sd0.07297456040021652, 32'sd-0.0020171414000609922, 32'sd0.07667502580976335, 32'sd-0.062299790833407996, 32'sd0.07203051930691531, 32'sd-0.003055561427207006, 32'sd-0.056275321669370736, 32'sd-0.004723904639257268, 32'sd-0.00883422678209033, 32'sd0.061718176330525634, 32'sd0.05009427021519832, 32'sd0.03169672074331485, 32'sd-0.01694062898933757, 32'sd0.053336424793713366, 32'sd-0.05372714848706701, 32'sd-0.03200636916053689, 32'sd0.08143507333683117, 32'sd0.12466159076941839, 32'sd0.11089222931621415, 32'sd-0.03911550451310419, 32'sd0.004781702476749762, 32'sd-0.12358403967774999, 32'sd-0.16489447399811638, 32'sd-0.10120998001983508, 32'sd0.0280983200164669, 32'sd0.17726634614402031, 32'sd0.07961122975516721, 32'sd0.03376522440661536, 32'sd-0.13687928527116433, 32'sd0.09815522819144436, 32'sd0.1800519082059435, 32'sd0.008144729364159107, 32'sd0.06099386115588935, 32'sd-0.01918010617949231, 32'sd-0.06633085656175172, 32'sd0.09410635862590352, 32'sd-0.10684546077029061, 32'sd0.01731588653741332, 32'sd0.047926811562369234, 32'sd-0.06001682810550237, 32'sd0.08319296588552257, 32'sd-0.012522918611827714, 32'sd0.08274262290957096, 32'sd0.037576568185824236, 32'sd0.1545859249922277, 32'sd0.07087476949327319, 32'sd0.04075509671566342, 32'sd-0.04265400851156395, 32'sd-0.13318646513616741, 32'sd-0.13776323776112095, 32'sd-0.08411921198648724, 32'sd0.009719767769362158, 32'sd0.10910234697233835, 32'sd0.20489541534912642, 32'sd0.23616649245182597, 32'sd0.07968404910715102, 32'sd0.0435890393128808, 32'sd0.08102034158913422, 32'sd0.14068528845319495, 32'sd0.039762259548704354, 32'sd-0.07888792893553216, 32'sd-0.030875282165340797, 32'sd0.022149052548738123, 32'sd0.09876039098142185, 32'sd0.02998350370463386, 32'sd0.06000738522084237, 32'sd-1.8802532012087867e-122, 32'sd-0.014541269197455887, 32'sd-0.021466292253360185, 32'sd0.03312382349729794, 32'sd0.1853360151261256, 32'sd-0.08734339153286107, 32'sd0.0029440633173815223, 32'sd-0.04460568077095483, 32'sd-0.05626999607037482, 32'sd-0.12670487686289994, 32'sd-0.2001144909034323, 32'sd-0.14320355268734336, 32'sd-0.09318725476945723, 32'sd0.1310729781505856, 32'sd0.07995623319410194, 32'sd0.2139161278046574, 32'sd0.13963503675556146, 32'sd0.13805339603259723, 32'sd0.1527662490635455, 32'sd0.1265080653279485, 32'sd0.06978457580082086, 32'sd0.11939607190205621, 32'sd0.01596669347958524, 32'sd-0.006571675246890213, 32'sd0.018377036796447966, 32'sd0.10857032639932991, 32'sd0.07589251656733188, 32'sd0.0007065780453279033, 32'sd-0.032225402997552534, 32'sd0.03837391972803526, 32'sd0.022200149846985765, 32'sd-0.05475479176195075, 32'sd0.13656258352697476, 32'sd0.07587369878926109, 32'sd-0.008226687488402424, 32'sd0.008491917223479868, 32'sd-0.07464639733990346, 32'sd-0.06681674175193986, 32'sd-0.23272400099258927, 32'sd-0.12694631306373344, 32'sd0.030401730700500573, 32'sd0.08296396312401473, 32'sd0.11228424923472827, 32'sd0.11621596649812524, 32'sd0.234315192863541, 32'sd0.14099006215979554, 32'sd0.1970391017090274, 32'sd0.061096380382837726, 32'sd-0.006070862825358539, 32'sd0.07324005268489704, 32'sd-0.07769777694466046, 32'sd-0.03036028755759828, 32'sd0.06514497582933765, 32'sd0.12492034994203109, 32'sd0.053429340651685524, 32'sd0.028296749414330066, 32'sd0.07629200606130893, 32'sd0.0024396618248079547, 32'sd0.021559023313247116, 32'sd-0.11331510981676045, 32'sd-0.015344933937780386, 32'sd-0.0026959820597748916, 32'sd-0.005183632128642236, 32'sd0.04000096591927722, 32'sd0.07071737248575745, 32'sd-0.03573467201097021, 32'sd-0.20878588470871312, 32'sd-0.090493175317191, 32'sd-0.01733144560249251, 32'sd-0.08554393225138518, 32'sd0.09414325921768366, 32'sd0.1300809077436957, 32'sd0.0900955294384123, 32'sd0.11662857728520286, 32'sd0.003345899653143116, 32'sd-0.03773916119761759, 32'sd-0.03306671238336415, 32'sd-0.0002709792317446375, 32'sd-0.007869756344123242, 32'sd-0.05864428159438761, 32'sd0.041369087034235676, 32'sd0.0563900766362289, 32'sd0.013534169237471734, 32'sd0.004916025496155612, 32'sd6.146650287399228e-123, 32'sd0.011033562852543808, 32'sd0.035993560693300286, 32'sd-0.030534567102296996, 32'sd-0.06434771597819625, 32'sd-0.05793204434489491, 32'sd-0.015939202113288954, 32'sd0.07261232449012636, 32'sd-0.022820644612021528, 32'sd-0.0909681403460422, 32'sd-0.0460441434171768, 32'sd-0.05660901382396114, 32'sd-0.02241261956401064, 32'sd-0.12898368590517023, 32'sd0.058441079984521485, 32'sd0.046749536314460306, 32'sd0.10041804394120384, 32'sd0.09619877173692455, 32'sd0.11165717504160179, 32'sd-0.09988935967383834, 32'sd-0.13451436731168698, 32'sd-0.03493114948151885, 32'sd-0.046380250402303314, 32'sd0.06482379029787512, 32'sd0.0923677827461755, 32'sd0.036698941580113935, 32'sd0.02733881138022018, 32'sd-0.014336900658305252, 32'sd0.039401100257847814, 32'sd0.010158834402135782, 32'sd0.03773431197097204, 32'sd-0.0479499242071388, 32'sd-0.06389724991273081, 32'sd-0.016154572925272843, 32'sd-0.00688468381519133, 32'sd-0.02085830764304346, 32'sd-0.06400146751595998, 32'sd0.04928553666108343, 32'sd0.05780618036160132, 32'sd-0.03989632900135403, 32'sd-0.0007162873183298167, 32'sd0.030205432838195156, 32'sd-0.1609630145835419, 32'sd-0.08032916095345166, 32'sd-0.08890746784528124, 32'sd0.008640342682419332, 32'sd-0.005588325157310364, 32'sd0.051163126296770736, 32'sd-0.07347284515443263, 32'sd-0.040982878654173605, 32'sd0.019772642624555387, 32'sd-0.07351559428274236, 32'sd-0.0029859875265329265, 32'sd0.060505906533139836, 32'sd0.019718404442514267, 32'sd0.018579394301555422, 32'sd0.0753907408481112, 32'sd0.020787832512993855, 32'sd-0.036899886491533154, 32'sd0.0855241768219811, 32'sd-0.03725440860873983, 32'sd0.05757045538713509, 32'sd-0.007143259216007687, 32'sd-0.0875032394038952, 32'sd-0.038322890755541184, 32'sd0.05248054063467618, 32'sd-0.02791178296797648, 32'sd-0.14082418229337543, 32'sd-0.09554676493486773, 32'sd-0.08975002017090637, 32'sd-0.1840523696742381, 32'sd-0.038829837754071735, 32'sd-0.02839750391343872, 32'sd-0.09414549843944325, 32'sd0.04362296622599796, 32'sd0.09124362016828148, 32'sd0.08156055770807684, 32'sd0.05484343313632175, 32'sd-0.020697025841099986, 32'sd-0.01005405341874877, 32'sd-0.12569169720695986, 32'sd-0.08508195421029448, 32'sd0.0018500273047104233, 32'sd0.08437796578416566, 32'sd-6.62862277745553e-115, 32'sd0.06877663451493696, 32'sd-0.03395938902374761, 32'sd0.03655948821577288, 32'sd-0.05005866300222775, 32'sd-0.03779937089439215, 32'sd0.01817780960201789, 32'sd0.05067337495145256, 32'sd-0.0686351959956483, 32'sd0.0426501531609473, 32'sd-0.015146627676597073, 32'sd-0.15962844254092476, 32'sd-0.1013096740109791, 32'sd-0.04240777412723759, 32'sd-0.0884031602665361, 32'sd-0.10433523191884123, 32'sd-0.06910284266092023, 32'sd0.0028067570439143075, 32'sd-0.06286550734602325, 32'sd0.0771076110834516, 32'sd0.11726445508605951, 32'sd0.005089779753594165, 32'sd0.049252629249053964, 32'sd0.11430120869875876, 32'sd-0.04062826842828151, 32'sd0.055834510803387326, 32'sd0.04696949254463962, 32'sd-9.633382925851645e-122, 32'sd-2.7483824512823315e-119, 32'sd1.567525073146903e-116, 32'sd0.004958887885027342, 32'sd0.07327617694825417, 32'sd-0.006045769624615327, 32'sd-0.10159913023713936, 32'sd0.006639531366034875, 32'sd0.03011429702435981, 32'sd0.06650207588630923, 32'sd0.07214711135796487, 32'sd0.05946605679724541, 32'sd0.12134348326933116, 32'sd-0.009041237171008151, 32'sd-0.011274510922765164, 32'sd-0.018076900820138977, 32'sd-0.025838314862520338, 32'sd-0.10678133145957004, 32'sd-0.09016122922437246, 32'sd0.0259454980783874, 32'sd0.03489440205662709, 32'sd-0.02353564765722443, 32'sd0.04358615867452636, 32'sd-0.05285915326047164, 32'sd0.025348559617216274, 32'sd-0.052244293858008314, 32'sd0.0836039359081435, 32'sd0.05512108606343826, 32'sd9.331926325841184e-120, 32'sd5.402440529201756e-118, 32'sd-3.0245766085548165e-116, 32'sd0.028103742505873726, 32'sd0.008491738635405172, 32'sd0.006723175192658088, 32'sd0.0013996992699028877, 32'sd0.048431697385744, 32'sd0.04751221971162642, 32'sd0.0016372097813271479, 32'sd0.15853155785476697, 32'sd0.053416064221272735, 32'sd0.033489689993986375, 32'sd0.03869342770652228, 32'sd-0.10397475661957233, 32'sd0.00021498401307551868, 32'sd-0.11357528278682628, 32'sd-0.0195294540131615, 32'sd-0.012962097342980131, 32'sd0.035517588553231026, 32'sd-0.008790717220091428, 32'sd-0.10638415063009365, 32'sd-0.06994939048100392, 32'sd-0.0160048524354986, 32'sd-0.0022493292514855676, 32'sd0.06966887826358552, 32'sd0.05477922604659946, 32'sd0.03284441684188517, 32'sd-7.789930207668379e-116, 32'sd6.886073167978332e-126, 32'sd8.234370205910937e-117, 32'sd1.315564012927728e-126, 32'sd0.06457393706975344, 32'sd0.01931256617620656, 32'sd-0.1454857486181714, 32'sd-0.08602239857576188, 32'sd-0.1065249739851626, 32'sd0.0008455690315284452, 32'sd0.054798143542530535, 32'sd-0.08381274905883422, 32'sd-0.030706844096334167, 32'sd-0.008447135907182407, 32'sd0.045373518669113065, 32'sd-0.06247451573870981, 32'sd-0.10767698599265524, 32'sd-0.08626704066104314, 32'sd0.001443967340328672, 32'sd-0.026013032190388183, 32'sd0.047166381801083644, 32'sd0.04884389422476916, 32'sd-0.01834531346317637, 32'sd-0.020647888389963755, 32'sd0.05095481354829341, 32'sd0.004395742001334539, 32'sd0.056059329509285764, 32'sd1.4818029900676935e-127, 32'sd-1.3092296301516125e-122, 32'sd8.946923864786878e-121, 32'sd3.358810912311843e-121, 32'sd-1.988805857071391e-127, 32'sd-1.2312577558811232e-118, 32'sd0.10080827036301647, 32'sd0.09129143435153832, 32'sd-0.03119596530314137, 32'sd0.07500276736641463, 32'sd0.028388495488249944, 32'sd0.07896186411973738, 32'sd0.021156134287207813, 32'sd-0.03238145119076726, 32'sd-0.02750366976376669, 32'sd-0.04987920843487872, 32'sd-0.0833564860090264, 32'sd-0.09641521491279247, 32'sd-0.07895981024358215, 32'sd0.04380528913546615, 32'sd-0.023180289162959368, 32'sd-0.052882206278483834, 32'sd0.03265965636641009, 32'sd0.025259918202898635, 32'sd0.017245798974866458, 32'sd0.07813303810354066, 32'sd2.5701916493151344e-124, 32'sd-2.3593664610041577e-115, 32'sd1.6491478815884706e-125, 32'sd-5.192189711910885e-126},
        '{32'sd-1.2632119948826054e-118, 32'sd-6.212192474086582e-121, 32'sd5.272827299902052e-115, 32'sd-1.056497547134726e-115, 32'sd6.256767027857393e-115, 32'sd1.0738337622954053e-121, 32'sd1.4295483422493779e-118, 32'sd-5.178511943437897e-118, 32'sd3.3133868384056965e-121, 32'sd2.661263943028022e-121, 32'sd6.584135275690422e-122, 32'sd-2.922239646503552e-127, 32'sd0.11477305173003548, 32'sd-0.008604961997367626, 32'sd0.13133712033815909, 32'sd0.11876757721239382, 32'sd5.673042506691292e-124, 32'sd3.751792178938703e-122, 32'sd1.0469383502943241e-121, 32'sd8.025003013208594e-128, 32'sd-4.922297764105187e-115, 32'sd2.9619261752362764e-116, 32'sd-4.6009549860357564e-120, 32'sd8.766436195277392e-127, 32'sd-1.097824458383773e-122, 32'sd-1.3205479158834292e-118, 32'sd-1.8551043022462763e-117, 32'sd-1.0753033384584543e-122, 32'sd-3.8048904425143626e-128, 32'sd2.665654734626809e-124, 32'sd9.32007172022629e-123, 32'sd4.6953938932054495e-118, 32'sd0.03219730148072553, 32'sd0.05787856354049059, 32'sd0.05235183379009955, 32'sd0.06186958571760502, 32'sd0.010711370019830633, 32'sd0.10099120724617959, 32'sd0.014044711782421792, 32'sd0.09707628098603625, 32'sd0.053493554407512474, 32'sd0.13510162636781037, 32'sd0.03454433947796546, 32'sd-0.035101402509119785, 32'sd0.01643251035591967, 32'sd-0.015833460464553563, 32'sd0.07177596172074156, 32'sd0.07860064020832794, 32'sd0.03626581859516537, 32'sd0.0963121049563851, 32'sd0.011930276789669035, 32'sd0.05372957536878699, 32'sd6.38826114267345e-116, 32'sd3.5798553726081003e-122, 32'sd-2.820177002419549e-125, 32'sd3.2229219164280607e-122, 32'sd9.588459467462813e-121, 32'sd6.889062099427269e-126, 32'sd0.03302351480974692, 32'sd0.04239658500640603, 32'sd-0.04424592922805636, 32'sd-0.037512674893072265, 32'sd0.02616898308248274, 32'sd0.12199209522020775, 32'sd0.12794582949547487, 32'sd0.12935855422917616, 32'sd0.1253355085229376, 32'sd0.12339326874520994, 32'sd0.09635878461379273, 32'sd0.03203735303827327, 32'sd0.10831340186373095, 32'sd-0.04126254160579518, 32'sd-0.027879430190648997, 32'sd0.04201783142248265, 32'sd0.0907035380547175, 32'sd-0.07373099503201261, 32'sd-0.058489535542261877, 32'sd0.07678075808185517, 32'sd0.09333898692766522, 32'sd-0.07712871394004363, 32'sd0.15603277260208176, 32'sd0.04056012432156338, 32'sd-8.150488877992631e-127, 32'sd1.8174343509099506e-123, 32'sd-7.070800728528066e-127, 32'sd-3.4460534497386106e-120, 32'sd-0.03990102226791011, 32'sd0.05711682980452324, 32'sd0.04085528744613543, 32'sd0.05265389143271018, 32'sd0.04909721177650505, 32'sd0.027217765373052278, 32'sd0.05027163283948124, 32'sd0.11136333601662568, 32'sd-0.06563328170162556, 32'sd-0.05348564412951993, 32'sd0.10649709184456703, 32'sd0.017648380646542505, 32'sd-0.02724776370333632, 32'sd-0.06199409140919145, 32'sd0.033697429017667195, 32'sd0.04850701450417253, 32'sd-0.05980753724215671, 32'sd0.013488754229001029, 32'sd-0.03571257977511635, 32'sd-0.028643584091891404, 32'sd-0.016600093406976654, 32'sd0.007807400914583927, 32'sd0.04447591539539362, 32'sd-0.021980396356666966, 32'sd-0.10493573168312237, 32'sd2.1107820037378376e-117, 32'sd-1.2513083396296395e-126, 32'sd0.031191447692091166, 32'sd0.054689970058417435, 32'sd-0.0197453596423577, 32'sd-0.021355122822709488, 32'sd-0.03830961641326224, 32'sd-0.06336851119166613, 32'sd0.05136334344152161, 32'sd-0.015092363940424217, 32'sd0.0701413123119583, 32'sd0.12029289199043292, 32'sd0.09771030955030484, 32'sd-0.01778195879227922, 32'sd0.11546027959575425, 32'sd0.03964285987916159, 32'sd-0.01658747284084377, 32'sd0.03471473408075684, 32'sd0.002563576806857017, 32'sd0.03774406245355098, 32'sd-0.009991375382802797, 32'sd-0.0050136227571538515, 32'sd-0.02409909819424544, 32'sd-0.08470482680892708, 32'sd-0.03927584918360136, 32'sd-0.026754931407634786, 32'sd0.010981111155747505, 32'sd-0.007853234919516743, 32'sd0.06099781811255309, 32'sd1.8876112506135976e-117, 32'sd0.0179725907115296, 32'sd0.06402621456619918, 32'sd-0.004502379284393134, 32'sd0.09267406643909364, 32'sd0.02491691262796336, 32'sd-0.05967270060224607, 32'sd0.023706678976731073, 32'sd0.10127136719452005, 32'sd-0.042231735266521846, 32'sd-0.014765485010884247, 32'sd-0.0749500525089982, 32'sd0.08493473918002659, 32'sd0.12841167322966063, 32'sd-0.06512780531060744, 32'sd-0.027823618941893315, 32'sd-0.03095479382886945, 32'sd-0.16236420241743546, 32'sd-0.08364502899773041, 32'sd0.03555070685686365, 32'sd-0.001798745867058919, 32'sd-0.01753226781557077, 32'sd-0.1368944426428247, 32'sd0.010116021872436803, 32'sd0.048908083869843404, 32'sd-0.017927863622423417, 32'sd0.012839103392751459, 32'sd0.0033305133032357913, 32'sd-4.470160088573217e-126, 32'sd0.06091511138792931, 32'sd-0.08063770941926925, 32'sd0.08137684731096533, 32'sd-0.006844156395001961, 32'sd0.042235430851786465, 32'sd-0.07376970227018664, 32'sd0.02476152072871838, 32'sd-0.050769239650532136, 32'sd-0.014829712287606005, 32'sd0.07239357428818607, 32'sd0.08120356356823769, 32'sd0.05298466871903339, 32'sd0.09748663549887455, 32'sd0.014526775538360844, 32'sd-0.029519352328891146, 32'sd-0.06588711759102382, 32'sd-0.0754324014334323, 32'sd-0.06719979460717532, 32'sd-0.103064121038642, 32'sd-0.00028293364989824104, 32'sd-0.12560448894741147, 32'sd0.011457158930716093, 32'sd-0.11824663079424758, 32'sd-0.04039941451447599, 32'sd-0.06346493579549763, 32'sd0.02231843454540404, 32'sd-0.09853057407875344, 32'sd0.06788478084174673, 32'sd0.08928382143034304, 32'sd-0.10255671864875127, 32'sd0.08335175596216543, 32'sd-0.009503917794816612, 32'sd-0.08454906350602828, 32'sd-0.1371784113116162, 32'sd-0.042869772959470906, 32'sd-0.007020623107195301, 32'sd0.0923612555453764, 32'sd0.009175324575379264, 32'sd-0.011582626441839617, 32'sd0.07302921685449726, 32'sd0.07203909887290005, 32'sd0.03726816984005285, 32'sd0.12995523358774996, 32'sd-0.09589105562444089, 32'sd-0.03453462606113657, 32'sd0.034847079535890606, 32'sd-0.045675301582158094, 32'sd-0.14689462436156905, 32'sd-0.05083628743383114, 32'sd0.02535518087852435, 32'sd-0.030026642895495496, 32'sd-0.18685375101290022, 32'sd-0.026641337259047625, 32'sd0.0737534610955281, 32'sd0.011683253803156214, 32'sd0.08353422613241189, 32'sd0.10704070600825567, 32'sd-0.10509770372830998, 32'sd-0.0003439471939121241, 32'sd0.11274782751628705, 32'sd-0.09408138804798814, 32'sd-0.08114059774976767, 32'sd-0.04673499371444947, 32'sd0.05764857106609883, 32'sd0.025183191154518496, 32'sd0.09880161769737102, 32'sd-0.03539129896056346, 32'sd-0.026150664753799395, 32'sd0.06923049801668624, 32'sd0.06092339901160825, 32'sd0.04777524138799746, 32'sd0.05669739963410401, 32'sd0.004164764801159864, 32'sd-0.11230896846446484, 32'sd-0.018796023490434806, 32'sd-0.05230189332766924, 32'sd-0.03144130446716913, 32'sd-0.135844428695093, 32'sd-0.016083939258083706, 32'sd-0.15525374825699093, 32'sd0.0033147174083254004, 32'sd0.038368888308947136, 32'sd-0.05011143841641864, 32'sd0.01085253004571585, 32'sd-0.015325521953960215, 32'sd-0.04760982303651218, 32'sd-0.07109212915815027, 32'sd-0.05116727650510107, 32'sd0.09540332256056505, 32'sd0.07122616794501828, 32'sd0.05145567939454138, 32'sd0.04814284679204255, 32'sd-0.014574626402038271, 32'sd-0.12050109584509554, 32'sd-0.012741185498468035, 32'sd-0.09339311572137768, 32'sd-0.016021830481951594, 32'sd0.05675524936413545, 32'sd-0.07146721936380322, 32'sd-0.02572546558404731, 32'sd0.046301191240693575, 32'sd0.0025470577675949786, 32'sd-0.08023746153585527, 32'sd-0.10742061035659559, 32'sd-0.035162173816087536, 32'sd-0.0858023356613045, 32'sd-0.09321136240450445, 32'sd-0.014328939019644259, 32'sd-0.055836293084705085, 32'sd-0.036438476268791056, 32'sd0.053629245110727884, 32'sd0.07043152506669102, 32'sd0.06791214580965609, 32'sd0.081773342264173, 32'sd-0.07309443518972898, 32'sd-0.10337077530266893, 32'sd0.07523225482704754, 32'sd0.07446769764883687, 32'sd-0.026792690437848172, 32'sd-0.11627924550841154, 32'sd-0.18834637488402475, 32'sd-0.14580011218738081, 32'sd-0.13283370231492328, 32'sd-0.08622981377986229, 32'sd-0.08976510274541472, 32'sd-0.06040090878742653, 32'sd-0.13103250129230193, 32'sd-0.08286044780027291, 32'sd-0.007436553503197439, 32'sd0.011505820491510013, 32'sd0.06568673416030728, 32'sd-0.059417751837686585, 32'sd-0.0431640344965853, 32'sd-0.1007289583497915, 32'sd-0.05552429603342363, 32'sd-0.007432905088046186, 32'sd-0.07076135901209758, 32'sd-0.08526328230810712, 32'sd0.044909933222204955, 32'sd0.006661070812336623, 32'sd-0.05683275812694933, 32'sd-0.05416387244047572, 32'sd-0.057108529687700284, 32'sd-0.018316202724524135, 32'sd-0.06450866226693468, 32'sd0.04997085931670643, 32'sd-0.11886434560467114, 32'sd-0.0689448135101736, 32'sd-0.19574581033222552, 32'sd-0.0600297745909929, 32'sd-0.17741270689971386, 32'sd-0.256017597146746, 32'sd-0.04876129132846338, 32'sd0.04652650940661038, 32'sd0.09020922969963723, 32'sd-0.06392319628569876, 32'sd-0.10617234906282323, 32'sd-0.06329585341006956, 32'sd-0.13424956112169506, 32'sd-0.03504635295148883, 32'sd-0.008615141365906924, 32'sd-0.031083950936237198, 32'sd-0.04665608815736158, 32'sd-0.03984986800095331, 32'sd0.0723185313037107, 32'sd-0.03817270637885884, 32'sd0.0010584679798219324, 32'sd0.036113990417300706, 32'sd-0.06753323507674594, 32'sd-0.10455073011583098, 32'sd-0.057075452709477635, 32'sd-0.04993675724544559, 32'sd-0.13379937070574474, 32'sd-0.20998541473249926, 32'sd-0.1867830899691432, 32'sd-0.1365521055297516, 32'sd-0.1514923774124687, 32'sd-0.11782966338201711, 32'sd-0.10781210284790416, 32'sd-0.040946686841600244, 32'sd-0.01691575992539355, 32'sd0.23859026483485135, 32'sd0.09336156245386815, 32'sd-0.006939060313391315, 32'sd-0.00013071136423307736, 32'sd0.07193317344186803, 32'sd-0.10306824826630635, 32'sd-0.009750042564961946, 32'sd0.05294915637818535, 32'sd-0.044544438563216965, 32'sd0.01806445432851766, 32'sd-0.05460594909972647, 32'sd0.015012337057935237, 32'sd-0.018415863917215284, 32'sd0.011997590317005901, 32'sd0.06346207039884802, 32'sd0.00550601827544963, 32'sd0.014829657326034506, 32'sd0.0037309849154659176, 32'sd-0.009728549724157567, 32'sd-0.07244481469116953, 32'sd-0.11209334433636671, 32'sd-0.12452840595287469, 32'sd-0.07035923953634862, 32'sd0.011419972452932114, 32'sd0.07286701534650711, 32'sd-0.04502497708157328, 32'sd0.029777121933223082, 32'sd0.055973538583571125, 32'sd0.14892837951214968, 32'sd0.0663220022808894, 32'sd-0.028252531069335108, 32'sd-0.04135753830079024, 32'sd0.055326676338398925, 32'sd0.1004743706069583, 32'sd0.041705744543591085, 32'sd0.07284023232419701, 32'sd0.024495161924403337, 32'sd-0.07674093238846845, 32'sd0.07776914338477423, 32'sd0.07309117920317745, 32'sd-0.048355919441449166, 32'sd0.0257028492177999, 32'sd0.03032179905703149, 32'sd-0.022677217805332626, 32'sd-0.059654852791463264, 32'sd0.07842900427025788, 32'sd-0.04298545704740212, 32'sd0.028427427529961784, 32'sd-0.08142224695709357, 32'sd-0.03212502364131507, 32'sd-0.05157567110502926, 32'sd0.08173709869974863, 32'sd0.09391050823000102, 32'sd0.16541923260354724, 32'sd0.12621061778692935, 32'sd0.03470917231144301, 32'sd0.07913900890733158, 32'sd-0.15472914678423227, 32'sd0.03296845429581107, 32'sd-0.11196803798483017, 32'sd0.015553935218826842, 32'sd0.13736456374036304, 32'sd0.07820720673731571, 32'sd0.08766355984257211, 32'sd0.06447699129413989, 32'sd-0.091210116896212, 32'sd-0.0689197405012285, 32'sd0.025938337228828053, 32'sd-0.10991772473430432, 32'sd0.12126399047766317, 32'sd0.07296455627534354, 32'sd0.020001901515167043, 32'sd-0.02687480821021577, 32'sd0.008967157705370718, 32'sd0.010467933604950028, 32'sd-0.030863135979499537, 32'sd-0.036001231302941826, 32'sd0.07805382366110306, 32'sd0.04279922166687895, 32'sd0.09799511635165654, 32'sd0.15940311580706712, 32'sd0.1960117539110516, 32'sd0.020189622952807195, 32'sd0.08358592889664583, 32'sd0.011095134203989804, 32'sd-0.18276982488787596, 32'sd-0.10464959353367177, 32'sd-0.140979850248267, 32'sd0.04214485267056472, 32'sd0.06317278761961355, 32'sd-0.04538362281348213, 32'sd0.057906885574890196, 32'sd-0.0819287681636461, 32'sd0.021175744833741614, 32'sd0.06238299921688631, 32'sd0.04552194286107394, 32'sd-0.08610942706727553, 32'sd0.019857209536935927, 32'sd0.06993036704028255, 32'sd0.006475573663350398, 32'sd0.03089963325446701, 32'sd0.05338561063687468, 32'sd-0.022697780655723105, 32'sd0.07897292352704431, 32'sd-0.0019564668301514246, 32'sd0.10098909305604202, 32'sd0.07356164978133148, 32'sd0.1183204434549263, 32'sd0.1680085200012612, 32'sd0.0416168258304006, 32'sd0.00936994815147703, 32'sd-0.055946756250553564, 32'sd-0.04047231347129543, 32'sd-0.11743327705235064, 32'sd-0.16818727743761847, 32'sd-0.21783762235314247, 32'sd-0.14102695574313004, 32'sd-0.09265742738407401, 32'sd-0.010369246334831597, 32'sd0.011312059404078735, 32'sd-0.039322938599136846, 32'sd0.03140330271210896, 32'sd0.008685110734948275, 32'sd0.026797637629675082, 32'sd0.04048311500751471, 32'sd-0.030400303108510388, 32'sd-7.595362921849764e-116, 32'sd0.03530680923786458, 32'sd0.013291387966379261, 32'sd-0.08262020939541388, 32'sd-0.14565391983941456, 32'sd-0.08163246681365975, 32'sd0.03493963977757707, 32'sd-0.03390352340001073, 32'sd-0.023210511561991724, 32'sd0.08069857592070832, 32'sd0.13392522022547365, 32'sd0.04716851988218987, 32'sd-0.0205360641426287, 32'sd-0.10898463949316528, 32'sd-0.003070203670724716, 32'sd-0.1360849671040747, 32'sd-0.02671639078978968, 32'sd-0.0697215466315063, 32'sd-0.07626214759718376, 32'sd0.008296514440708357, 32'sd-0.0696104489859189, 32'sd0.08814293168074648, 32'sd0.13175036590360392, 32'sd0.12921300676528497, 32'sd-0.0067285092659756735, 32'sd0.08437800092776751, 32'sd0.03204517412977556, 32'sd0.04831616045558004, 32'sd-0.025687791309387843, 32'sd0.08548634650630593, 32'sd0.02692666370628877, 32'sd0.022800190304715143, 32'sd-0.0456992616527484, 32'sd-0.06639200266768765, 32'sd-0.028850973649089527, 32'sd0.003173551033916373, 32'sd0.0017213015006402376, 32'sd0.03572523613692788, 32'sd0.03963396536014193, 32'sd0.026691516584739294, 32'sd-0.005487761290324942, 32'sd0.10816785183265579, 32'sd0.05387086302981871, 32'sd0.04653627190100645, 32'sd0.03110923036565113, 32'sd-0.016407567582799595, 32'sd-0.045486044972422174, 32'sd-0.044458952217748746, 32'sd-0.04242890565823885, 32'sd-0.016782584181789125, 32'sd-0.002586873664185483, 32'sd0.003679870456890451, 32'sd-0.04718217639941391, 32'sd0.06326095096956844, 32'sd0.05801205675071982, 32'sd0.022946242231867784, 32'sd0.00466944111703012, 32'sd-0.00769721003210881, 32'sd-0.025252001636973578, 32'sd-0.11371650550148414, 32'sd-0.011619969721562484, 32'sd0.0020108893217611547, 32'sd-0.11489000000054822, 32'sd-0.04463952177595059, 32'sd-0.13821874733366143, 32'sd0.039948490250888924, 32'sd0.09285956986911223, 32'sd0.004704441278077987, 32'sd-0.026566639868243938, 32'sd-0.017953237914746033, 32'sd0.0376571674391749, 32'sd-0.03412161315084921, 32'sd0.0998023914871776, 32'sd0.1330473442061001, 32'sd0.04691787232931504, 32'sd-0.13030897444735154, 32'sd0.004592838490368306, 32'sd0.004648534983259883, 32'sd-0.009014059852064044, 32'sd0.03372901804274557, 32'sd-0.044336523935762075, 32'sd-0.07718852976978975, 32'sd0.029587743140834226, 32'sd0.003739500217739221, 32'sd6.354282839673584e-126, 32'sd0.001228893524239719, 32'sd0.005611621050579387, 32'sd-0.03356876014960032, 32'sd-0.10222599071635532, 32'sd0.011718795521780966, 32'sd-0.13657805441960472, 32'sd-0.1352059618607015, 32'sd0.01704902305449365, 32'sd0.051205864074954796, 32'sd0.12803099995843753, 32'sd0.0023786078536171497, 32'sd0.13455100680868456, 32'sd0.12160928943183082, 32'sd0.14070875220764698, 32'sd0.08107143655167016, 32'sd0.054458884827023976, 32'sd-0.020975511818725354, 32'sd0.03844773655166067, 32'sd-0.12436899123300804, 32'sd-0.08657815408467696, 32'sd-0.024868114686246234, 32'sd0.10157045735664483, 32'sd0.06862474510985582, 32'sd0.024900980473840244, 32'sd-0.05192551539341565, 32'sd-0.02405073210332726, 32'sd0.03898143537050889, 32'sd-0.0007100529759816713, 32'sd0.04925706940502636, 32'sd0.014394471262792446, 32'sd0.023902963764116825, 32'sd-0.004984051642141772, 32'sd-0.1393636122101173, 32'sd-0.20410218386419818, 32'sd-0.03030203761514881, 32'sd-0.04068119912100703, 32'sd0.09549500743406783, 32'sd0.12825276419424794, 32'sd0.15095264215027804, 32'sd0.06154396126427061, 32'sd0.14355585210788935, 32'sd0.10633620594814573, 32'sd0.07958538271174653, 32'sd0.06996522117213465, 32'sd0.07936034912500718, 32'sd0.0418641747653847, 32'sd-0.07014368539765763, 32'sd-0.09065092419265178, 32'sd-0.006296093013646136, 32'sd0.04316629431242862, 32'sd0.002154708926362225, 32'sd-0.022983685443896902, 32'sd-0.011264151794126364, 32'sd-0.03296760432416462, 32'sd0.02774666602560213, 32'sd0.08862314258936864, 32'sd0.02214843297033745, 32'sd-0.02264559824714762, 32'sd0.04784117397155621, 32'sd-0.06906602923974146, 32'sd-0.04894653281753249, 32'sd-0.011033706774198859, 32'sd-0.06788300447748008, 32'sd0.007390487901994619, 32'sd0.10664105105716723, 32'sd0.07296863129750342, 32'sd0.0461912572972595, 32'sd0.07123292867940094, 32'sd0.06390050326153783, 32'sd-0.00839831458638208, 32'sd0.10671233530058592, 32'sd-0.053754443433102476, 32'sd-0.09529710723767308, 32'sd-0.02344471605021392, 32'sd0.06518885028154561, 32'sd0.08674899551521736, 32'sd0.07145520159917056, 32'sd0.1266234201300514, 32'sd0.013950204285532394, 32'sd0.015554538748740993, 32'sd-0.028030094539002227, 32'sd0.0006358260021609874, 32'sd0.02306015106126097, 32'sd-1.3675569804084744e-115, 32'sd0.05083165573711474, 32'sd-0.027690332017908194, 32'sd0.02519070728779492, 32'sd-0.06839202833169422, 32'sd0.04508785397835571, 32'sd-0.0023162969729203712, 32'sd-0.1037944722938346, 32'sd-0.030041599529707814, 32'sd0.05609726550148109, 32'sd0.08328124695947724, 32'sd0.044214109380483264, 32'sd0.026133634984120906, 32'sd0.07341700536922653, 32'sd0.03033811993219861, 32'sd0.009982807581956231, 32'sd0.09528536629154094, 32'sd-0.019067446450980678, 32'sd-0.11717697793965759, 32'sd0.06396560859087973, 32'sd0.07732510553427484, 32'sd0.020635361593963425, 32'sd0.009961205179931478, 32'sd-0.04939506294139287, 32'sd-0.12922583453759293, 32'sd-0.07683771447724876, 32'sd-0.0065236074793059195, 32'sd1.1652773589123896e-115, 32'sd-1.028853043136807e-121, 32'sd-3.748102086692695e-125, 32'sd-0.048099067169002446, 32'sd0.006941042682043252, 32'sd0.02764923679682711, 32'sd-0.04378909695857376, 32'sd-0.15025478647725285, 32'sd-0.08307415371815544, 32'sd-0.13969315678626038, 32'sd-0.05904056792711762, 32'sd-0.06596450519473786, 32'sd-0.04807620872212205, 32'sd0.014925356004403574, 32'sd-0.018247569321976898, 32'sd0.0396248020850006, 32'sd-0.1488232572026946, 32'sd-0.07969097252348237, 32'sd-0.04992631802633285, 32'sd0.006354365699504653, 32'sd0.001727525967722831, 32'sd0.03658792192083506, 32'sd-0.07266596459282035, 32'sd-0.03286919283710404, 32'sd-0.11006005091256103, 32'sd-0.11957806733173834, 32'sd0.09197643990486112, 32'sd0.04397688666311039, 32'sd-1.47073801808452e-125, 32'sd-5.882615344212454e-116, 32'sd1.1801779396655673e-122, 32'sd0.05495299442463913, 32'sd-0.01190958628398516, 32'sd0.014167489014865973, 32'sd-0.05168599661532712, 32'sd0.02893817077362166, 32'sd0.0008455083055439099, 32'sd0.028632271872844877, 32'sd-0.10386257958275309, 32'sd-0.055471764430378635, 32'sd0.09830248225656453, 32'sd0.10824660779905697, 32'sd-0.04948804600379477, 32'sd0.006307250788623148, 32'sd-0.18998779924956702, 32'sd-0.02065513561306184, 32'sd0.017475517450536673, 32'sd0.08705582707430845, 32'sd-0.08150743352768369, 32'sd0.06962377040920885, 32'sd-0.016791166975461673, 32'sd-0.1520436626700795, 32'sd-0.15508229247885238, 32'sd0.03563985324096545, 32'sd0.04829683601534712, 32'sd0.03166795644739569, 32'sd1.2108285115748392e-118, 32'sd-2.812350004645831e-123, 32'sd2.3642883400113497e-120, 32'sd1.0513488058240353e-124, 32'sd0.05107973926068816, 32'sd0.02572555036296623, 32'sd0.045336703659489205, 32'sd-0.029332565105962487, 32'sd0.0020933676161752706, 32'sd0.09383213643783299, 32'sd0.03299025604764448, 32'sd0.06356596684641697, 32'sd-0.005293841337644102, 32'sd-0.09235170245960533, 32'sd-0.06109851716769185, 32'sd0.02283155041793886, 32'sd-0.00045505256102045536, 32'sd-0.01663148157649815, 32'sd0.02504666551197397, 32'sd0.06627810909274147, 32'sd0.005626615302601489, 32'sd-0.09817930954588582, 32'sd-0.020374357871178722, 32'sd0.030909024195278523, 32'sd0.054780990778190916, 32'sd-0.06122457856978755, 32'sd0.05180996613682335, 32'sd-2.0588252755033167e-117, 32'sd1.2522446153429601e-127, 32'sd1.506443175871455e-123, 32'sd-3.410120164577566e-122, 32'sd-2.0983557049202707e-115, 32'sd2.111655180359786e-123, 32'sd0.05333176480529639, 32'sd0.03336762916565186, 32'sd0.0713844940875065, 32'sd0.0591338386693144, 32'sd0.048102420138897685, 32'sd0.06278865829813465, 32'sd0.003073319870962174, 32'sd0.03246464466267818, 32'sd0.08158823727942643, 32'sd0.02901952712972267, 32'sd0.025935647965202552, 32'sd0.07884669707768283, 32'sd0.016814950663790955, 32'sd0.05845642139468718, 32'sd-0.021324219906411136, 32'sd0.00017987218780637923, 32'sd0.007984945891316035, 32'sd-0.07293636806704053, 32'sd0.05202451427871185, 32'sd-0.008317033343780629, 32'sd1.2291154369230574e-125, 32'sd5.872513930269198e-117, 32'sd6.140387766738671e-122, 32'sd2.0860619587894913e-117},
        '{32'sd2.9313017561411223e-120, 32'sd2.3360499178175216e-123, 32'sd-1.0617023602828847e-124, 32'sd1.1250056314533696e-122, 32'sd2.63554063687015e-119, 32'sd-4.583025128570006e-120, 32'sd-9.589555386655525e-125, 32'sd2.600366129654179e-126, 32'sd-1.096288425529853e-115, 32'sd3.333265754382256e-127, 32'sd-1.7738670756923004e-117, 32'sd3.3515433409414926e-122, 32'sd-0.002688758718231045, 32'sd-0.05060010359254344, 32'sd0.03820214540240084, 32'sd0.07963422177801574, 32'sd4.438244619359013e-122, 32'sd6.8292660883912774e-127, 32'sd-1.2495021379400236e-122, 32'sd-2.7508757997410616e-118, 32'sd-3.274551334133792e-119, 32'sd7.5611574482267765e-115, 32'sd-1.6698994747134124e-127, 32'sd-2.2432226415279992e-123, 32'sd-5.57497207315024e-115, 32'sd-2.219590984359807e-118, 32'sd3.6478636167658804e-116, 32'sd-3.395468102630127e-120, 32'sd-9.8129963750385e-127, 32'sd2.8941421680084875e-115, 32'sd-4.2973923148157234e-125, 32'sd1.3713026577342463e-121, 32'sd0.07196273752291675, 32'sd0.05148984468125656, 32'sd0.011261480505607152, 32'sd-0.02419171997230052, 32'sd0.056637959061152716, 32'sd0.06606843568928039, 32'sd0.04913241819980691, 32'sd0.005390043621349914, 32'sd-0.04460342401462784, 32'sd0.02005567089164763, 32'sd0.012403537713586115, 32'sd0.06303185887641877, 32'sd0.016045103733724385, 32'sd0.039194739890453204, 32'sd0.043323706062261366, 32'sd0.03152117434872604, 32'sd0.07912907021823883, 32'sd0.09215865994790362, 32'sd-0.04385720118542152, 32'sd-0.0015124538127613601, 32'sd-1.1923558641426191e-122, 32'sd1.438501202965997e-125, 32'sd2.7118059388987535e-118, 32'sd-2.1818495160059153e-119, 32'sd-3.1553017571477015e-127, 32'sd-1.0197908946342433e-121, 32'sd0.011608845741643848, 32'sd-0.013784381717804469, 32'sd0.0742371125220075, 32'sd0.04890184062629287, 32'sd0.00815659945427684, 32'sd-0.05516791411620837, 32'sd0.03761463063696357, 32'sd0.042599808292886766, 32'sd-0.03533940796517295, 32'sd0.03886112883415623, 32'sd0.004357298647115225, 32'sd0.052330674049247405, 32'sd0.12324763428355946, 32'sd0.09819630071339061, 32'sd0.06691288879163565, 32'sd0.11276974091516359, 32'sd0.10997249158216874, 32'sd0.13408785801861267, 32'sd0.03546625800623412, 32'sd0.16525851336093872, 32'sd0.09261242891435992, 32'sd0.01576914952835637, 32'sd0.0429149304122266, 32'sd0.06585358936409359, 32'sd-2.016262563697165e-127, 32'sd6.789800464764009e-120, 32'sd8.053380635472189e-124, 32'sd1.036302570877936e-121, 32'sd0.05450527017657402, 32'sd-0.018145372410450878, 32'sd-0.007270254168093677, 32'sd-0.03803300460196371, 32'sd0.06323477830135868, 32'sd-0.1409363688414879, 32'sd-0.0280415759668852, 32'sd-0.005111777946301863, 32'sd-0.1142456574732842, 32'sd-0.011769977970596361, 32'sd0.08293414452823948, 32'sd0.1732023874652036, 32'sd-0.010563305608691459, 32'sd-0.010542387810660131, 32'sd0.0008429625566553766, 32'sd0.13338537176954463, 32'sd0.009299688929645604, 32'sd0.024199431425757357, 32'sd-0.011766692312203165, 32'sd-0.016686767289547315, 32'sd-0.009015411685637856, 32'sd0.044039428483183374, 32'sd0.05934401772497222, 32'sd-0.014423712004335025, 32'sd0.051439246340299845, 32'sd-8.100715838349625e-118, 32'sd-1.678988847513335e-125, 32'sd0.04238570724857934, 32'sd-0.003775731982581644, 32'sd0.013186681773976767, 32'sd-0.037877562447075776, 32'sd-0.0027478650021653703, 32'sd-0.010737525067536988, 32'sd-0.08665582489312157, 32'sd-0.07211097116360711, 32'sd-0.05017179237533146, 32'sd0.010929214860051259, 32'sd-0.04663404467669843, 32'sd-0.07056569009044968, 32'sd0.014848592435090914, 32'sd-0.021029391764236963, 32'sd0.04545480249071853, 32'sd0.07780772763600233, 32'sd0.0556252188482935, 32'sd-0.027735646101721988, 32'sd-0.013286416465135316, 32'sd-0.13105066549856068, 32'sd-0.02381944631306257, 32'sd0.021051665542586653, 32'sd0.013391367852775808, 32'sd0.0022811260622211324, 32'sd-0.0952234178123985, 32'sd0.02333496911236121, 32'sd0.03701877407217549, 32'sd-1.0228074642748839e-127, 32'sd0.018320239980771796, 32'sd-0.06340510468822594, 32'sd0.019692903442491794, 32'sd-0.10774274343179373, 32'sd-0.040524642268454314, 32'sd-0.10972455892013726, 32'sd-0.03824284683159884, 32'sd-0.01986358249716249, 32'sd-0.1791055478026411, 32'sd-0.07595168889394932, 32'sd-0.06793991930522279, 32'sd-0.18918507575430446, 32'sd-0.02632381649365069, 32'sd0.1757186894582572, 32'sd0.1611447391097109, 32'sd0.016826564846388406, 32'sd0.021350036260099525, 32'sd-0.05897174620045077, 32'sd-0.10219294257330507, 32'sd-0.04174077666752582, 32'sd-0.0029656704517059965, 32'sd-0.08463528911418411, 32'sd0.006205576595757523, 32'sd0.05511564213406706, 32'sd0.08043083077392393, 32'sd0.047716518263169715, 32'sd-0.05412394685197404, 32'sd-3.680317920275457e-120, 32'sd0.03338028558318394, 32'sd-0.03546793451122081, 32'sd-0.09989062937760708, 32'sd-0.18802387405983073, 32'sd-0.029319222318224824, 32'sd-0.06483731352130565, 32'sd-0.04813614525735698, 32'sd-0.12959618049182722, 32'sd-0.1258284624813938, 32'sd0.007617944391368918, 32'sd0.014096773321986361, 32'sd0.006235905902625548, 32'sd0.12883920997110637, 32'sd0.16615709685838156, 32'sd0.15135166140773687, 32'sd-0.03562826273911439, 32'sd-0.05814951693027028, 32'sd-0.10343043169510134, 32'sd-0.1905192553018307, 32'sd-0.1428035401866436, 32'sd-0.0825325482396491, 32'sd0.0011404071823229828, 32'sd-0.13140398979811443, 32'sd0.04558454513580522, 32'sd-0.08199940347863295, 32'sd0.02518995940169785, 32'sd-0.12552708963391065, 32'sd0.04061573133344123, 32'sd0.006855928703875608, 32'sd-0.07638122974758033, 32'sd-0.026259170264515175, 32'sd-0.033381249408310325, 32'sd-0.04928582227314082, 32'sd-0.024690426587970778, 32'sd-0.07203740833649984, 32'sd-0.03105562940291587, 32'sd0.06768588681746206, 32'sd-0.014561269748498704, 32'sd0.11591372317848196, 32'sd0.1052726288619942, 32'sd0.012341297461816595, 32'sd0.04113504731419889, 32'sd0.13716896928111155, 32'sd-0.026468150483564074, 32'sd0.0114574963586505, 32'sd0.045742903626135895, 32'sd-0.0420503080137502, 32'sd-0.20565746251565126, 32'sd-0.15612347958650152, 32'sd-0.017926994164052072, 32'sd0.012286146756979192, 32'sd0.12036635158134637, 32'sd0.06024167527595078, 32'sd0.01261509363726615, 32'sd-0.08723042639107148, 32'sd-0.004604293444833551, 32'sd0.07662098166492017, 32'sd0.10572538650975229, 32'sd-0.0598129355717662, 32'sd-0.08587778877635106, 32'sd-0.030879265949407275, 32'sd-0.007430612388622816, 32'sd0.004884538997696441, 32'sd0.14563971475009282, 32'sd-0.04976314010270029, 32'sd0.04242728675449793, 32'sd-0.027196678507110054, 32'sd0.017642728428930346, 32'sd0.007162063546275615, 32'sd0.2006061867103664, 32'sd0.24840518535304237, 32'sd-0.04845177691134986, 32'sd-0.02103383362103763, 32'sd0.055354657108962986, 32'sd-0.10080959001123757, 32'sd-0.19994014810439675, 32'sd0.0043816967291087855, 32'sd-0.020125429738033242, 32'sd0.05564132557529052, 32'sd0.06484358183013601, 32'sd0.0755910051782356, 32'sd0.039978472002002136, 32'sd-0.043335472241607845, 32'sd-0.015951206037269947, 32'sd-0.0011943296982075084, 32'sd0.17134236550168144, 32'sd-0.02417415377105783, 32'sd-0.027478846929566092, 32'sd0.08677113565067246, 32'sd0.06711715692296549, 32'sd0.07338479502867953, 32'sd0.045029497877820034, 32'sd0.0036438114487816115, 32'sd-0.062306399393522206, 32'sd-0.12036047320989497, 32'sd-0.08935130693137662, 32'sd0.05137446256011948, 32'sd0.18505780177497175, 32'sd0.05263247009114566, 32'sd-0.0732952062494098, 32'sd-0.06390760191229096, 32'sd-0.07800356327966579, 32'sd-0.06770815598567173, 32'sd-0.004050488245666926, 32'sd-0.009203540835449915, 32'sd0.08745477200737263, 32'sd0.08636087656661458, 32'sd-0.030801610813391812, 32'sd0.07160146036045642, 32'sd-0.043564530728729504, 32'sd0.021510528746828215, 32'sd0.006214444896540003, 32'sd0.004036199275404754, 32'sd0.0785822545365269, 32'sd0.02369392428305564, 32'sd0.045468239327979776, 32'sd-0.012890687051246554, 32'sd-0.011918925068314636, 32'sd-0.02882089610207615, 32'sd-0.10258446763983327, 32'sd-0.18288641670358424, 32'sd-0.2210473790357171, 32'sd-0.1826807232445733, 32'sd-0.02932944128294436, 32'sd0.08467580296062506, 32'sd0.12661212412347495, 32'sd0.11572068747578178, 32'sd-0.06597620730370418, 32'sd-0.08195193035311639, 32'sd-0.1339443185812244, 32'sd-0.09272150032306506, 32'sd0.03300607746830144, 32'sd0.05288748157190298, 32'sd0.1448201576746813, 32'sd0.08775045973653184, 32'sd-0.01638577292641201, 32'sd0.0008388210704563611, 32'sd0.06537675789656101, 32'sd0.08021533495009095, 32'sd-0.035827825206658385, 32'sd0.039779161556081584, 32'sd0.09713840639600897, 32'sd0.07671981309169212, 32'sd0.026478467285703675, 32'sd-0.05952628205560711, 32'sd0.003937195209555193, 32'sd-0.08517661530672171, 32'sd-0.16504112438728086, 32'sd-0.1705575115441677, 32'sd-0.21617990585505223, 32'sd-0.11502049769445753, 32'sd0.12309808003068813, 32'sd0.20900933892263224, 32'sd-0.002931174597785622, 32'sd-0.13415088970337058, 32'sd-0.15381736441049124, 32'sd-0.07255187807872786, 32'sd-0.16795384545215591, 32'sd-0.07652564361056788, 32'sd0.0641176384385244, 32'sd0.00025335613704295824, 32'sd0.12908611730029046, 32'sd0.0338075673236336, 32'sd0.06449210793030781, 32'sd0.06111204384488711, 32'sd0.0005616749019945692, 32'sd-0.05732753558539063, 32'sd-0.014007119015228251, 32'sd-0.01124077556830814, 32'sd-0.03519825412634655, 32'sd-0.051751728680006756, 32'sd-0.03820657713019898, 32'sd-0.11938102634658727, 32'sd-0.10542049885109875, 32'sd-0.09594391922982135, 32'sd-0.20923880202844672, 32'sd-0.14109422343246975, 32'sd-0.04352143637279238, 32'sd0.01154226395518136, 32'sd0.20057762589325556, 32'sd0.09741140537421981, 32'sd-0.07047160281547837, 32'sd-0.20612230406415008, 32'sd-0.22422549230294916, 32'sd-0.04616819380624278, 32'sd-0.03811081783890316, 32'sd-0.0038519432181512267, 32'sd-0.02090294010302905, 32'sd0.07298284509031808, 32'sd0.0695100794748778, 32'sd-0.003038542595707051, 32'sd0.10563990244670475, 32'sd0.036467083886489775, 32'sd0.017102577760606648, 32'sd0.08229406986120862, 32'sd0.014472988971834003, 32'sd0.03549495302661004, 32'sd-0.06532730141453776, 32'sd0.10960863215718984, 32'sd-0.0008470424788002398, 32'sd-0.09563553566960628, 32'sd-0.10264244183652384, 32'sd-0.010541484834496507, 32'sd0.08363656532404697, 32'sd0.04564912317250692, 32'sd0.11864458685363936, 32'sd0.18531069831833533, 32'sd0.12096008136184896, 32'sd0.032419661273775456, 32'sd-0.15121187443261483, 32'sd-0.21706291534377148, 32'sd-0.2071248866472616, 32'sd-0.04842167666149869, 32'sd0.04453426858087564, 32'sd0.11783642542327363, 32'sd-0.05506108087264559, 32'sd0.01531621261416285, 32'sd-0.0001229046805661683, 32'sd0.048552058074258685, 32'sd0.09513277293261402, 32'sd0.029363473910890937, 32'sd0.07323344478923598, 32'sd0.08224614247303944, 32'sd0.0024980853538743453, 32'sd0.025019664166884784, 32'sd-0.028027953942766314, 32'sd-0.02839221684012952, 32'sd0.016675796955781204, 32'sd0.07799209682847699, 32'sd-0.0248000247587122, 32'sd-0.05903499511099343, 32'sd0.05066376930803405, 32'sd0.1255870553537877, 32'sd0.08583614524506525, 32'sd0.095631226063466, 32'sd-0.010832657273516675, 32'sd-0.18360492643752455, 32'sd-0.16612701063091595, 32'sd-0.12347986255659488, 32'sd-0.08242325250109878, 32'sd-0.053087617565025384, 32'sd-0.010137964148894191, 32'sd0.0621964176098696, 32'sd-0.008122497093045715, 32'sd-0.07290768373961222, 32'sd0.0013476893023517925, 32'sd0.020750476378143562, 32'sd-0.00012347968645754146, 32'sd0.04295572785772555, 32'sd-0.03926078477436198, 32'sd0.08018479741762982, 32'sd0.009129676577403914, 32'sd-0.0436682808613578, 32'sd-0.07062633069494212, 32'sd-0.003482750117942484, 32'sd-0.12277433798058518, 32'sd0.022182763473875693, 32'sd-0.02270216080728572, 32'sd0.05008343838875661, 32'sd0.13083145490001838, 32'sd0.11181650503593459, 32'sd0.11476933334661768, 32'sd0.10560936236500675, 32'sd-0.014220234473303972, 32'sd-0.1975505836050371, 32'sd-0.20438333001466746, 32'sd-0.05200270090018927, 32'sd0.04651791047654116, 32'sd0.02923228107273175, 32'sd-0.0013032561623162293, 32'sd0.0248064536452797, 32'sd0.04541582697296768, 32'sd0.059291220925465814, 32'sd0.0870027471718558, 32'sd-0.07527431422941828, 32'sd-0.0033761912234427285, 32'sd0.011536964417722752, 32'sd-0.06989597418710759, 32'sd0.051353696033844064, 32'sd0.01885656225388125, 32'sd0.041565793925170215, 32'sd0.005678997372707455, 32'sd-0.006056118100125468, 32'sd-0.03375274264388658, 32'sd-0.005819276158178773, 32'sd-0.06359717709031586, 32'sd0.07404245373892561, 32'sd0.020501630612881228, 32'sd0.13716436041455707, 32'sd0.1134950476825054, 32'sd0.12319165044684302, 32'sd-0.08964725330589644, 32'sd-0.09882973201354245, 32'sd-0.16306501358255918, 32'sd-0.0022309729500894224, 32'sd0.05168699278473339, 32'sd0.0025210542867161625, 32'sd-0.10186268424747404, 32'sd-0.07941163078461205, 32'sd-0.03885844002984639, 32'sd0.026551563018912656, 32'sd0.07862209297254971, 32'sd0.037217172312366625, 32'sd0.0770043449213511, 32'sd0.04600735557189159, 32'sd0.0360116129457003, 32'sd0.06094598574447507, 32'sd2.492663789046834e-124, 32'sd-0.01510383789200047, 32'sd-0.054959255388781006, 32'sd-0.091797424806818, 32'sd0.03743258874543743, 32'sd0.06638718934443474, 32'sd0.10077660367323145, 32'sd0.007718142136234714, 32'sd-0.059492856949704104, 32'sd0.058967781878566626, 32'sd-0.05022256998678545, 32'sd-0.03453529715072514, 32'sd-0.0028528650827904603, 32'sd-0.07730586322435679, 32'sd-0.03520956673744757, 32'sd0.013235020078603697, 32'sd0.08177680754426021, 32'sd-0.040069418797949535, 32'sd-0.03879170712205264, 32'sd0.036037940495053, 32'sd-0.030744786176366033, 32'sd-0.04578861490155507, 32'sd0.02529251168918913, 32'sd0.022470282900329704, 32'sd-0.02269315169349284, 32'sd0.07209338186119404, 32'sd-0.08691214029176637, 32'sd0.06642708631612042, 32'sd-0.019539157838436457, 32'sd-0.07083962847527232, 32'sd-0.03940143469475267, 32'sd-0.19734346214035245, 32'sd-0.023975929277679525, 32'sd-0.043730114833775625, 32'sd0.013476384301051922, 32'sd0.01728241959471892, 32'sd0.06517259267767785, 32'sd0.15337352325964035, 32'sd-0.0335585722096319, 32'sd-0.03162991356447593, 32'sd-0.09063286442085565, 32'sd-0.06402452332559033, 32'sd-0.12715506815785613, 32'sd0.03990494470789327, 32'sd0.002894544488875275, 32'sd-0.08001019973886438, 32'sd0.06264733101939227, 32'sd-0.0758389344207973, 32'sd0.036309490838859794, 32'sd0.025028675806259375, 32'sd0.08281959385402551, 32'sd-0.060279699455815884, 32'sd-0.02358620964415892, 32'sd-0.04276298907153606, 32'sd-0.1304088311468277, 32'sd-0.042813039608740965, 32'sd0.016404052635425364, 32'sd0.045006784380180256, 32'sd-0.0938824234638588, 32'sd-0.1550580475060216, 32'sd0.03042955253406563, 32'sd0.0471714491354866, 32'sd-0.014623355251575277, 32'sd0.046510366045825355, 32'sd0.09242169361124385, 32'sd0.056811523317426, 32'sd0.037753900245763486, 32'sd-0.012719431322690636, 32'sd-0.053112719851825065, 32'sd0.03386012931436534, 32'sd-0.10538825998568287, 32'sd0.05368683320144061, 32'sd0.06716646874826704, 32'sd-0.043660357413677284, 32'sd0.007470466452041713, 32'sd0.013843586164611826, 32'sd-0.06739800269681404, 32'sd0.05939513345764739, 32'sd0.15900522973853112, 32'sd0.06207959429367826, 32'sd-0.09233115897708938, 32'sd0.04835449305955214, 32'sd-0.022423558037321958, 32'sd-0.057099669366516864, 32'sd-3.538410702995874e-123, 32'sd-0.07540238146107474, 32'sd0.01035837874493754, 32'sd-0.08944345598662638, 32'sd-0.09248593175137881, 32'sd-0.060560318057419266, 32'sd0.0839792033594662, 32'sd0.1996528948973235, 32'sd0.012272085597946113, 32'sd0.15316915023610167, 32'sd0.09260635642687967, 32'sd0.08021501077983387, 32'sd0.13478378360361612, 32'sd-0.025096816868071553, 32'sd-0.04963901740141492, 32'sd0.08224952611384889, 32'sd0.025993150389292573, 32'sd-0.0069739272139860255, 32'sd0.06497943213649772, 32'sd-0.00535966147982957, 32'sd0.1091210340265389, 32'sd0.030045397527364768, 32'sd0.017258642918928365, 32'sd0.07569013880410694, 32'sd-0.10300808608701206, 32'sd0.04195898196827074, 32'sd0.04549785224818813, 32'sd-0.027586664911310857, 32'sd0.018653894482635203, 32'sd0.054148904392192734, 32'sd-0.015048858819229093, 32'sd-0.0871469900746716, 32'sd0.02812838753127792, 32'sd-0.00023793319390441223, 32'sd-0.010716724084897941, 32'sd-0.050364696946622434, 32'sd0.09491262942140996, 32'sd0.042585795996731415, 32'sd0.011763071268753396, 32'sd0.08326878553857522, 32'sd0.07802599311158014, 32'sd0.039970595145399926, 32'sd0.05025228483874861, 32'sd-0.012257696432612953, 32'sd0.03007972495054461, 32'sd0.017321410150490085, 32'sd0.037705600325699154, 32'sd-0.008278791933347884, 32'sd-0.07341429118807194, 32'sd0.05449886621555759, 32'sd0.11973356624738066, 32'sd0.038636097512729096, 32'sd0.021104614252049292, 32'sd0.003964575784715716, 32'sd0.05652639135509126, 32'sd0.010115332514295267, 32'sd0.09901967607817079, 32'sd0.035413932443835505, 32'sd-0.052584728914924786, 32'sd0.0031055704211163456, 32'sd-0.027823831380632373, 32'sd0.06384708937181693, 32'sd0.04289503316189593, 32'sd0.017424844862438605, 32'sd0.12006126740202609, 32'sd0.06989055551422006, 32'sd0.0884474890225944, 32'sd0.03808824124460049, 32'sd0.16373168894896228, 32'sd0.004299806579399168, 32'sd-0.16859809100364936, 32'sd-0.08712833302217311, 32'sd-0.16330248038883086, 32'sd-0.032271354783813065, 32'sd-0.08021014868025612, 32'sd0.01687616213395323, 32'sd-0.07132947579756416, 32'sd-0.06209952465204639, 32'sd0.09994221036894058, 32'sd-0.08180591453881011, 32'sd-0.03642532500363561, 32'sd-0.014433014699678878, 32'sd0.13663949525420474, 32'sd0.06242947804223187, 32'sd9.258753267014289e-125, 32'sd-0.010129486392803972, 32'sd0.08207741795878376, 32'sd-0.14480232891371428, 32'sd-0.016151724567706704, 32'sd-0.06829317236002713, 32'sd-0.033571633283782404, 32'sd0.1332537278334417, 32'sd0.06108412615900618, 32'sd0.07765695183221383, 32'sd0.10603226889514995, 32'sd0.07275614629800516, 32'sd0.1291902497593952, 32'sd-0.12773202110516965, 32'sd-0.18414463888036, 32'sd-0.06061540637465712, 32'sd-0.1264710809952274, 32'sd-0.01630185533402457, 32'sd-0.07670289320944904, 32'sd-0.08163745320494308, 32'sd0.0031597772600749636, 32'sd0.023658039664252794, 32'sd-0.04082843163371374, 32'sd-0.07289177433424204, 32'sd-0.09046857709525874, 32'sd-0.08515645190734362, 32'sd0.06940000579281523, 32'sd2.9152947373504837e-118, 32'sd-1.8817078164860737e-116, 32'sd-8.428378169707815e-127, 32'sd0.04935566093928025, 32'sd-0.04635616699842677, 32'sd0.009626181531086159, 32'sd-0.04443972380475168, 32'sd-0.012164821495439683, 32'sd0.1417540597907269, 32'sd0.10178321091016254, 32'sd0.004147711123909863, 32'sd-0.02694185349338169, 32'sd-0.01076940581531361, 32'sd0.14017432371423333, 32'sd0.0713205173839097, 32'sd0.068891371550164, 32'sd0.011150703841591222, 32'sd0.07543561205049192, 32'sd-0.023952156318225528, 32'sd0.06510309753790768, 32'sd-0.06994501471260844, 32'sd-0.0283128209261342, 32'sd0.03551413280968465, 32'sd0.06944841784926964, 32'sd0.00327684050726355, 32'sd-0.03397476212121883, 32'sd0.048960753245530404, 32'sd0.019698276865771927, 32'sd-2.1067274919915848e-117, 32'sd6.955675148512945e-124, 32'sd1.1308097230568152e-123, 32'sd-0.06045165961802962, 32'sd-0.0037658314726676597, 32'sd-0.13236763017624895, 32'sd-0.05150016227084248, 32'sd-0.028402715203722596, 32'sd-0.1488851081537192, 32'sd-0.10120131875101766, 32'sd0.04807010228252789, 32'sd-0.05567979389198061, 32'sd0.021785094351281505, 32'sd0.009647816684171513, 32'sd-0.012606438182345773, 32'sd0.0369118603769308, 32'sd-0.03388080061961866, 32'sd-0.05585868298241141, 32'sd-0.07963814186781787, 32'sd-0.008176452472100233, 32'sd0.01869528460968002, 32'sd-0.04448352847425879, 32'sd-0.05637231610393929, 32'sd-0.043242567090360194, 32'sd0.01890675223648466, 32'sd-0.12250055005025762, 32'sd0.012121403475307718, 32'sd0.012027608745500446, 32'sd-6.135334784875849e-120, 32'sd2.6725186653179833e-116, 32'sd4.003412823929464e-117, 32'sd-4.642548355070391e-123, 32'sd-0.02302385372195275, 32'sd0.002759649858982522, 32'sd-0.028852397606547585, 32'sd-0.05938470959899635, 32'sd-0.126511126461825, 32'sd-0.10908843999611645, 32'sd0.016048158619317864, 32'sd0.03359772607203593, 32'sd0.07944502444812185, 32'sd-0.08065535249082838, 32'sd0.0404875510304554, 32'sd0.17784045690910996, 32'sd0.08490259539532641, 32'sd0.009717399678887642, 32'sd0.028660693374358077, 32'sd-0.03866513065084094, 32'sd-0.06144663175355087, 32'sd-0.04015872486676443, 32'sd-0.05524034447210688, 32'sd-0.11801788047045049, 32'sd0.008658254676868779, 32'sd-0.015933449214962498, 32'sd0.021399161276003817, 32'sd-2.048655200330604e-123, 32'sd-2.4971476780771603e-121, 32'sd-2.1734584769623024e-129, 32'sd1.1932364709020175e-115, 32'sd5.0903412645017075e-118, 32'sd-9.700653350363623e-116, 32'sd0.03223439029079471, 32'sd0.06275001179903811, 32'sd-0.026780480519919263, 32'sd0.08181678639575973, 32'sd-0.041969380263101014, 32'sd0.03297026744573003, 32'sd-0.01920122314273957, 32'sd-0.09602048671494001, 32'sd0.02362487525035807, 32'sd-0.0006871032866776843, 32'sd-0.06864850946577751, 32'sd-0.056815328045222754, 32'sd-0.028857177803597776, 32'sd0.050484629442009904, 32'sd0.017443458893933204, 32'sd-0.0730974403845754, 32'sd-0.07210634990688695, 32'sd0.05450853871377071, 32'sd-0.020529402480981326, 32'sd0.04767544084916264, 32'sd5.452044507301409e-125, 32'sd2.184366350320381e-124, 32'sd-7.621517806096445e-117, 32'sd8.885005786173608e-121},
        '{32'sd-3.240665501028214e-120, 32'sd4.4012795860065996e-126, 32'sd3.078001508304444e-120, 32'sd-5.038696803742111e-127, 32'sd4.56299337274266e-115, 32'sd7.83483348955286e-127, 32'sd-5.998992121071872e-122, 32'sd1.2412594350549148e-122, 32'sd9.244104026048972e-117, 32'sd3.084064980105206e-120, 32'sd5.900579048319467e-128, 32'sd-1.6266485241329497e-129, 32'sd0.06776540206468787, 32'sd0.02407670691130675, 32'sd0.08870357805314047, 32'sd0.10567450952529756, 32'sd1.1265122361428118e-125, 32'sd-3.0774963290359674e-115, 32'sd-4.027646210561138e-125, 32'sd1.3171894359021536e-124, 32'sd1.9076464554893573e-127, 32'sd-9.711466542317547e-120, 32'sd-1.4449762513919002e-127, 32'sd-4.772102535683861e-126, 32'sd7.696039617037839e-125, 32'sd6.744009337117375e-120, 32'sd-3.437668984000198e-119, 32'sd8.903000179006208e-127, 32'sd-1.4451715530808757e-124, 32'sd9.28869001172705e-116, 32'sd1.187674136071224e-119, 32'sd-7.413865147227947e-125, 32'sd-0.005180823742589016, 32'sd0.06264806789402716, 32'sd0.08883684350714292, 32'sd0.06878110124065273, 32'sd0.14488762444615097, 32'sd0.0921872677940548, 32'sd0.07026831576698277, 32'sd0.00786473221633302, 32'sd-0.05309395561408194, 32'sd-0.0721139096478592, 32'sd0.05406716205789488, 32'sd0.09413466872992723, 32'sd0.04914902822714999, 32'sd0.08042473819594144, 32'sd0.07068586723733547, 32'sd-0.0029778118784716976, 32'sd0.07158436162248613, 32'sd0.019398306527192113, 32'sd0.04728701076599192, 32'sd0.024670520276806517, 32'sd-3.1597315756376816e-127, 32'sd1.208082560478609e-126, 32'sd1.98302687871506e-124, 32'sd1.9443208360014226e-121, 32'sd8.420776511402211e-127, 32'sd8.56204802382248e-117, 32'sd0.03753778812815017, 32'sd-0.06675705226224142, 32'sd-0.01766075141713048, 32'sd-0.03493473266976704, 32'sd0.004895618839252238, 32'sd-0.013419472190571317, 32'sd-0.052166851534449506, 32'sd0.035893878018494994, 32'sd-0.04013378737098, 32'sd0.01384363152414875, 32'sd0.01693368872040713, 32'sd-0.04422809384956522, 32'sd0.050006608675438616, 32'sd-0.006915472943136098, 32'sd0.017339343821592898, 32'sd0.02887892416732262, 32'sd-0.027090280600443738, 32'sd0.1169350521986451, 32'sd0.011272729035705796, 32'sd0.08196058913397217, 32'sd-0.043189787428345894, 32'sd0.014820894548596688, 32'sd-0.024933791638038924, 32'sd0.07897146313354515, 32'sd-2.6271607231712654e-121, 32'sd-1.6890007111944687e-117, 32'sd-2.9215472520836527e-120, 32'sd4.676976183888614e-118, 32'sd0.03519897952018394, 32'sd0.037872584583272764, 32'sd0.03647773903952399, 32'sd-0.026475753883284006, 32'sd-0.028116765654588777, 32'sd-0.05109006452826851, 32'sd-0.1098705853105652, 32'sd-0.029291862225538506, 32'sd-0.008489678738666106, 32'sd-0.11087778973470126, 32'sd-0.15156555962130547, 32'sd0.09741276234550522, 32'sd0.025821492147755396, 32'sd0.08544280049353445, 32'sd0.10136295191879664, 32'sd0.08629912720222847, 32'sd0.12198005363074285, 32'sd-0.07150722704243262, 32'sd0.06774315669497012, 32'sd0.07180729201902848, 32'sd0.0766323586173854, 32'sd-0.007471276557429867, 32'sd-0.01823263416146566, 32'sd0.11464231618003348, 32'sd-0.006310783600915259, 32'sd4.224703118753213e-126, 32'sd8.676329916714895e-123, 32'sd0.026240974423920677, 32'sd0.02809603455970035, 32'sd-0.09145924447347245, 32'sd0.02168367012704453, 32'sd0.02080222606739322, 32'sd0.05548606324992523, 32'sd0.0644626003803633, 32'sd0.08550398329857113, 32'sd0.1163577163009922, 32'sd0.03249144351407616, 32'sd-0.023179176656914446, 32'sd-0.016075509267860416, 32'sd0.10058078638573961, 32'sd-0.11452419759144321, 32'sd0.07104987522969208, 32'sd0.11088092941611126, 32'sd0.06075281541889218, 32'sd0.07143733792866344, 32'sd0.05581404328737195, 32'sd0.10974011434067749, 32'sd0.06355920999305967, 32'sd0.058610377425079914, 32'sd0.03565922803311429, 32'sd-0.023239534780042995, 32'sd-0.02449435250582217, 32'sd-0.03181428059838787, 32'sd0.050727090924935055, 32'sd4.737210974508376e-125, 32'sd0.014991856603223122, 32'sd-0.058054326008616645, 32'sd0.08642170161642822, 32'sd0.11253117315070482, 32'sd0.0690434231941508, 32'sd0.07704208028239425, 32'sd-0.07168441730193967, 32'sd0.05604531290924023, 32'sd0.024052934596300528, 32'sd0.11345705356025848, 32'sd0.05999815923496066, 32'sd-0.022042521870827742, 32'sd0.1702238407299445, 32'sd0.12075698293552153, 32'sd0.11844511237415509, 32'sd0.025572320176195238, 32'sd0.006831876032085212, 32'sd0.07408166578978706, 32'sd0.1945381533515496, 32'sd0.07478651723976788, 32'sd0.08066103344554418, 32'sd0.14585248625370908, 32'sd-0.04909406284191784, 32'sd-0.0871516233057625, 32'sd-0.002346475870379279, 32'sd-0.0037147823006340413, 32'sd-0.03798381041769667, 32'sd2.5415179280112362e-124, 32'sd0.02105065688763607, 32'sd0.00954602659690377, 32'sd0.058999676314781244, 32'sd-0.0442301838800051, 32'sd-0.022337994516456853, 32'sd0.06181309930319304, 32'sd0.12857759748254446, 32'sd0.057980401089239623, 32'sd0.12627295398160118, 32'sd0.07432745914580798, 32'sd0.10894649781179033, 32'sd-0.031383306451824466, 32'sd0.005697401813897483, 32'sd-0.12670520827589915, 32'sd0.09201048108216468, 32'sd0.07549286392843754, 32'sd0.10610451584910004, 32'sd0.07238358231172264, 32'sd0.13635050352907344, 32'sd0.12258864821457673, 32'sd0.014063502022822949, 32'sd0.037721107437761615, 32'sd-0.060570696688671974, 32'sd-0.022653068061970465, 32'sd-0.0034447083332071627, 32'sd-0.06505764720032353, 32'sd0.03184359872865716, 32'sd0.06945221685245817, 32'sd-0.05842342631853409, 32'sd0.023623556653943036, 32'sd-0.06141342710347416, 32'sd0.07355658263427083, 32'sd0.0904555004593026, 32'sd0.15565166647588133, 32'sd-0.013590235339597963, 32'sd0.0027773348487436307, 32'sd-0.027793188677161084, 32'sd0.16344482466958501, 32'sd0.05256106008699197, 32'sd-0.031180194790527648, 32'sd-0.034277902444321336, 32'sd-0.11356840574561945, 32'sd-0.05939656351172965, 32'sd0.053608771118231216, 32'sd0.06223731366951034, 32'sd0.027557315743778038, 32'sd0.05393461363792984, 32'sd0.06502811355488224, 32'sd0.037431037663202, 32'sd0.067139096227876, 32'sd-0.014446319904069204, 32'sd-0.02473158590917092, 32'sd0.03642954833815239, 32'sd-0.05477010059293085, 32'sd0.00524132032219, 32'sd0.06423871129113412, 32'sd0.06375930890943234, 32'sd0.09474710215128247, 32'sd-0.05914423548746257, 32'sd-0.025774018687011534, 32'sd0.17979479525991324, 32'sd0.08423538236311859, 32'sd-0.048738383272110025, 32'sd0.07050739281490812, 32'sd-0.05078823549684757, 32'sd0.0001311715459795713, 32'sd-0.04794124782563018, 32'sd-0.1337835446495903, 32'sd-0.15852637030364308, 32'sd-0.06126675921130122, 32'sd0.07860260491774926, 32'sd-0.07779834084487863, 32'sd-0.00733625237585327, 32'sd0.08615685334216959, 32'sd0.05662839055708095, 32'sd0.060539625994445595, 32'sd0.06962786126235206, 32'sd0.031088922113054147, 32'sd0.023689969586137435, 32'sd-0.060911181639753065, 32'sd-0.013700649387261874, 32'sd-0.07170385201887713, 32'sd0.02814527176056745, 32'sd-0.018590065393432016, 32'sd0.05030380939509467, 32'sd-0.06839661920781628, 32'sd-0.15730763384780186, 32'sd-0.01372011205908838, 32'sd0.0003873454882936999, 32'sd0.0035903728542301112, 32'sd-0.0011655850778995499, 32'sd0.11870706398670257, 32'sd0.0021346407642312544, 32'sd0.015523777219978508, 32'sd-0.0716576252986682, 32'sd-0.17457498234688415, 32'sd-0.03406401078797121, 32'sd-0.13611791660021513, 32'sd-0.07917942865739837, 32'sd-0.20586917241772626, 32'sd-0.08161033947327384, 32'sd-0.027275337845681293, 32'sd-0.005643273223303845, 32'sd-0.046386134873998175, 32'sd0.06411913353135776, 32'sd0.018651048986473906, 32'sd-0.09479812660402198, 32'sd-0.029084897691627618, 32'sd0.07184238842725967, 32'sd-0.02803553988984342, 32'sd0.03455707265304665, 32'sd0.03138451389689034, 32'sd0.014667698315320821, 32'sd0.08708108145174438, 32'sd-0.05155758232166133, 32'sd0.13514059191056638, 32'sd-0.01906342035142479, 32'sd-0.03161357129451335, 32'sd0.024186834537695014, 32'sd0.1111098608068568, 32'sd0.07941403276883092, 32'sd0.0472697345073487, 32'sd-0.0797352044902002, 32'sd-0.10036694528303979, 32'sd-0.2118065701150333, 32'sd-0.19581856299479516, 32'sd-0.19240316914854186, 32'sd-0.17396885684873659, 32'sd-0.1322608787576082, 32'sd-0.12225057498028098, 32'sd-0.15084142122674338, 32'sd-0.19068246094668193, 32'sd0.07081522437207234, 32'sd0.025614517501815745, 32'sd-0.004896287736825556, 32'sd0.03436488821040707, 32'sd0.05894349915996314, 32'sd-0.08872353558100575, 32'sd0.022328807311546503, 32'sd-0.0654108837028816, 32'sd0.059699403235155296, 32'sd0.10297472014983754, 32'sd-0.03901233228657122, 32'sd-0.06738359872333341, 32'sd0.01385529531476435, 32'sd-0.010675858496442148, 32'sd0.05469880839422502, 32'sd-0.09034043459000804, 32'sd-0.050692468861976064, 32'sd-0.08210535983936458, 32'sd-0.2046817237119232, 32'sd-0.0975293927922182, 32'sd-0.20698416247310514, 32'sd-0.22006228229760283, 32'sd-0.25261645897910046, 32'sd-0.16031105584995728, 32'sd-0.15092996082201424, 32'sd-0.09190363977470269, 32'sd-0.15821369540266073, 32'sd-0.14982385593419367, 32'sd-0.003110190748023571, 32'sd0.03814491090720061, 32'sd0.10343829358041749, 32'sd0.0700757109758764, 32'sd-0.05117122396552156, 32'sd-0.09238478223103432, 32'sd0.04587525132551279, 32'sd0.022564257845749423, 32'sd0.052560707315619556, 32'sd-0.02757549302264631, 32'sd0.07632473489805303, 32'sd-0.08102214929017298, 32'sd-0.003444286297488722, 32'sd0.03908932546981935, 32'sd0.07534929677510106, 32'sd0.014959397012598246, 32'sd-0.0914008742678363, 32'sd-0.048448971606251535, 32'sd-0.12944569221565136, 32'sd-0.0823859388522039, 32'sd-0.2254757747841496, 32'sd-0.1737864220899649, 32'sd-0.16625146387066295, 32'sd-0.09605355335387943, 32'sd-0.06717652252573203, 32'sd-0.21458990415090437, 32'sd-0.014376104792183752, 32'sd-0.03302365035330528, 32'sd-0.0010470633011244036, 32'sd0.06646655561043857, 32'sd-0.06875902599921382, 32'sd-0.01236682142567848, 32'sd-0.04443240074347073, 32'sd-0.03756888508246696, 32'sd0.09179060491104576, 32'sd0.027993459492136358, 32'sd-0.00949254225426792, 32'sd0.05327743207245217, 32'sd0.10332873843153782, 32'sd0.10946126748955567, 32'sd-0.015272510525999186, 32'sd-0.006550653464553599, 32'sd-0.04514925060821941, 32'sd-0.03226088022283908, 32'sd-0.09221866510937887, 32'sd0.013746185703034628, 32'sd-0.01903014970801248, 32'sd-0.1534204648901737, 32'sd-0.14780605588767906, 32'sd-0.12859870814361693, 32'sd-0.12294999106366249, 32'sd-0.07481505999466231, 32'sd-0.029983510932389174, 32'sd-0.10197045714501264, 32'sd0.058672297721640426, 32'sd0.008620729775797042, 32'sd0.0986589337740321, 32'sd0.09887253086871998, 32'sd0.03203301501048326, 32'sd-0.04155400756854403, 32'sd0.03474632304748105, 32'sd0.012496878871746832, 32'sd0.09967252475518311, 32'sd0.09693525526324856, 32'sd0.032675778969016946, 32'sd-0.03443123597648443, 32'sd0.05967026542661951, 32'sd0.047282118186344244, 32'sd0.07828349009837883, 32'sd-0.030261049633378494, 32'sd0.07727875801789005, 32'sd0.061339822665080514, 32'sd-0.0030314478572134227, 32'sd0.006622083383188942, 32'sd-0.02824214482181797, 32'sd0.029181353340589623, 32'sd0.08396117950259577, 32'sd0.07732633165257204, 32'sd0.037183343650140505, 32'sd-0.11373970312378397, 32'sd-0.02526580245549448, 32'sd-0.021654486617336394, 32'sd0.04944142335367599, 32'sd0.1253659088169299, 32'sd0.09660171922273635, 32'sd0.037462482886981625, 32'sd0.00036007436658738555, 32'sd0.05032845882074473, 32'sd-0.007552724250836088, 32'sd0.11211244446995575, 32'sd0.03420026320380839, 32'sd0.11304808759610414, 32'sd0.05911188722156361, 32'sd0.04945799647742169, 32'sd0.04684495462972143, 32'sd-0.01048665111115588, 32'sd-0.048009190673418925, 32'sd-0.026131967923215087, 32'sd-0.06694463736707718, 32'sd0.04259317337658216, 32'sd0.10078709903694232, 32'sd0.020921422608987304, 32'sd0.009927189637097432, 32'sd0.01412671868017608, 32'sd0.033074153977239326, 32'sd0.04188265931616959, 32'sd0.022912188354264094, 32'sd-0.08709677165137653, 32'sd-0.06236051471904174, 32'sd0.059831195868660876, 32'sd0.14418299190683356, 32'sd0.04682476600387682, 32'sd0.13604988549600502, 32'sd0.09308452450979439, 32'sd-0.06522549847351498, 32'sd0.03137865649254227, 32'sd0.0661034872346219, 32'sd-0.00034258634150552723, 32'sd-0.03402207592652362, 32'sd0.02462873443540521, 32'sd-0.060790076852675415, 32'sd-0.037459913049981156, 32'sd0.017158779692601614, 32'sd0.03785914885921072, 32'sd0.043246314926405446, 32'sd0.03913103620301927, 32'sd-0.03399736469735068, 32'sd-0.005289526385165513, 32'sd-0.03667070824433848, 32'sd-0.06918853427708609, 32'sd0.007522083943752863, 32'sd-0.08061689572110187, 32'sd-0.06749934446439111, 32'sd-0.05923589102677276, 32'sd-0.1410131976331141, 32'sd-0.20392081608586646, 32'sd-0.15322868426584785, 32'sd0.0414495254518439, 32'sd-0.017223021135021537, 32'sd0.13704699230733508, 32'sd0.1537201338220622, 32'sd-0.03206056384168175, 32'sd-0.04611414156643235, 32'sd-0.10105633540650344, 32'sd0.04173065844097361, 32'sd0.07867304758205279, 32'sd-0.015690523307676518, 32'sd-1.18966173708401e-115, 32'sd-0.09039968443076929, 32'sd-0.12049633936235322, 32'sd-0.015874357784288716, 32'sd-0.06322904871143573, 32'sd-0.02034251693014082, 32'sd0.11078957690721794, 32'sd0.15826793486649224, 32'sd0.041936774743630195, 32'sd-0.0726592162071078, 32'sd-0.01255218875790153, 32'sd-0.1305599647482046, 32'sd-0.039826913766633776, 32'sd-0.15136633834739027, 32'sd-0.16431074310931587, 32'sd-0.26004206035378236, 32'sd-0.20637881293801555, 32'sd0.02499941424756796, 32'sd0.10182245347387224, 32'sd-0.0034497695240505066, 32'sd0.12276665332106362, 32'sd0.01312250739591902, 32'sd-0.023906974019717697, 32'sd-0.06468522606119405, 32'sd-0.028695767028622386, 32'sd-0.014958935824360009, 32'sd0.02144069861379, 32'sd0.07382821306845767, 32'sd0.01821670663711176, 32'sd0.042514568472609315, 32'sd-0.082182739968143, 32'sd0.11015505803561293, 32'sd0.0461678129440564, 32'sd-0.07477889831167638, 32'sd0.1507941655488783, 32'sd0.21250628293160306, 32'sd-0.009524490793376096, 32'sd0.01758935774801351, 32'sd0.13393284794279803, 32'sd-0.08398574361239673, 32'sd-0.11084444137979194, 32'sd-0.19039308425375367, 32'sd-0.13668952945972063, 32'sd-0.14220913348280909, 32'sd-0.018229893664441856, 32'sd0.11518087771569223, 32'sd0.08129022768634193, 32'sd0.02625189570925672, 32'sd0.047381891940005944, 32'sd-0.05640420266203791, 32'sd-0.08509271222014743, 32'sd-0.13648599750098223, 32'sd-0.12753535596420573, 32'sd0.01701246275052848, 32'sd0.0759261950869767, 32'sd0.005909882251844572, 32'sd0.0322400432251717, 32'sd0.0552075084925947, 32'sd-0.07487890962705492, 32'sd0.1256661055027753, 32'sd-0.010238150353930987, 32'sd-0.08418766609165607, 32'sd0.1844359172751793, 32'sd0.090223324824212, 32'sd0.01983741386313445, 32'sd0.12412867388519182, 32'sd0.0437663340510874, 32'sd-0.07721824410243218, 32'sd0.014697791545378177, 32'sd-0.1402977422893857, 32'sd0.03613441223740489, 32'sd0.040818395646669475, 32'sd0.06481367304053531, 32'sd0.06654746085452215, 32'sd0.09219490199120164, 32'sd-0.011990316568534335, 32'sd-0.06650163137297256, 32'sd0.012035329745424572, 32'sd0.08512332607941629, 32'sd-0.07977807994434913, 32'sd-0.008284095238579875, 32'sd0.0011338609534620031, 32'sd-0.016999773730656368, 32'sd-0.09100856025440042, 32'sd6.581071482336339e-125, 32'sd-0.01659596730046565, 32'sd0.00291140856935477, 32'sd0.06554881362162288, 32'sd-0.027798181924364545, 32'sd0.07746736184048213, 32'sd0.14380267648913303, 32'sd0.07570229975800606, 32'sd0.07992144255574675, 32'sd0.11675982760901361, 32'sd-0.013281619257271313, 32'sd0.05690100307113245, 32'sd-0.01470573013902841, 32'sd-0.04159087746407891, 32'sd-0.05904455657703429, 32'sd-0.04652239150390706, 32'sd0.13654230510174883, 32'sd0.17058151518847234, 32'sd0.16319720613693428, 32'sd0.061174879698791054, 32'sd-0.01458377236841608, 32'sd0.09352904477498979, 32'sd0.04399071175143389, 32'sd0.027243570704999127, 32'sd-0.0393346288974756, 32'sd-0.09409570867280394, 32'sd0.010282351092822198, 32'sd0.008975551308194708, 32'sd0.06509559287354465, 32'sd0.06171082572403689, 32'sd0.04053445427101858, 32'sd0.1646830385659133, 32'sd-0.04997196111848175, 32'sd-0.05615677092087981, 32'sd0.08524717960334022, 32'sd0.12455907548640008, 32'sd0.04505798021602537, 32'sd-0.018500650153502954, 32'sd-0.09163902609460627, 32'sd-0.06586151598098837, 32'sd-0.01382927133688308, 32'sd-0.0026178452546771346, 32'sd0.1167868153460381, 32'sd0.05844647258911142, 32'sd0.14927329651815557, 32'sd0.10245769124284107, 32'sd0.019745365077993342, 32'sd0.028142883813963526, 32'sd-0.009968023018779698, 32'sd-0.017775862694613873, 32'sd0.05687183991885041, 32'sd-0.021506006240201006, 32'sd0.08833207241343297, 32'sd0.07512033938884895, 32'sd-0.02405425073505126, 32'sd-0.028018921738711747, 32'sd0.12619028615894007, 32'sd0.08754879815506111, 32'sd0.0005667387471404612, 32'sd0.09443829128409303, 32'sd-0.003244530321049782, 32'sd-0.01814732570291302, 32'sd-0.023577556061188477, 32'sd-0.007303664032874494, 32'sd0.05025312321287429, 32'sd0.03886491256369777, 32'sd0.021681305498294046, 32'sd0.10662561705396359, 32'sd-0.02615787956588689, 32'sd0.11500523084354201, 32'sd0.172223529700139, 32'sd0.10381404313836129, 32'sd0.1598183001071028, 32'sd0.12395117820377177, 32'sd0.13481805162759994, 32'sd0.0575147251835471, 32'sd-0.005801491117122854, 32'sd-0.04264589898689943, 32'sd0.08395792035868223, 32'sd0.11071902721442195, 32'sd0.142813109558638, 32'sd0.018048175921405455, 32'sd-0.014975206541076513, 32'sd0.04158301039899237, 32'sd-3.03394887020631e-121, 32'sd0.07809569715294282, 32'sd0.107350442880922, 32'sd-0.03515147269543502, 32'sd-0.09060767261777691, 32'sd-0.012815743921514525, 32'sd-0.029537075492014314, 32'sd-0.07691303588062093, 32'sd-0.06975438942819043, 32'sd0.1151508586806157, 32'sd0.15379220487403256, 32'sd0.15891325059850028, 32'sd0.11997464559589643, 32'sd0.14973467162852278, 32'sd0.16051508894061278, 32'sd0.05919524045572089, 32'sd0.14176077302927306, 32'sd0.12288762870684547, 32'sd0.09740296328284351, 32'sd0.012626120531059187, 32'sd0.006138889483865777, 32'sd0.040696557538415605, 32'sd0.035769740391531045, 32'sd-0.020254701452638225, 32'sd0.08029030065856406, 32'sd0.06941962890989879, 32'sd-0.02965691110385554, 32'sd7.90453324015144e-116, 32'sd1.0302051382561982e-124, 32'sd1.0289850347827491e-123, 32'sd-0.012309529692344537, 32'sd0.03863412721394797, 32'sd-0.04666662577492928, 32'sd-0.010468695021549993, 32'sd-0.04574456255566794, 32'sd-0.001316545607182459, 32'sd0.06374250351453528, 32'sd-0.05570530550213413, 32'sd-0.049961908546416356, 32'sd-7.326534438984006e-05, 32'sd0.1331478542886261, 32'sd0.15848946101652886, 32'sd0.014299011531461075, 32'sd0.028515046355621278, 32'sd-0.029396089734939925, 32'sd0.02239866875683448, 32'sd-0.049057916685209424, 32'sd-0.03860469442641551, 32'sd0.035141555570305044, 32'sd0.010099418520142006, 32'sd-0.0010931170984358066, 32'sd-0.0003207060430258924, 32'sd0.058787607107765025, 32'sd0.06710748524972686, 32'sd0.034978821132771856, 32'sd-4.8736563400949885e-123, 32'sd1.129097342029341e-126, 32'sd6.366346878032835e-123, 32'sd0.010505699020166839, 32'sd0.0471545682480218, 32'sd-0.0561423852966071, 32'sd-0.03913188216768695, 32'sd-0.05338226329135654, 32'sd-0.007332583774914353, 32'sd0.04869273218198257, 32'sd-0.031126932470952853, 32'sd0.05581680680077605, 32'sd-0.10718817072509006, 32'sd-0.15218202572700276, 32'sd0.04864278422901274, 32'sd-0.0017001153482612244, 32'sd-0.09413302979910726, 32'sd-0.1596114694428621, 32'sd-0.027807442020946305, 32'sd0.12088906812832571, 32'sd0.04346533788655879, 32'sd-0.056807755714951766, 32'sd-0.1315381785741247, 32'sd-0.01003820167825313, 32'sd0.06953207121533975, 32'sd0.03132884503269094, 32'sd0.02179015339819554, 32'sd0.06085542896756886, 32'sd-8.311491919285865e-123, 32'sd-2.6135712826120903e-126, 32'sd-3.743045241008681e-127, 32'sd3.1188663313633034e-120, 32'sd0.07597252545386544, 32'sd0.05713540661321133, 32'sd-0.04676829066046748, 32'sd0.02337019936435559, 32'sd-0.018795863429522518, 32'sd0.007111905115855266, 32'sd0.07527183531247254, 32'sd-0.007994841115108115, 32'sd-0.11896310308686565, 32'sd-0.1216704695656923, 32'sd0.02156898013178349, 32'sd-0.05612037125459343, 32'sd-0.14854805513082164, 32'sd-0.04266049814842687, 32'sd-0.2137423639881859, 32'sd-0.07991727535148815, 32'sd-0.039745423640986356, 32'sd-0.11789850601844819, 32'sd-0.011636214864159522, 32'sd-0.03629988875219671, 32'sd-0.0020717588657507223, 32'sd0.06387462411173968, 32'sd0.004830326037340855, 32'sd1.2640118268854483e-118, 32'sd-2.122425235156819e-121, 32'sd-2.588697693239618e-116, 32'sd1.464529847985974e-120, 32'sd-4.0923160823674976e-125, 32'sd1.2385317905540645e-115, 32'sd0.0807054702940671, 32'sd-0.035336116768873584, 32'sd0.06636266050101354, 32'sd0.029570690178111838, 32'sd-0.023324548018830448, 32'sd0.03886606931835652, 32'sd0.03655504426360724, 32'sd0.05281318242283286, 32'sd0.07748648617876305, 32'sd-0.004712732176412739, 32'sd0.049860743869417544, 32'sd0.0888236543008512, 32'sd-0.013896709610987943, 32'sd0.021251233274080593, 32'sd0.01744356499742246, 32'sd-0.06734974412441906, 32'sd0.06283824480440685, 32'sd-0.027989443442095824, 32'sd-0.03171060108511211, 32'sd0.02956883991971249, 32'sd-3.895188767423505e-119, 32'sd-3.674731163541698e-122, 32'sd2.2219216762585404e-125, 32'sd-1.0761670835812245e-121},
        '{32'sd1.4117942195477076e-115, 32'sd1.3368938554304955e-115, 32'sd2.8702186222436487e-126, 32'sd-3.3585674353920623e-116, 32'sd-1.1236371372917827e-121, 32'sd9.769611380600383e-122, 32'sd-1.915637013071747e-120, 32'sd9.382706106579807e-121, 32'sd-9.110355799764342e-125, 32'sd-5.750901379011186e-115, 32'sd-2.690238065591152e-124, 32'sd-1.069942647835447e-124, 32'sd-0.03469596074344458, 32'sd0.009238310064277444, 32'sd-0.011059752693600248, 32'sd-0.04026176742240364, 32'sd-1.083173327552841e-118, 32'sd4.241619013766339e-127, 32'sd4.2053721058433927e-125, 32'sd2.1067416959929275e-122, 32'sd-2.082568829774215e-121, 32'sd-3.5754004138972235e-121, 32'sd-1.8621091086593783e-127, 32'sd-3.9649265608368336e-122, 32'sd-6.270232954911613e-117, 32'sd-2.116410627518233e-117, 32'sd-2.202418023465433e-126, 32'sd4.051595821958935e-125, 32'sd-1.324052189032389e-122, 32'sd4.249558659570662e-123, 32'sd-5.349192411599794e-118, 32'sd2.554580398685585e-128, 32'sd-0.03129514044859363, 32'sd-0.10700226603352753, 32'sd-0.025862009049350508, 32'sd0.005275337600681409, 32'sd-0.12277916823795221, 32'sd0.0190458409823686, 32'sd-0.06365498154507383, 32'sd-0.07354461437676457, 32'sd-0.017962388474910013, 32'sd-0.040461485169955624, 32'sd0.014695741095446205, 32'sd-0.049279638895291196, 32'sd-0.0673244595754259, 32'sd-0.08267836070778731, 32'sd-0.019023112307613305, 32'sd-0.014831304911860868, 32'sd0.08400202123767793, 32'sd0.01719385920137871, 32'sd-0.05291582220103466, 32'sd0.0005368598391261649, 32'sd2.0519661225982025e-124, 32'sd5.408855863421269e-125, 32'sd-6.175350657341765e-118, 32'sd1.5163542268576845e-123, 32'sd1.3506867781909e-118, 32'sd2.1078126434356984e-122, 32'sd0.006378557252295727, 32'sd0.03069199998934296, 32'sd-0.03198913877266428, 32'sd-0.023639552121463698, 32'sd-0.04111663370608376, 32'sd-0.03385178996892281, 32'sd-0.046492308889744434, 32'sd-0.017262928369329585, 32'sd-0.12442492896777657, 32'sd-0.04782806806061345, 32'sd-0.016891614549964927, 32'sd-0.030659210174770014, 32'sd-0.10377526820886473, 32'sd-0.009025482066227717, 32'sd0.0367750722727985, 32'sd-0.03622572301854637, 32'sd-0.003687164822186321, 32'sd0.026866339087519876, 32'sd0.011378902871167385, 32'sd0.035544043716016265, 32'sd-0.028855600971015544, 32'sd0.11195422944709808, 32'sd0.07823697394437665, 32'sd1.2441815682141307e-05, 32'sd-1.0778600622939835e-126, 32'sd-3.548982782650111e-116, 32'sd-1.3212258136412756e-122, 32'sd4.2955244652044923e-128, 32'sd-0.03239931749114535, 32'sd0.00868982373261709, 32'sd-0.06865722354031668, 32'sd-0.014729955599598964, 32'sd0.0223428929647035, 32'sd-0.07566458661093486, 32'sd-0.08129834008114933, 32'sd0.04365029671780554, 32'sd-0.07244104927907509, 32'sd-0.14079429513526848, 32'sd-0.09372294837370737, 32'sd-0.19091935195779575, 32'sd-0.18099999904830125, 32'sd-0.10792201612621424, 32'sd0.15956684613642494, 32'sd0.14251242047577073, 32'sd0.07482759562709668, 32'sd0.004410416478002794, 32'sd-0.1262373376272488, 32'sd-0.08323908981278648, 32'sd-0.03217733569299241, 32'sd-0.02882332333806656, 32'sd-0.029604263003309296, 32'sd-0.02427268639743643, 32'sd0.021059236787206004, 32'sd8.312083610390825e-125, 32'sd-3.1399072585307964e-124, 32'sd0.05221493172490639, 32'sd-0.029538334035862236, 32'sd0.05269798619858627, 32'sd0.027146863264662008, 32'sd0.03901639109209571, 32'sd-0.07451045232673546, 32'sd-0.08469812171643663, 32'sd-0.050544652534782075, 32'sd-0.0026986202105801237, 32'sd-0.02827346644933179, 32'sd-0.04373233712250373, 32'sd-0.0846811157541598, 32'sd-0.1939614225793293, 32'sd-0.10855985211050155, 32'sd-0.06766181512561871, 32'sd-0.04776117750914246, 32'sd0.052366425935215365, 32'sd0.016204124622723214, 32'sd0.023287983988404325, 32'sd-0.10350269237888507, 32'sd-0.08022033464137472, 32'sd-0.17439891917983852, 32'sd-0.20858399629781726, 32'sd-0.14074953183860114, 32'sd0.053926417728772866, 32'sd-0.105370796292209, 32'sd0.04670050370599013, 32'sd-8.50169224413204e-120, 32'sd-0.0007847994982116549, 32'sd-0.03053863780816876, 32'sd0.001171783221073884, 32'sd0.03609382101774484, 32'sd0.0320901274374676, 32'sd0.041439277831183174, 32'sd-0.0322067373496605, 32'sd0.08137479606596103, 32'sd-0.007137420083831034, 32'sd0.11327599007467141, 32'sd0.11767924366645297, 32'sd0.038550505304272197, 32'sd0.09068603636877137, 32'sd-0.004711230602764603, 32'sd0.014517900185803696, 32'sd-0.06920363751353384, 32'sd-0.10693582851455818, 32'sd0.01438284291325534, 32'sd0.038908041818744264, 32'sd-0.09493832102270074, 32'sd-0.011005365335055172, 32'sd-0.11248849385060468, 32'sd-0.03094285327137837, 32'sd-0.02483090313546802, 32'sd0.04983650806551961, 32'sd-0.001460598446156618, 32'sd0.005210140232456165, 32'sd2.948513739153002e-125, 32'sd-0.04376857895007163, 32'sd0.011596885423643982, 32'sd0.006847620147691114, 32'sd-0.09683779549789763, 32'sd-0.03377913054125415, 32'sd0.04110538597635078, 32'sd0.014090901802243722, 32'sd-0.021547459121425885, 32'sd0.03382024422400085, 32'sd0.015163385574254186, 32'sd0.07528663636969957, 32'sd0.07812265635674162, 32'sd0.07817072063743213, 32'sd-0.022554478558932563, 32'sd-0.05492130540664344, 32'sd-0.06804660401125906, 32'sd0.03172583989781015, 32'sd0.0224072958403468, 32'sd0.1226847927711871, 32'sd0.04759035645942051, 32'sd0.17081857725455715, 32'sd-0.10086046085694128, 32'sd-0.017714925561851946, 32'sd-0.07462887554220642, 32'sd-0.005850792328253539, 32'sd-0.036905161497316236, 32'sd-0.021533993608056416, 32'sd-0.03397112421252305, 32'sd-0.036328134000113414, 32'sd-0.03265038291679891, 32'sd0.06381110784607763, 32'sd0.015469473813371708, 32'sd-0.06312013542845656, 32'sd0.11289737959398682, 32'sd0.0831181194807045, 32'sd0.04390589804756981, 32'sd0.07808205406984337, 32'sd0.0211329157723791, 32'sd-0.02677719433141947, 32'sd-0.003798884399528897, 32'sd-0.10094024866507995, 32'sd-0.09800140663593661, 32'sd-0.05029707141842713, 32'sd0.10419983796726888, 32'sd0.015435618967786438, 32'sd0.1341460350472342, 32'sd0.08126075635508423, 32'sd0.08075262984448059, 32'sd0.10391117757640117, 32'sd0.02611608691334545, 32'sd0.04040812343990247, 32'sd-0.016180991148830825, 32'sd0.015336465347537936, 32'sd0.05439384089882402, 32'sd-0.02439692487562228, 32'sd0.03347664760182765, 32'sd0.07348179628972683, 32'sd-0.02052587354079598, 32'sd-0.043217997149101156, 32'sd0.08660693012213033, 32'sd-0.03806912424948667, 32'sd0.008853357432971783, 32'sd-0.04325067974822726, 32'sd0.153269624650187, 32'sd0.1225712562643312, 32'sd-0.06812332397874371, 32'sd-0.09777564008103756, 32'sd-0.003710569176202863, 32'sd-0.043991847462914506, 32'sd0.026735106249201394, 32'sd0.06388290101444899, 32'sd0.06483118984564479, 32'sd-0.07180590023141571, 32'sd0.06495430782900972, 32'sd-0.029751936314267365, 32'sd0.034601100595730454, 32'sd0.04867804043158417, 32'sd0.035517733722256375, 32'sd0.007058740150033106, 32'sd-0.01230854530466385, 32'sd-0.044961574006375606, 32'sd-0.0009649336384494146, 32'sd0.056163044530512615, 32'sd-0.026843539205147364, 32'sd0.014267807518254533, 32'sd-0.02759875802512561, 32'sd-0.029549012451285012, 32'sd0.12232807955664729, 32'sd0.05339828330206907, 32'sd0.05486395209909811, 32'sd-0.026393723984941147, 32'sd-0.015899536338002652, 32'sd-0.04998903995173092, 32'sd-0.05255735066978271, 32'sd-0.041479337568294784, 32'sd-0.013106602069768733, 32'sd-0.006321651717849793, 32'sd-0.008356247258647663, 32'sd-0.058340817613204574, 32'sd0.08575705677121763, 32'sd0.03741685075726053, 32'sd-0.018614655546254882, 32'sd-0.05384171525086337, 32'sd0.03482064922790585, 32'sd0.01815457762384892, 32'sd-0.008485024042509157, 32'sd-0.04519417644896281, 32'sd0.03236008794621444, 32'sd0.02547590840097697, 32'sd0.003526214994872415, 32'sd0.005026800925224995, 32'sd0.035514539829704296, 32'sd-0.03596072757694881, 32'sd0.005896176821265064, 32'sd-0.09162972741402485, 32'sd-0.025657633805300926, 32'sd0.0497947784934599, 32'sd0.07939614855883229, 32'sd0.05023112015847193, 32'sd0.10229208883858404, 32'sd0.12628036061836137, 32'sd-0.027108102821263243, 32'sd-0.06321332469010135, 32'sd-0.02800883336891695, 32'sd0.0062421344489531376, 32'sd0.02785407760070589, 32'sd-0.0940040996150065, 32'sd0.07057564215604237, 32'sd0.051558324451332266, 32'sd-0.06153887270488033, 32'sd0.008288392601369923, 32'sd-0.0942553692275621, 32'sd0.011178159000835425, 32'sd0.10748649342933805, 32'sd0.09090198005065574, 32'sd0.07341187794139087, 32'sd0.019825579386333645, 32'sd0.04672163963147574, 32'sd-0.009786381196467844, 32'sd0.018234876890729838, 32'sd0.02347313848783905, 32'sd0.06519575923949547, 32'sd0.029471989879946658, 32'sd0.05160357871222244, 32'sd-0.0327482489223259, 32'sd-0.016591930296748037, 32'sd0.056295318283362095, 32'sd0.03495847572290543, 32'sd0.10033753251950872, 32'sd0.178048293708623, 32'sd-0.009247166897295147, 32'sd-0.051785662425174586, 32'sd-0.08635614045314023, 32'sd-0.00032293557223885894, 32'sd-0.06676410899486272, 32'sd-0.06064282137626739, 32'sd-0.0881001981810355, 32'sd-0.06168628155572242, 32'sd-0.08052798819515482, 32'sd-0.05615894159332503, 32'sd0.02216373630251297, 32'sd0.12312727092733486, 32'sd-0.04520825522506211, 32'sd0.09576619319302701, 32'sd-0.02410851946919704, 32'sd-0.023459902347105478, 32'sd-0.14795049210401437, 32'sd0.04429116802915695, 32'sd0.04633311668725986, 32'sd0.0025666522138192275, 32'sd0.10218632021087841, 32'sd0.00040717508214317954, 32'sd-0.0196405385263276, 32'sd-0.008631035058767365, 32'sd0.016478087658497946, 32'sd-0.007578120208033755, 32'sd0.02391640186436873, 32'sd0.11176789980970643, 32'sd-0.04201362121077849, 32'sd0.013341849928972164, 32'sd-0.03169184153509547, 32'sd-0.16132261776628712, 32'sd-0.053969137513220466, 32'sd-0.055878999901689014, 32'sd0.020679643870184023, 32'sd0.03517417204478283, 32'sd-0.03780344015768225, 32'sd0.01018171623432889, 32'sd-0.009912057943372634, 32'sd0.1188916814307142, 32'sd0.0649674338203929, 32'sd0.14859706510474144, 32'sd-0.09815066976903046, 32'sd-0.12094138888987578, 32'sd-0.054233619317541455, 32'sd-0.022917185099910035, 32'sd0.07782939547642936, 32'sd0.042042320974585295, 32'sd0.09913494875116247, 32'sd0.03141037518172129, 32'sd0.03962162186268716, 32'sd0.067941166008618, 32'sd0.051311363203203474, 32'sd0.026968889198068842, 32'sd-0.013961465588999779, 32'sd0.04660773334741982, 32'sd-0.07190976828170999, 32'sd-0.1255050977721374, 32'sd-0.14208154063733447, 32'sd-0.12739655820583942, 32'sd-0.025161349472856264, 32'sd-0.011265227231241065, 32'sd0.05917828846252453, 32'sd-0.09073307790038614, 32'sd0.036651151412460115, 32'sd0.047132672033666105, 32'sd0.16824287460854614, 32'sd0.209588083426967, 32'sd0.053602575485500924, 32'sd-0.024636459412325597, 32'sd-0.05451176167103469, 32'sd0.01665918673880054, 32'sd-0.011083805059454433, 32'sd-0.025539186879000746, 32'sd0.00629225297329379, 32'sd-0.0054095868335865644, 32'sd-0.022986171331744458, 32'sd-0.050880406575164655, 32'sd0.07415692431769967, 32'sd0.02448382605969555, 32'sd-0.013847938682793404, 32'sd-0.05535439434769383, 32'sd0.009642823265666053, 32'sd-0.07002721800355277, 32'sd-0.03500036698468971, 32'sd0.04914016102230101, 32'sd-0.04155182410389172, 32'sd-0.03826051498611326, 32'sd0.042409227708119945, 32'sd-0.04582438149516118, 32'sd0.16415492475325422, 32'sd0.15177215172305755, 32'sd0.11330283503320396, 32'sd0.09759295933839757, 32'sd0.16102213941207236, 32'sd0.05051870584635265, 32'sd-0.008072159661848386, 32'sd0.01289413345456395, 32'sd0.0341545747245124, 32'sd0.11320862703900779, 32'sd0.03456758334987557, 32'sd-0.03170571306918835, 32'sd0.0361367511065038, 32'sd0.05895263762980802, 32'sd0.10441207633723527, 32'sd-0.0854997956655314, 32'sd0.05905596418393938, 32'sd0.004329804196461364, 32'sd0.05038783601359426, 32'sd-0.0552062006124544, 32'sd-0.03800404105849155, 32'sd-0.12299220385079239, 32'sd0.03900745446682585, 32'sd-0.047875403091056264, 32'sd0.031946584103182844, 32'sd0.06814889872409507, 32'sd0.1471781191233388, 32'sd-7.645703928145675e-05, 32'sd0.19456996320069514, 32'sd0.052906357443848806, 32'sd0.007229461157975628, 32'sd0.06877584343131903, 32'sd0.04279512861351362, 32'sd-0.016131029421637817, 32'sd0.023811395709688925, 32'sd0.11739301786005835, 32'sd0.09675995915561642, 32'sd0.10143364501071196, 32'sd0.052609290804743906, 32'sd0.013608371097725433, 32'sd-0.06345616193328418, 32'sd-0.019918938745476768, 32'sd0.0037978269438019383, 32'sd0.07331325793588792, 32'sd0.09898652082136306, 32'sd0.011169577612420933, 32'sd-0.00031416182502090595, 32'sd-0.01708484452474883, 32'sd-0.26283254638792575, 32'sd-0.11400614650417226, 32'sd0.0031186412088919447, 32'sd0.05567550259502682, 32'sd0.00585588287867915, 32'sd0.02973314914942224, 32'sd0.010173122657918303, 32'sd0.1291707223066652, 32'sd0.08986516575852542, 32'sd0.05703665136143746, 32'sd0.0023399816977019167, 32'sd0.0803607623165927, 32'sd0.1274428732949785, 32'sd-0.057109075058271765, 32'sd0.042634424600728554, 32'sd-0.01251610281734707, 32'sd-0.06911882853649051, 32'sd0.018124658265996133, 32'sd-0.059570519669813776, 32'sd3.788061182168619e-122, 32'sd-0.013272692961700083, 32'sd-0.002030168491324841, 32'sd0.03983292976514528, 32'sd0.0855039169482871, 32'sd0.04220191077270811, 32'sd-0.029284656376958533, 32'sd-0.14301471536242719, 32'sd-0.13989028464464406, 32'sd-0.27792288408320437, 32'sd-0.1497557799429238, 32'sd0.15622971163824256, 32'sd0.1415268995900721, 32'sd0.03026879780276285, 32'sd0.04662960810559801, 32'sd0.09421552831632024, 32'sd0.06630523804840147, 32'sd-0.036356426265746304, 32'sd-0.030984165741081763, 32'sd0.10785419158877516, 32'sd0.037102166740808525, 32'sd0.04638915838318394, 32'sd0.11386896058485363, 32'sd0.024033742337854033, 32'sd0.012443636310684963, 32'sd0.06569331111664473, 32'sd0.14055966375502976, 32'sd0.11698035228956595, 32'sd-0.029196428648312404, 32'sd0.029835050166905425, 32'sd-0.06598142182502817, 32'sd0.034360789894824995, 32'sd-0.0823293573727161, 32'sd-0.030580573030405, 32'sd-0.04232950385457567, 32'sd-0.13884389345534803, 32'sd-0.20906268194585093, 32'sd-0.1461547320471339, 32'sd-0.03599234008338555, 32'sd0.13037579255014572, 32'sd0.16084597677426668, 32'sd0.13417399675156597, 32'sd0.03122056216667076, 32'sd-0.003105952830877577, 32'sd-0.048881557025298034, 32'sd-0.0070457815226130805, 32'sd-0.05083803494453259, 32'sd-0.04446264145461484, 32'sd0.03240110425896578, 32'sd0.08406640893442908, 32'sd-0.0008170200100534254, 32'sd-0.07558805044520593, 32'sd-0.015135394996066562, 32'sd-0.061845652072794625, 32'sd0.07658804413010621, 32'sd0.10003369583021748, 32'sd-0.012707253767565796, 32'sd0.059635114678902305, 32'sd0.008576243427251783, 32'sd-0.02190505060278061, 32'sd-0.11913525119180243, 32'sd-0.08763080019519635, 32'sd-0.21847056282553215, 32'sd-0.16256252712168942, 32'sd-0.15930553697719962, 32'sd0.080036907493302, 32'sd0.2561494011810254, 32'sd0.09684402508976561, 32'sd0.025465356361188945, 32'sd0.013373897640388864, 32'sd-0.04267237325646952, 32'sd-0.014335069891282899, 32'sd-0.004247035242122709, 32'sd-0.12345519003561964, 32'sd-0.11281728894116358, 32'sd-0.055288367954703696, 32'sd-0.10637026854999995, 32'sd0.0031046687744216575, 32'sd-0.13181030422847112, 32'sd-0.1753411137225778, 32'sd-0.010095992713012049, 32'sd-0.07799864169778738, 32'sd0.04184657882758699, 32'sd0.09669565660171967, 32'sd-5.190121040873655e-126, 32'sd0.025338399030416757, 32'sd0.06006844275866861, 32'sd-0.05226697806086315, 32'sd-0.14351711897572508, 32'sd-0.06353608515145757, 32'sd-0.16212441102288158, 32'sd-0.1496934495495052, 32'sd0.0364202248228993, 32'sd0.045324097548750435, 32'sd0.21475123620565076, 32'sd0.14995131263745817, 32'sd0.0025892516136188813, 32'sd-0.05768162483695361, 32'sd-0.0008575409915156672, 32'sd-0.04697088804932632, 32'sd-0.07296026656436304, 32'sd-0.16178367923351997, 32'sd-0.05304297136094979, 32'sd-0.11853730925514026, 32'sd-0.14124235073590918, 32'sd-0.05270687901972784, 32'sd-0.08441753179370397, 32'sd-0.1410153557911142, 32'sd0.0747356699264056, 32'sd0.03496040064806836, 32'sd-0.04813884270815047, 32'sd-0.00407350734972006, 32'sd0.015528707550645159, 32'sd-0.03774034239684382, 32'sd-0.10472302487317019, 32'sd0.04381369704829911, 32'sd-0.04313234738425808, 32'sd-0.13152538862679417, 32'sd-0.1869378501354205, 32'sd-0.22661929940667394, 32'sd-0.004286575802560995, 32'sd0.028483808371741876, 32'sd0.04924100855658302, 32'sd0.0635907884283013, 32'sd0.08869948369986727, 32'sd0.07074922597265484, 32'sd-0.10672292611252429, 32'sd-0.1259805531892049, 32'sd-0.05945551697245658, 32'sd-0.14865136408668705, 32'sd-0.18484863886725703, 32'sd-0.09851231511056202, 32'sd-0.08689283363030105, 32'sd-0.11735588120741827, 32'sd-0.10902620236776484, 32'sd-0.08009629529980936, 32'sd0.08569059177528321, 32'sd-0.10680502348864905, 32'sd-0.07854154646513126, 32'sd-0.0388722063588, 32'sd-0.03090150916608771, 32'sd-0.02669833613939058, 32'sd0.01744583781423786, 32'sd-0.05786538555636111, 32'sd-0.10049044319662602, 32'sd-0.14801022532956634, 32'sd-0.1663742969102224, 32'sd-0.09976273466454412, 32'sd-0.12738961259721698, 32'sd-0.010937178579709675, 32'sd-0.016738072011813678, 32'sd0.06523892507131436, 32'sd0.24173887153021942, 32'sd0.22486775808708395, 32'sd0.05531703255102936, 32'sd-0.027044546436862164, 32'sd-0.10582237446501722, 32'sd-0.13391187429593487, 32'sd-0.12809858686654302, 32'sd-0.10610392910130255, 32'sd-0.0710613869881648, 32'sd-0.0151137107507002, 32'sd-0.016938793479881774, 32'sd0.036305117231332534, 32'sd-0.005597847149141926, 32'sd0.013395172007255927, 32'sd0.050003724457355084, 32'sd0.02306477238525109, 32'sd-2.8856111386590087e-118, 32'sd-0.006290668772678584, 32'sd0.0028942541402350143, 32'sd-0.11245453952084407, 32'sd0.04371345772235889, 32'sd-0.1064573646238209, 32'sd-0.10809337641727172, 32'sd-0.04130054926611075, 32'sd-0.04002692516312351, 32'sd-0.025611322765485698, 32'sd-0.10071385696142661, 32'sd0.017346239186123, 32'sd0.2064484995778113, 32'sd0.2832553386800496, 32'sd0.07872854026040625, 32'sd0.01686296927673428, 32'sd-0.06977984378646251, 32'sd-0.12288904385536269, 32'sd-0.10875765001332437, 32'sd-0.20597814093811412, 32'sd-0.10694182415000406, 32'sd0.05892825577502276, 32'sd0.0375335884845136, 32'sd0.02776535718745787, 32'sd-0.031265049520188146, 32'sd-0.07536715358502241, 32'sd-0.024397761522185108, 32'sd-5.074742310279872e-126, 32'sd4.975729926257557e-122, 32'sd2.543129513744851e-122, 32'sd0.051483137152896874, 32'sd0.029889249177197895, 32'sd0.07386460299092311, 32'sd-0.02846912703517154, 32'sd-0.06066277391790461, 32'sd-0.024933572478779437, 32'sd-0.07626594712884333, 32'sd-0.09158907532708016, 32'sd0.03212495355113316, 32'sd0.02941463131452683, 32'sd0.06020100526890884, 32'sd0.027700839803874912, 32'sd0.06388017988877653, 32'sd0.19154058707039964, 32'sd0.14652232008951868, 32'sd-0.0345095645691636, 32'sd-0.09608790959963702, 32'sd0.044180120961063545, 32'sd-0.0016104327881990878, 32'sd-0.017080159825853432, 32'sd0.06001669052374031, 32'sd0.04849189254388889, 32'sd-0.11661829817021539, 32'sd-0.06362052533677318, 32'sd-0.028597522515119628, 32'sd8.83037574888375e-119, 32'sd6.892296715116216e-126, 32'sd-1.8505304056139444e-124, 32'sd-0.03141328151861367, 32'sd-0.03942931382858348, 32'sd-0.1056281739792676, 32'sd-0.12600682411959485, 32'sd-0.029625185668487885, 32'sd-0.02922516859869248, 32'sd0.016519518176253793, 32'sd0.07377373183278539, 32'sd0.027055659137940787, 32'sd0.0011071914647239206, 32'sd-0.016761064748002378, 32'sd-0.05076615995564639, 32'sd0.13822459811401305, 32'sd0.039226567587717, 32'sd0.10875655496938097, 32'sd-0.07692387391722488, 32'sd0.019991629590663616, 32'sd-0.05282560547237352, 32'sd-0.043756364638926265, 32'sd-0.13258977803299515, 32'sd-0.07058571939869299, 32'sd0.013628869817905764, 32'sd0.03934338374540712, 32'sd0.02030155011707172, 32'sd-0.03373575201646809, 32'sd-2.8071456842339226e-119, 32'sd-2.529659600241268e-118, 32'sd3.2219845253278536e-122, 32'sd2.0335476628903614e-126, 32'sd0.027578679036532817, 32'sd0.035060528849212944, 32'sd0.04499033114068926, 32'sd-0.030473457345680507, 32'sd0.006888772363461276, 32'sd-0.10043915650107782, 32'sd0.05181623922744935, 32'sd0.037820937516490113, 32'sd-0.06386894099333087, 32'sd-0.06088818926864873, 32'sd0.08316227765997614, 32'sd0.06637811790282831, 32'sd0.02043462303514434, 32'sd0.03014201174951393, 32'sd0.03895003050070339, 32'sd0.02843532497075155, 32'sd-0.023035640015681386, 32'sd0.03218085881746865, 32'sd0.00013842694411607176, 32'sd-0.034131885386066596, 32'sd0.037928311267532974, 32'sd0.055778078193592595, 32'sd0.023784082097445133, 32'sd-7.209704007528278e-116, 32'sd-3.294341443185005e-121, 32'sd1.0629749948735199e-117, 32'sd5.913972254531722e-119, 32'sd-4.1521553995218526e-122, 32'sd-9.505450230741546e-123, 32'sd0.022731968663795597, 32'sd-0.0521606092604153, 32'sd-0.01605035629169006, 32'sd0.06801967616906968, 32'sd-0.016657164321589504, 32'sd0.000864541920034482, 32'sd0.0259093775084212, 32'sd0.047626980218567525, 32'sd-0.04722964125511902, 32'sd-0.022545012576452413, 32'sd0.007346965645988375, 32'sd-0.048251266286500644, 32'sd-0.010685464434821325, 32'sd0.12170293905194396, 32'sd0.08081911757209694, 32'sd-0.03297359293374846, 32'sd0.0001302841429348301, 32'sd-0.04027325700702636, 32'sd-0.1063929690317608, 32'sd0.021175303703128458, 32'sd3.543980962489353e-124, 32'sd2.1636121710504068e-124, 32'sd-2.8086046805546996e-119, 32'sd-5.241390394816233e-119},
        '{32'sd4.6433754615646315e-123, 32'sd-1.1340327730737704e-116, 32'sd4.702665365467718e-124, 32'sd-1.0070608969445509e-120, 32'sd3.606690184383097e-120, 32'sd-7.459771966869434e-119, 32'sd-6.223033608865225e-126, 32'sd2.836163061178848e-128, 32'sd5.056434692567939e-115, 32'sd-2.1866606636417408e-122, 32'sd2.4735159183696384e-125, 32'sd-9.14174340745035e-118, 32'sd0.012097782738146165, 32'sd-0.058474521883702085, 32'sd0.0018840450918207804, 32'sd-0.009371343201637933, 32'sd4.15259922924705e-125, 32'sd-1.3338887374491557e-122, 32'sd8.315533065205253e-124, 32'sd2.584234542706565e-121, 32'sd-2.569240638797327e-122, 32'sd-9.596106258401144e-123, 32'sd-3.133375098941123e-114, 32'sd-6.951804217669219e-124, 32'sd-1.0144903317865415e-119, 32'sd-1.9096433171473773e-127, 32'sd-3.8946873450821643e-119, 32'sd3.16968372353518e-121, 32'sd3.289058398152577e-120, 32'sd2.0425650185162766e-123, 32'sd1.7665350961913292e-124, 32'sd1.0725362086198634e-117, 32'sd-0.0175619250550619, 32'sd-0.03357724596726092, 32'sd0.039446402542039544, 32'sd-0.04217765296133062, 32'sd-0.03806624732854416, 32'sd0.04463888914705489, 32'sd0.0015732414101534973, 32'sd-0.07353475351583831, 32'sd-0.10592965263012018, 32'sd-0.12053899951667905, 32'sd-0.09508861695992457, 32'sd0.02020260666139985, 32'sd0.05962994369579021, 32'sd0.017849277079482195, 32'sd0.09836771699846739, 32'sd0.02705623247915918, 32'sd-0.06641455842061723, 32'sd-0.03658730559944723, 32'sd-0.01780044979211872, 32'sd0.06190181686589166, 32'sd-4.920605503044737e-123, 32'sd-4.4133799287938067e-128, 32'sd1.8002078461146824e-123, 32'sd6.28107934379999e-117, 32'sd1.700555769729873e-121, 32'sd1.108450819626654e-121, 32'sd-0.05191364713438205, 32'sd0.02452450479971923, 32'sd-0.05078258025449789, 32'sd-0.05442857710897695, 32'sd0.022090944138951796, 32'sd-0.07601385917273155, 32'sd0.06196824003735346, 32'sd0.1219469516147499, 32'sd-0.03043628478315825, 32'sd0.12159334816254652, 32'sd0.014614623955810143, 32'sd0.07207105953655457, 32'sd0.10360850595248627, 32'sd0.14357110612076224, 32'sd-0.01569284499160827, 32'sd0.0767442772138019, 32'sd0.013888182224026734, 32'sd0.056555531961734885, 32'sd0.07097528599140203, 32'sd0.11946112420742869, 32'sd0.022184051941586826, 32'sd-0.009224115845233166, 32'sd-0.04582506371991865, 32'sd-0.06423302945321391, 32'sd-8.896394226918965e-127, 32'sd1.0430145703877987e-124, 32'sd6.375243469471148e-122, 32'sd3.860770168510245e-124, 32'sd-0.03720811327289867, 32'sd0.03294386837475674, 32'sd-0.003919753183209947, 32'sd0.033553859944756036, 32'sd0.007644523375618836, 32'sd-0.08472702467134172, 32'sd0.07953517444353836, 32'sd-0.05127243714068126, 32'sd0.054276442869266896, 32'sd0.10600311127430502, 32'sd0.0968388744165247, 32'sd0.08023578578242598, 32'sd-0.022585678718748177, 32'sd0.04660880818240071, 32'sd-0.01645227286974095, 32'sd-0.02501556996622075, 32'sd0.08338108245850698, 32'sd-0.009182650903060781, 32'sd0.02564294171844547, 32'sd-0.12252106463688942, 32'sd-0.16380037057329416, 32'sd0.03133199361074385, 32'sd0.047694935538299406, 32'sd0.006506224644227748, 32'sd-0.05927995316589588, 32'sd4.763824875003954e-123, 32'sd1.0745384236515145e-124, 32'sd0.07464956560316867, 32'sd-0.047517424520154374, 32'sd0.009466481133640962, 32'sd0.021287846065386952, 32'sd-0.11214082148307782, 32'sd-0.09257445858540776, 32'sd-0.018919875318967, 32'sd0.11926820616168125, 32'sd0.03243638955598886, 32'sd0.08884404568688731, 32'sd0.0593553963743456, 32'sd0.08570698637065945, 32'sd0.13402998551598824, 32'sd0.07048596559925374, 32'sd0.02983232335858595, 32'sd0.1770759994127599, 32'sd-0.023491097174411918, 32'sd-0.012368446811710777, 32'sd0.021433763186762905, 32'sd-0.05993694714948575, 32'sd0.0095834106708642, 32'sd-0.05416023065732105, 32'sd-0.01720584704075071, 32'sd-0.011472799509346624, 32'sd-0.1373499757059419, 32'sd0.03808657821712927, 32'sd-0.023077531345802756, 32'sd3.610969214889359e-116, 32'sd-0.04264686103630654, 32'sd-0.028747401516012735, 32'sd-0.06556141956519324, 32'sd-0.07530720567934203, 32'sd-0.0955482333238644, 32'sd0.017371676670797316, 32'sd0.07118009985911775, 32'sd0.05039349433482907, 32'sd0.04466874160620324, 32'sd0.08526258284617247, 32'sd0.048437148878532024, 32'sd0.00028800100588608797, 32'sd0.1126783161397757, 32'sd0.02333260299482112, 32'sd-0.00862255026511698, 32'sd0.08041003545869325, 32'sd-0.05883929154254494, 32'sd-0.04021978503280515, 32'sd0.06569063877702898, 32'sd-0.02434831281408969, 32'sd-0.0800116662711733, 32'sd0.0039696813034683, 32'sd0.0657344059214463, 32'sd-0.054478775292170795, 32'sd-0.08830557881003517, 32'sd-0.00459267225436546, 32'sd-0.05845753053075106, 32'sd-1.5407087014101113e-117, 32'sd-0.05931497909324912, 32'sd0.047636292974150486, 32'sd0.06904200338388247, 32'sd0.0712026024237135, 32'sd0.04754958836389751, 32'sd-0.01425747572661854, 32'sd0.026489825186169734, 32'sd-0.04903558879180322, 32'sd0.08805334536124027, 32'sd0.1327707117966137, 32'sd-0.03377293610751775, 32'sd-0.012432713841901111, 32'sd0.02653747123165877, 32'sd-0.09959330111586524, 32'sd0.03504619262366983, 32'sd-0.11106504815858774, 32'sd-0.012362138250413903, 32'sd0.02049698301135507, 32'sd-0.05024671302147548, 32'sd0.0029307804103398272, 32'sd0.06465177218982034, 32'sd0.020433062028813294, 32'sd-0.04668378529720749, 32'sd-0.06812508803837593, 32'sd-0.07599547754195907, 32'sd-0.012338497097536993, 32'sd-0.058820508085579114, 32'sd-0.017181462521880724, 32'sd-0.015103382600844322, 32'sd-0.027082202507635406, 32'sd0.14129461920055547, 32'sd0.11358880923538169, 32'sd-0.06062666060962684, 32'sd0.07016027142887032, 32'sd0.11769211158251022, 32'sd0.04653993649361376, 32'sd-0.019261044232605194, 32'sd0.12887867589410984, 32'sd-0.04451952709077416, 32'sd-0.032108596608861145, 32'sd-0.1059854758956593, 32'sd-0.059222905415128764, 32'sd-0.1326878974778584, 32'sd0.00245730975202251, 32'sd0.019858016367710816, 32'sd-0.08022038939200332, 32'sd-0.062096206813428485, 32'sd-0.056409098987394594, 32'sd-0.060180664442133075, 32'sd-0.039239252735694875, 32'sd-0.08000289769387588, 32'sd-0.08346486363910698, 32'sd0.011858531644537023, 32'sd0.015237150633305383, 32'sd0.025378554674525954, 32'sd-0.0012573038397105623, 32'sd-0.02154433258045437, 32'sd-0.0889248393044998, 32'sd-0.08605297013524525, 32'sd-0.04945153322656812, 32'sd0.025385671165905205, 32'sd0.03883659273677517, 32'sd-0.008279954356369754, 32'sd-0.07244095670469891, 32'sd-0.01794106354866295, 32'sd-0.11453638563883287, 32'sd-0.08860927819501832, 32'sd-0.0168337953439172, 32'sd-0.03435884609403593, 32'sd-0.01906212342326245, 32'sd0.06508062549751151, 32'sd0.09002285629117575, 32'sd0.028691329907652784, 32'sd-0.1391557925101526, 32'sd-0.05079529314945538, 32'sd-0.011663996363839396, 32'sd0.017397297015360736, 32'sd0.08098656102399733, 32'sd-0.00602021389760993, 32'sd-0.06656544857214337, 32'sd-0.037666588855313446, 32'sd0.001383161595766032, 32'sd-0.014562582513639346, 32'sd-0.0434864121858838, 32'sd0.051054365500864306, 32'sd0.041542985376501244, 32'sd-0.05551486350403954, 32'sd0.03079911067722169, 32'sd0.03608085428110174, 32'sd-0.11323018380284934, 32'sd0.01153743518481986, 32'sd-0.12493519926755599, 32'sd-0.13111103277470967, 32'sd-0.14008759923117092, 32'sd-0.11025695566690824, 32'sd0.048208445861122384, 32'sd0.09276659310564049, 32'sd0.1299534506136483, 32'sd0.08327775514059482, 32'sd-0.012999475567727686, 32'sd0.009172629044853242, 32'sd-0.09451497278134974, 32'sd-0.03967732368784298, 32'sd0.1266718940934761, 32'sd-0.032966047349080894, 32'sd0.1397713618284829, 32'sd0.17062453699870242, 32'sd-0.0005648590003250115, 32'sd0.08218721677879987, 32'sd-0.11549786995285609, 32'sd-0.034278240188283, 32'sd0.006481037868984487, 32'sd-0.07274039853082039, 32'sd0.005607175462108145, 32'sd0.017660953203858083, 32'sd-0.07109395409274699, 32'sd-0.06772448069035866, 32'sd-0.058995299264463556, 32'sd-0.13106460521701085, 32'sd-0.08062747697831274, 32'sd0.016196543246484806, 32'sd0.0017802950524272061, 32'sd0.0475801759127249, 32'sd0.04007859000279864, 32'sd0.26444691193481396, 32'sd0.019055859861372475, 32'sd-0.06481404447283515, 32'sd-0.01220857126077142, 32'sd-0.04145527488103207, 32'sd0.03827084240398408, 32'sd-0.09726953938212278, 32'sd0.0882111854861416, 32'sd0.12463087374450287, 32'sd0.14868888564876145, 32'sd0.15640247864879736, 32'sd0.062362382059239156, 32'sd-0.02898712001696435, 32'sd-0.07361127289987013, 32'sd-0.031238737030340205, 32'sd-0.04209318044064888, 32'sd0.135308792673756, 32'sd-0.061149392778213546, 32'sd-0.07524410513319667, 32'sd-0.09446818202842966, 32'sd-0.1235229812142152, 32'sd-0.08242681240626068, 32'sd-0.05901793881218876, 32'sd0.02824523940409996, 32'sd0.08292160206998858, 32'sd0.18665275102021794, 32'sd0.13744321313693222, 32'sd0.20441192130128671, 32'sd0.016440895141554137, 32'sd-0.1430456973776424, 32'sd-0.1336486752943061, 32'sd-0.1938738529851878, 32'sd-0.1299177123175415, 32'sd0.004333649458080073, 32'sd0.05023511050251598, 32'sd0.10481971835025843, 32'sd-0.006016963618223263, 32'sd0.021055692560391925, 32'sd0.02824633726289697, 32'sd0.09944510913220103, 32'sd-0.0531017886913656, 32'sd-0.01454984528474227, 32'sd-0.0324297829046434, 32'sd-0.011136634660990425, 32'sd-0.036482679239509194, 32'sd-0.05223314186702635, 32'sd-0.012079013713824943, 32'sd-0.07858655308267179, 32'sd0.0034320302512611442, 32'sd-0.0035832191504722184, 32'sd0.22228827273088805, 32'sd0.17447648953415143, 32'sd0.24792806278504737, 32'sd0.2720227512828546, 32'sd0.1502735115227222, 32'sd0.08678901337062832, 32'sd-0.19577549702304378, 32'sd-0.14573595447239368, 32'sd-0.21695526157100872, 32'sd-0.003425207732684847, 32'sd-0.04685871410631576, 32'sd-0.08362050745168013, 32'sd-0.12820397838167988, 32'sd-0.1093214656607154, 32'sd-0.014918251307378848, 32'sd0.04765545363868992, 32'sd-0.026267893572586822, 32'sd-0.037637142881964174, 32'sd-0.0025761979219750637, 32'sd-0.054187900913212385, 32'sd-0.00809494465008196, 32'sd0.055553025247319456, 32'sd0.03177474114868432, 32'sd-0.08275368584300766, 32'sd-0.030423654086940425, 32'sd0.005162882557109174, 32'sd-0.1079456928194577, 32'sd0.018238535547461056, 32'sd0.20449986096819078, 32'sd0.30268327325832745, 32'sd0.279074360086884, 32'sd0.07566893295971425, 32'sd0.0003771543896726235, 32'sd-0.18255881912938204, 32'sd-0.22200578757126227, 32'sd-0.0826936145654714, 32'sd-0.17321022385676102, 32'sd-0.030556209448835445, 32'sd0.017776086901890448, 32'sd-0.14905975330811497, 32'sd-0.27124809796218124, 32'sd-0.04553040983387404, 32'sd-0.0570448929056887, 32'sd-0.0010388353075652809, 32'sd0.06232781916491182, 32'sd-0.03183400682438558, 32'sd0.0025627212460022793, 32'sd0.06625810515616379, 32'sd0.038233036591825725, 32'sd-0.04001292981601421, 32'sd-0.013112186843657078, 32'sd-0.07412394819752556, 32'sd-0.03290856372760838, 32'sd-0.044054488772046395, 32'sd0.04045556950356683, 32'sd-0.014906082541330454, 32'sd-0.0032609761244260824, 32'sd0.10841171448557736, 32'sd-0.04512863259514536, 32'sd-0.15630994726318714, 32'sd-0.23151667256132477, 32'sd-0.2463000243739733, 32'sd-0.12790590490658227, 32'sd-0.13512206977126923, 32'sd-0.08998551741592622, 32'sd-0.057866391990557646, 32'sd-0.05619097339069958, 32'sd-0.05632853339692022, 32'sd-0.18204125141747146, 32'sd-0.08067777647534113, 32'sd0.06227278180760741, 32'sd0.027096123312610305, 32'sd-0.010639495452773377, 32'sd0.024512938842204988, 32'sd0.07765199148008906, 32'sd0.05809371501695851, 32'sd0.11107871670674736, 32'sd-0.05341650314348836, 32'sd0.002706670185023084, 32'sd-0.05704816075176413, 32'sd0.02471488184423095, 32'sd-0.03791850931514885, 32'sd0.05959030091941185, 32'sd-0.09286392216473013, 32'sd0.07955010416946484, 32'sd0.019228670783633568, 32'sd-0.09895059672614184, 32'sd-0.2958323645092953, 32'sd-0.28783420544696536, 32'sd-0.35582651710768376, 32'sd-0.1329364467841359, 32'sd-0.11205077655601722, 32'sd-0.09507942062713891, 32'sd0.034933915517359894, 32'sd-0.10686592211453444, 32'sd-0.10574949890569185, 32'sd-0.15695055939287866, 32'sd-0.02977943897910146, 32'sd0.007146025830371193, 32'sd0.05940804405431967, 32'sd-0.0738922688707908, 32'sd0.05171824072832578, 32'sd0.030867465435901763, 32'sd0.029657308350459783, 32'sd-0.07229702796795619, 32'sd-0.0232608776681362, 32'sd0.0746162136021987, 32'sd-0.014495533537495069, 32'sd0.050765762473017575, 32'sd-0.09344787728915285, 32'sd-0.06050321566599803, 32'sd-0.11646634369205981, 32'sd-0.0873358408002996, 32'sd-0.11716646912234893, 32'sd-0.09956169907505492, 32'sd-0.16300707277087972, 32'sd-0.20336316200840707, 32'sd-0.25216478200877096, 32'sd-0.22945274383487907, 32'sd-0.04109258462245113, 32'sd-0.025201138105358126, 32'sd0.0578644146054298, 32'sd-0.1609192470592226, 32'sd-0.1500523333070679, 32'sd-0.17210871480542494, 32'sd-0.05560501413875561, 32'sd0.02892245457259513, 32'sd-0.014492156411542258, 32'sd0.05479226885486707, 32'sd0.11735917611344229, 32'sd0.030557965587010596, 32'sd-0.04407993478533036, 32'sd-0.013991254204450469, 32'sd1.61535049853804e-129, 32'sd-0.03009057051110312, 32'sd0.1050072157818738, 32'sd-0.024140514904995882, 32'sd0.09781110488993382, 32'sd0.05326115738490582, 32'sd-0.12617617010311624, 32'sd-0.0034739522529062144, 32'sd-0.1398189461861402, 32'sd-0.11395422992309902, 32'sd-0.1428383903334312, 32'sd-0.24280482051660748, 32'sd-0.1252665737025551, 32'sd-0.061304868819224013, 32'sd-0.14204388648722285, 32'sd-0.07781897694384644, 32'sd0.11695181202562954, 32'sd-0.07959926711490706, 32'sd-0.10396478375814282, 32'sd-0.054817801113968466, 32'sd0.03268838816325455, 32'sd-0.0013496355308831073, 32'sd0.02457205627395095, 32'sd0.10916652360632578, 32'sd0.13958705667514254, 32'sd0.048005316894328895, 32'sd-0.0553190845667017, 32'sd0.05250937692309014, 32'sd-0.023786881891832617, 32'sd0.016915942058948898, 32'sd-0.03233482816649286, 32'sd0.031075101784046065, 32'sd-0.007805050000926127, 32'sd0.1047960593067653, 32'sd0.02209975428127143, 32'sd0.002915276264379503, 32'sd-0.04309780314440171, 32'sd0.015644771264322652, 32'sd-0.07088319092195046, 32'sd-0.19226479705340951, 32'sd-0.07135773001048672, 32'sd-0.016451597579864, 32'sd-0.20855850435335627, 32'sd-0.12143937479357068, 32'sd0.09438752260581998, 32'sd-0.0783091948769262, 32'sd0.008732883563169928, 32'sd-0.04487106011343875, 32'sd-0.043780685947693306, 32'sd0.08135453589726103, 32'sd0.023326187960820876, 32'sd0.10039563290276153, 32'sd0.01707074167475144, 32'sd-0.16166755529785123, 32'sd-0.003252094732899301, 32'sd-0.058752116158208245, 32'sd-0.04192221331415031, 32'sd-0.04544529593816779, 32'sd-0.0010343858004305548, 32'sd0.02755542879922351, 32'sd-0.04140634239232949, 32'sd0.08464896685785116, 32'sd0.06643033306240943, 32'sd0.10956931868826572, 32'sd0.0067593687143529734, 32'sd0.009027295017593475, 32'sd-0.06042245931909018, 32'sd0.04949521053006598, 32'sd-0.09900367623923853, 32'sd0.008712799902405822, 32'sd0.019121394821764538, 32'sd-0.00016039372646943514, 32'sd0.027552614985238526, 32'sd-0.01801533613077797, 32'sd0.06678767911715605, 32'sd0.04660917807783433, 32'sd0.07400465069427652, 32'sd0.028762088479719686, 32'sd-0.02849002176996354, 32'sd0.0009583459498481519, 32'sd0.02379530810732014, 32'sd-0.11610891685694377, 32'sd0.006942399043885257, 32'sd-0.03492658765825012, 32'sd-6.743107949951018e-124, 32'sd0.0217040176325013, 32'sd-0.09249872412765649, 32'sd-0.005373446191050569, 32'sd0.049132595330857655, 32'sd0.0209480636452975, 32'sd0.08086277401555349, 32'sd0.1468484094743887, 32'sd0.10555233715695053, 32'sd0.09648209286927055, 32'sd0.10161310880671376, 32'sd0.10272135679999236, 32'sd-0.08017502096366966, 32'sd-0.017690252373771462, 32'sd0.0732321803883528, 32'sd0.1086879174371804, 32'sd0.10620652961544014, 32'sd0.05155330157575591, 32'sd0.08772551303692602, 32'sd0.03417289478673393, 32'sd0.07389402110849086, 32'sd0.09543312622070338, 32'sd-0.007003175995682612, 32'sd0.010312886856925578, 32'sd0.005818940592986555, 32'sd-0.009017916795838453, 32'sd0.019810984519811378, 32'sd-0.028620549855141314, 32'sd-0.033654535389170376, 32'sd-0.02023808792408753, 32'sd-0.006265238972522462, 32'sd-0.02277157634008396, 32'sd0.04714827636778055, 32'sd-0.044138925610793925, 32'sd-0.009732346042257119, 32'sd0.057438226547842634, 32'sd0.05832106194888012, 32'sd-0.02696588020560685, 32'sd0.06716207189728682, 32'sd0.13066658727675337, 32'sd-0.0848836585001681, 32'sd0.008060937552316313, 32'sd0.17888563645823133, 32'sd0.03429075911779032, 32'sd0.13200894839125216, 32'sd0.13924685491025265, 32'sd0.0887689968771226, 32'sd0.056153835990220176, 32'sd-0.06148948733790911, 32'sd-0.0824510229835014, 32'sd0.03791862022838161, 32'sd0.062481113441418996, 32'sd-0.10469100625195776, 32'sd0.04339608751576746, 32'sd-0.060391364806888725, 32'sd0.04231392744969116, 32'sd0.012875993714740656, 32'sd-0.04746753031356404, 32'sd-0.03242798425244649, 32'sd-0.0013941498619446724, 32'sd-0.030453146852460762, 32'sd0.052769335424768214, 32'sd0.015528593039943278, 32'sd-0.033999032872977085, 32'sd0.029699838537242267, 32'sd-0.019289558987095484, 32'sd0.06123372233902092, 32'sd0.05858877637372539, 32'sd0.1304439611721468, 32'sd0.009127757953527018, 32'sd0.005350985610262782, 32'sd0.11489636907888574, 32'sd-0.04084775600013167, 32'sd0.07751824130508794, 32'sd0.023956078473650288, 32'sd0.015074978995368507, 32'sd0.03368897064797143, 32'sd-0.01982596157217678, 32'sd0.11882805229518764, 32'sd0.07602945153845685, 32'sd0.000964171665959192, 32'sd-0.06529622048728384, 32'sd0.002641149996940608, 32'sd0.039714945762253026, 32'sd-1.963218722075315e-127, 32'sd-0.030980332670035464, 32'sd0.00959317951778368, 32'sd-0.1364001458146386, 32'sd-0.0018388312784245763, 32'sd0.005574199371166847, 32'sd0.02066004415146606, 32'sd0.07655015610445501, 32'sd-0.01905463403404196, 32'sd0.06400742531102842, 32'sd0.06267759112453754, 32'sd0.11327197666319815, 32'sd0.05021949987191368, 32'sd0.03821058470695453, 32'sd-0.11115870130505638, 32'sd0.16909155806939802, 32'sd0.09191164043387111, 32'sd0.0021706427909681456, 32'sd0.012504913746944004, 32'sd-0.15053384656059987, 32'sd-0.03888910777117049, 32'sd-0.04599182061754768, 32'sd-0.09038663112791268, 32'sd0.09101599879998865, 32'sd0.08099250678562848, 32'sd-0.010298685617619529, 32'sd-0.02090080273962191, 32'sd-8.90028259181015e-127, 32'sd-3.1877281951914905e-121, 32'sd3.443478334483743e-125, 32'sd-0.001766035629957014, 32'sd0.0026509503763404675, 32'sd0.04955941453800267, 32'sd-0.012503852979275299, 32'sd-0.01450261905198768, 32'sd0.15300783506281665, 32'sd0.0402571044645047, 32'sd0.12112728399883495, 32'sd0.011419027124802378, 32'sd0.02993787648276551, 32'sd-0.0013090161886908811, 32'sd-0.0794660546629054, 32'sd0.02762653036875541, 32'sd0.11654661645304573, 32'sd-0.016204818752572594, 32'sd0.05073916761722424, 32'sd0.05375513586559266, 32'sd-0.044066881651615965, 32'sd-0.15851827897055362, 32'sd-0.0010151878029624772, 32'sd-0.020464837453906013, 32'sd0.008900941592871137, 32'sd0.016668919196533575, 32'sd-0.07744143884573912, 32'sd0.06712933103683646, 32'sd3.518326522396298e-122, 32'sd-3.303430897821872e-116, 32'sd8.665589424756164e-127, 32'sd-0.012335443906054502, 32'sd-0.0009968186609033312, 32'sd-0.06656128273488847, 32'sd0.012082579659737335, 32'sd-0.04162784762346911, 32'sd0.05430372526356447, 32'sd0.021824942579636405, 32'sd0.16149119179562269, 32'sd0.03235391966866773, 32'sd0.12965076281303217, 32'sd0.15607084509175337, 32'sd0.08377440383295318, 32'sd0.05890445594577108, 32'sd0.09894145576641336, 32'sd0.011699188616891343, 32'sd0.021897304520581314, 32'sd0.04848608027027524, 32'sd0.13005556678364544, 32'sd0.0826814186440432, 32'sd0.09666108148376598, 32'sd0.025853044405833685, 32'sd0.037297418336240624, 32'sd0.07993352690896267, 32'sd-0.005331614556646714, 32'sd-0.011668578148331507, 32'sd-8.011795973398454e-119, 32'sd2.5163139218016685e-124, 32'sd-6.862349685012604e-126, 32'sd-8.257790238659523e-127, 32'sd0.015043317230611619, 32'sd0.029225384093435603, 32'sd-0.027088799724574564, 32'sd0.05423981076521139, 32'sd0.044184986301689516, 32'sd-0.016769351934427593, 32'sd-0.08767723348937355, 32'sd0.05969772094691986, 32'sd0.03523971099670504, 32'sd0.09550974772020064, 32'sd0.042640262083783645, 32'sd0.01667405593195734, 32'sd0.09953107297440446, 32'sd0.13166537335616163, 32'sd0.07029578721561362, 32'sd0.018574031420021675, 32'sd0.08881226175200448, 32'sd0.017468672572418454, 32'sd0.032805992678387165, 32'sd0.04147844127775533, 32'sd0.035538331201242106, 32'sd-0.08773330898559467, 32'sd0.061283290571312536, 32'sd-6.715496729604391e-126, 32'sd4.8317059793884747e-123, 32'sd1.2170305558200285e-122, 32'sd-2.1075214623287694e-127, 32'sd-3.4261131870716813e-119, 32'sd1.3959680484672484e-123, 32'sd-0.017519176436139382, 32'sd-0.060896051877682406, 32'sd-0.022491501440730928, 32'sd-0.014767385885499565, 32'sd0.1082513418733462, 32'sd0.050210431361368685, 32'sd0.08364983703339099, 32'sd-0.06900234731931534, 32'sd0.05784155994119362, 32'sd0.034949812424660165, 32'sd-0.04254161716730026, 32'sd-0.0889845694128342, 32'sd-0.06793246994042584, 32'sd-0.008748217818807453, 32'sd0.03254012851254224, 32'sd0.0717403751973155, 32'sd0.0017141580640380374, 32'sd0.026463800163805232, 32'sd0.06321143012397197, 32'sd0.015468464235939833, 32'sd1.0896363904998383e-121, 32'sd-1.0561563496998545e-125, 32'sd-2.2653244652259684e-117, 32'sd2.1668068843474866e-127},
        '{32'sd-3.4160139336317256e-123, 32'sd8.241187566054829e-116, 32'sd-3.2899248310168434e-120, 32'sd-1.1684924359817252e-122, 32'sd2.516637603215059e-124, 32'sd-1.9664454910046562e-126, 32'sd3.7417554536227966e-125, 32'sd8.257291358039096e-127, 32'sd6.0736887734007664e-124, 32'sd-3.798652308399228e-122, 32'sd-1.6244166758567993e-115, 32'sd-2.8086469397145224e-121, 32'sd0.06098301818474711, 32'sd-0.0020941630750751367, 32'sd0.015221612116688519, 32'sd-0.0032328470018804876, 32'sd7.892712715119729e-126, 32'sd-1.2022229058792653e-125, 32'sd7.561857551613663e-117, 32'sd-5.044454032606161e-125, 32'sd4.6955828571180315e-124, 32'sd7.169724359805494e-122, 32'sd3.196422352732617e-118, 32'sd-2.56169447780046e-119, 32'sd-4.560125939879074e-126, 32'sd3.6358412714271306e-120, 32'sd-2.9824639572077817e-118, 32'sd-4.8351435017675895e-123, 32'sd-3.316752340228695e-120, 32'sd-4.078703603715929e-117, 32'sd-2.9877053039697226e-114, 32'sd1.8590517932420283e-117, 32'sd0.03224338685845786, 32'sd0.017524057975016324, 32'sd-0.020016401073893453, 32'sd-0.04517002208122701, 32'sd-0.07886696356977946, 32'sd0.0048303471990400445, 32'sd0.02852559210896045, 32'sd0.10551652035064046, 32'sd0.019295911461637512, 32'sd0.01726432584792724, 32'sd0.024844309017651185, 32'sd0.05308709581582108, 32'sd-0.02153985397438602, 32'sd0.08847377291178006, 32'sd-0.00031180750073502104, 32'sd0.07964312163200711, 32'sd0.06394535080774628, 32'sd0.04963905169702799, 32'sd0.07341778765170162, 32'sd0.00596146587288047, 32'sd-1.3053783202086833e-117, 32'sd-9.589559731846737e-127, 32'sd-9.92085400337851e-121, 32'sd-7.198748735253824e-115, 32'sd4.472071985248526e-118, 32'sd-1.516428888310551e-124, 32'sd0.022644400569213238, 32'sd0.009264221027086798, 32'sd0.07966775456727156, 32'sd-0.02378948703639703, 32'sd0.03263950001040027, 32'sd-0.05563556069461101, 32'sd-0.024585037243191516, 32'sd-0.05457445946439486, 32'sd-0.028039394729933585, 32'sd0.02908440792211543, 32'sd0.037759014388782826, 32'sd0.17696444689611496, 32'sd0.03861197912118736, 32'sd0.11198860403108958, 32'sd0.02488025582867566, 32'sd0.10270805795352062, 32'sd-0.031669828323206084, 32'sd0.02417783718891811, 32'sd-0.005087627232454065, 32'sd0.05387313895184951, 32'sd0.08729839505246673, 32'sd0.05139567264857201, 32'sd0.043545399785356216, 32'sd0.0037900594450402405, 32'sd3.809876755080611e-119, 32'sd5.4278267814864224e-126, 32'sd1.142560033471374e-118, 32'sd1.159330584959432e-122, 32'sd-0.015924123027744496, 32'sd-0.0562687244492705, 32'sd0.06625482699109977, 32'sd0.0016670053459725746, 32'sd0.04364507711498262, 32'sd0.034315915942507734, 32'sd-0.11506426533052298, 32'sd0.024855397865395826, 32'sd-0.08722008181797777, 32'sd-0.07021059269269776, 32'sd0.12159290345178285, 32'sd0.03644132653736434, 32'sd0.11283657145568282, 32'sd0.0357783985347852, 32'sd-0.02838074379538829, 32'sd-0.006806937949886989, 32'sd-0.04766000405049621, 32'sd-0.17174199754323757, 32'sd-0.1310141751483285, 32'sd-0.10307942265726963, 32'sd-0.09540176808378592, 32'sd-0.15428415729669454, 32'sd-0.02381111582171977, 32'sd-0.05521658209961822, 32'sd0.016424432690239254, 32'sd-3.88071832617934e-120, 32'sd2.8142580484287393e-118, 32'sd-0.0007235919224366144, 32'sd0.0560851069611941, 32'sd0.02807489563275831, 32'sd-0.10516611180613628, 32'sd0.000817425862536579, 32'sd-0.0017890229282014494, 32'sd-0.10779051448465732, 32'sd-0.06887792393799819, 32'sd-0.10141902877949502, 32'sd-0.16496351229439016, 32'sd0.15820919588667942, 32'sd0.1019215422497976, 32'sd0.09368637761077304, 32'sd-0.07880006683588765, 32'sd0.09112473527882785, 32'sd-0.10063281280997875, 32'sd-0.012386661707241033, 32'sd-0.009454972598136619, 32'sd-0.0992098852370448, 32'sd-0.05300438573681819, 32'sd-0.021212160629315226, 32'sd0.03991888844043522, 32'sd0.011008407850239233, 32'sd0.00694229168463897, 32'sd-0.07113904876733344, 32'sd0.028486164871162886, 32'sd0.022320689199852438, 32'sd2.526177760547026e-124, 32'sd0.03412338770866647, 32'sd0.06016016755726778, 32'sd-0.03790484714532443, 32'sd-0.0692940268070815, 32'sd-0.0456675646784582, 32'sd-0.15392865006334128, 32'sd-0.15567197047246675, 32'sd-0.05444662382355934, 32'sd-0.02344391883277061, 32'sd0.03595734619368335, 32'sd0.12054744818880311, 32'sd0.10103382822964933, 32'sd0.04002313685823526, 32'sd0.10168865307525904, 32'sd0.08873214496980812, 32'sd-0.05203450328988815, 32'sd-0.14441629497868833, 32'sd0.008724847392315849, 32'sd-0.05468145581858837, 32'sd-0.13442010751689074, 32'sd0.0320964178938141, 32'sd0.052673424111139566, 32'sd-0.05167774714775191, 32'sd0.10434596659998807, 32'sd-0.07313035624830899, 32'sd0.048151377391995466, 32'sd-0.018112401747881954, 32'sd-3.235887582503892e-124, 32'sd-0.009773311549896144, 32'sd0.003205168193451202, 32'sd0.008097568561478244, 32'sd-0.03944651077491577, 32'sd-0.02571351821870178, 32'sd-0.2140043824072195, 32'sd-0.1347308962386554, 32'sd-0.04718955051273923, 32'sd-0.11098747438748015, 32'sd-0.13805088852768274, 32'sd0.07612320180401397, 32'sd-0.0061325683948948405, 32'sd0.15463912760228424, 32'sd0.07860728419088836, 32'sd-0.08468180234053568, 32'sd-0.1285627489456648, 32'sd-0.13993424189654025, 32'sd-0.004345516468900883, 32'sd0.004697169171469806, 32'sd-0.013723025257602604, 32'sd0.09620536348577148, 32'sd0.13350258406391302, 32'sd0.08028941262122662, 32'sd0.17093529162698193, 32'sd0.1330160611561773, 32'sd0.11833666936272759, 32'sd0.07984742314780283, 32'sd0.011050640644197992, 32'sd0.02922314136227665, 32'sd0.002738722809598351, 32'sd9.568981313306847e-06, 32'sd-0.0038220200700603384, 32'sd-0.005932783657066491, 32'sd-0.08996307415704874, 32'sd-0.06049630378392414, 32'sd-0.2562174428295603, 32'sd-0.2183704478641762, 32'sd-0.006367395332802584, 32'sd0.19290754398807494, 32'sd0.1263523594058977, 32'sd0.13362104563250296, 32'sd-0.10071922912710271, 32'sd-0.006155450752319085, 32'sd0.0613950940897793, 32'sd0.012893029761894532, 32'sd0.14967110941069106, 32'sd0.11693142828548234, 32'sd0.1385577691126925, 32'sd0.13156424895791544, 32'sd0.13240271584680316, 32'sd0.13025853149257002, 32'sd0.11752357028470169, 32'sd0.14289337859308954, 32'sd0.015286011457057293, 32'sd-0.030385822960876278, 32'sd0.04932998470838147, 32'sd-0.008787807701834538, 32'sd-0.09889722698990196, 32'sd0.021309297989454072, 32'sd-0.04889477318368131, 32'sd0.09001303228056393, 32'sd-0.06018291703625693, 32'sd-0.06764119687407563, 32'sd-0.26117353046207276, 32'sd-0.011675936864098494, 32'sd-0.018514075430505678, 32'sd0.14096986442830106, 32'sd0.1781870509132302, 32'sd0.019215614824483467, 32'sd0.014945810436661043, 32'sd0.07176824754329894, 32'sd-0.022899785324040703, 32'sd0.12868606306321775, 32'sd0.14348905147198762, 32'sd0.06039812433316144, 32'sd-0.03700303866760343, 32'sd0.05563979860372619, 32'sd0.06086523091538555, 32'sd-0.06348260339102685, 32'sd0.04395973880715427, 32'sd-0.07438220434155465, 32'sd-0.03355262166949599, 32'sd-0.05810163812223761, 32'sd0.10599148666666937, 32'sd-0.02836042150187336, 32'sd-0.040815934870178955, 32'sd-0.02571847262213709, 32'sd0.045886883074201065, 32'sd0.07553980333231285, 32'sd-0.0728886268511051, 32'sd-0.18746846222400543, 32'sd-0.17101725756349564, 32'sd0.050334109259593904, 32'sd-0.06013884237771934, 32'sd0.11641128595529605, 32'sd0.11603346133630245, 32'sd0.03429728623408329, 32'sd-0.14394673913225367, 32'sd-0.02806619274105247, 32'sd-0.007315749183628124, 32'sd-0.1537814583844752, 32'sd-0.056732309625633824, 32'sd-0.13755563399792267, 32'sd-0.08903905417122097, 32'sd-0.10586434257591677, 32'sd-0.04179571372396901, 32'sd-0.05219534562075282, 32'sd-0.07991655937263277, 32'sd-0.1278204417333233, 32'sd-0.04575683883992207, 32'sd0.024015137671847, 32'sd-0.011322635412845134, 32'sd0.052804079185742654, 32'sd0.004121578799497579, 32'sd-0.02773706130092268, 32'sd-0.04642542832044473, 32'sd0.07206468319824362, 32'sd0.01991087345881009, 32'sd-0.09644550366676528, 32'sd-0.19542634094205025, 32'sd-0.03254557426778538, 32'sd0.07527419166542912, 32'sd0.18821116884666386, 32'sd0.07156642216391894, 32'sd-0.028947667216323032, 32'sd-0.056002876920965824, 32'sd-0.1263312228905468, 32'sd-0.17984569104411982, 32'sd-0.09544996775704391, 32'sd-0.08977886859583392, 32'sd-0.17422178672411504, 32'sd-0.25151261854988277, 32'sd-0.07364415883472246, 32'sd-0.016001701544176232, 32'sd-0.08950223108587056, 32'sd-0.030487706646216268, 32'sd-0.01491689519722314, 32'sd-0.07002489381463822, 32'sd-0.07909424587677281, 32'sd0.01644309551911268, 32'sd-0.08614124826223347, 32'sd-0.08613126768567264, 32'sd-0.049199194389833126, 32'sd-0.011972501944068445, 32'sd0.0007910266277277341, 32'sd-0.051131531151168065, 32'sd-0.007446989644426685, 32'sd-0.18224551701087294, 32'sd-0.09001214847183647, 32'sd0.007970514456147366, 32'sd0.029959287652994347, 32'sd-0.008809205825016023, 32'sd-0.061181134558748435, 32'sd-0.0316482564367456, 32'sd-0.2515568724316653, 32'sd-0.0297811252661737, 32'sd-0.007285099495518447, 32'sd-0.07876835804534023, 32'sd-0.06645486846245365, 32'sd-0.16686201745219925, 32'sd-0.0036671930299121947, 32'sd0.046516009494251734, 32'sd0.07256742150069558, 32'sd0.11555415764638002, 32'sd-0.08901436571499231, 32'sd0.06273229580611034, 32'sd-0.0501387563417601, 32'sd0.04203818901960083, 32'sd-0.04740511789037619, 32'sd0.0487230369092433, 32'sd-0.09151281890865266, 32'sd0.018083351522783373, 32'sd0.012005314303958552, 32'sd0.0325692998748546, 32'sd-0.10274743036845514, 32'sd-0.039774645073760995, 32'sd0.002195957989323485, 32'sd-0.013797027213799242, 32'sd0.10484505256328781, 32'sd-0.04045533484215332, 32'sd-0.040398636445677476, 32'sd-0.035515698006424234, 32'sd-0.066260473121448, 32'sd-0.19012084980018634, 32'sd0.013705956107966252, 32'sd0.09209051871891735, 32'sd0.018411678616819815, 32'sd-0.11038367481280596, 32'sd-0.06738089101699805, 32'sd-0.0627427406148529, 32'sd0.06673899579171648, 32'sd0.0266049103889605, 32'sd0.08863103961885117, 32'sd0.09705836992238327, 32'sd0.034971879712971256, 32'sd0.0431031838567855, 32'sd-0.005916282915549, 32'sd-0.044793643030154144, 32'sd-0.03504375305286337, 32'sd0.04613377213445071, 32'sd0.12678290804990536, 32'sd-0.040688455489335085, 32'sd0.05152430441292732, 32'sd-0.09991354208585956, 32'sd-0.10145388976336846, 32'sd0.023115079107448745, 32'sd-0.06401183779980175, 32'sd-0.04634629570550142, 32'sd-0.07187804297763607, 32'sd0.03856700633090791, 32'sd-0.009567690243050141, 32'sd-0.08004221561422348, 32'sd-0.0826365157969779, 32'sd-0.05505529626018594, 32'sd0.09380070600297856, 32'sd0.06021295494602984, 32'sd0.024294173448036083, 32'sd0.010733061030719807, 32'sd0.04034322970021143, 32'sd-0.04317662734034837, 32'sd0.04709780619751056, 32'sd0.042447638437721424, 32'sd-0.049301999936290065, 32'sd0.03441900110333585, 32'sd0.0797596660929326, 32'sd0.0459844843024552, 32'sd-0.013132205947767636, 32'sd0.031286080410206765, 32'sd0.029221875338904486, 32'sd-0.05172230438353881, 32'sd0.08686772738188538, 32'sd-0.035942260003673385, 32'sd0.06003994427425539, 32'sd-0.009501931609283296, 32'sd-0.09723316317176146, 32'sd-0.06081413947415334, 32'sd-0.03745606173582031, 32'sd0.014126143549641304, 32'sd0.11800600833287012, 32'sd0.03930990188872538, 32'sd0.046336245572101996, 32'sd-0.017099709283588144, 32'sd-0.007967308286086659, 32'sd-0.026671429126543928, 32'sd0.035267916981438815, 32'sd0.11342264445762462, 32'sd0.0953418092278435, 32'sd-0.032447716207621206, 32'sd0.09017589276631079, 32'sd0.012465827101674765, 32'sd0.029951232036813474, 32'sd0.11150896036144634, 32'sd-0.06662088687120749, 32'sd-0.08988741082914632, 32'sd0.03994927896500148, 32'sd-0.021730404904436722, 32'sd0.09299799338770566, 32'sd-0.09088191254640983, 32'sd-0.10282773614868815, 32'sd-0.08121844122713512, 32'sd0.029260458889585686, 32'sd0.07610410248426594, 32'sd0.05095349273855672, 32'sd0.10403551413160589, 32'sd-0.10004480238113726, 32'sd-0.07044591462437295, 32'sd0.0727426135246189, 32'sd-0.05373702978223123, 32'sd0.09049597879372011, 32'sd0.0333274984629985, 32'sd-0.1546158715885849, 32'sd-0.047727748047091074, 32'sd0.05550182147754711, 32'sd0.13976692942836078, 32'sd0.04161313319770833, 32'sd0.037739455558899605, 32'sd0.024301610695654927, 32'sd-0.006706843421135157, 32'sd0.024534082357079035, 32'sd0.017836114033546898, 32'sd-0.016714764936347448, 32'sd0.06545416270805618, 32'sd0.040828717059837656, 32'sd0.06235735756069538, 32'sd0.07538792361520971, 32'sd-0.02413835335152065, 32'sd0.04282101656228173, 32'sd-0.056788135473671626, 32'sd-0.08693746815165372, 32'sd-0.009145749062051211, 32'sd0.08980139272185401, 32'sd0.0011259657483438906, 32'sd-0.0798895598094352, 32'sd-0.06462755517825146, 32'sd-0.08368133197497074, 32'sd-0.041764473484273354, 32'sd-0.04440334367394549, 32'sd-0.015046032661817045, 32'sd-0.11209128070403097, 32'sd-0.050602067011427034, 32'sd0.047760563537989534, 32'sd0.1094863327086416, 32'sd0.016821127634785885, 32'sd-0.036747918081554885, 32'sd-0.025296246311784502, 32'sd-0.07068498563388062, 32'sd0.01233554805702218, 32'sd-1.1838991741610665e-126, 32'sd-0.004464188084108469, 32'sd0.06304538026889422, 32'sd-0.0015757289082508508, 32'sd0.020428930398369623, 32'sd0.033344184238885334, 32'sd-0.063513934726331, 32'sd-0.08130883872743117, 32'sd-0.02299091432237321, 32'sd-0.11701468353150735, 32'sd-0.005172420549285332, 32'sd0.028369418231663758, 32'sd-0.037550490643441334, 32'sd-0.008745859637007995, 32'sd-0.03519332321881584, 32'sd-0.15244571787731004, 32'sd0.0291837819645346, 32'sd0.03632410136858959, 32'sd-0.03950857589153225, 32'sd-0.16658286640994396, 32'sd-0.009874168414207017, 32'sd0.010557996555371431, 32'sd0.07473910683652106, 32'sd-0.010534783246376451, 32'sd-0.0271993015057297, 32'sd-0.04354067196035859, 32'sd-0.012150094334583292, 32'sd0.08561290742896836, 32'sd0.0563485683081023, 32'sd-0.03061234483450969, 32'sd-0.016235660146148023, 32'sd0.03088714499638526, 32'sd0.0646622480722488, 32'sd0.054472816069438414, 32'sd0.017544659208875785, 32'sd0.037948921995937676, 32'sd-0.047579433266613444, 32'sd-0.09327457140078432, 32'sd-0.16684970182817213, 32'sd-0.14021528291140195, 32'sd-0.06608255388645105, 32'sd-0.1688436352916836, 32'sd-0.10226871415187948, 32'sd-0.043991411130469185, 32'sd0.06204341217668981, 32'sd0.053933335378455086, 32'sd-0.10347545318245137, 32'sd0.007997268252104566, 32'sd0.02585502246902688, 32'sd0.052734128586905425, 32'sd-0.03445120073944198, 32'sd0.021779989802756795, 32'sd-0.10950950505033756, 32'sd-0.0069215127819918934, 32'sd-0.052522090054564305, 32'sd-0.03501878439109612, 32'sd0.056565937246411215, 32'sd0.023834965281539375, 32'sd-0.048674422846239844, 32'sd-0.07131547861628486, 32'sd-0.02975809343493863, 32'sd-0.004942299481404587, 32'sd0.015770047646178818, 32'sd0.02673485922588408, 32'sd0.06295276690879717, 32'sd-0.06854240120255539, 32'sd-0.15235544196274883, 32'sd-0.1501225625331208, 32'sd-0.08885048234679263, 32'sd-0.09065381992685467, 32'sd0.10549532898651723, 32'sd0.12886687831760255, 32'sd0.14497223814661095, 32'sd0.02150143798939338, 32'sd0.09065807584017804, 32'sd-0.07775104876779906, 32'sd0.032537804558248694, 32'sd-0.10402771784956369, 32'sd0.006977343597420168, 32'sd-0.03392859167862157, 32'sd-0.07193132135819025, 32'sd0.12658422619480947, 32'sd-0.11643978872439556, 32'sd0.0006224341932275135, 32'sd2.0423729795724607e-123, 32'sd0.038709682030162056, 32'sd0.01878211479726572, 32'sd-0.040211692575138354, 32'sd-0.1138421891193757, 32'sd-0.03454525275179122, 32'sd0.034423710318585314, 32'sd-0.05514748127947244, 32'sd0.07705809227844003, 32'sd0.011256984216850958, 32'sd0.014602344402722175, 32'sd-0.05046767051101915, 32'sd0.03267167435384521, 32'sd-0.03022596996595795, 32'sd0.11585256560475517, 32'sd0.06873006141722246, 32'sd-0.00441208273358555, 32'sd0.056527201996377605, 32'sd0.07972632420599055, 32'sd-0.013501765948029905, 32'sd-0.051440102713853866, 32'sd-0.12879149123296507, 32'sd0.05007844395600343, 32'sd-0.02035993010244613, 32'sd-0.005919567853226121, 32'sd0.047433458776779014, 32'sd-0.09339567507520281, 32'sd0.04455069283456344, 32'sd0.09450372879347228, 32'sd-0.07550299212786964, 32'sd0.03269772631515699, 32'sd-0.01632284159438125, 32'sd-0.12230386155993805, 32'sd-0.04502006984451715, 32'sd0.03999969712434302, 32'sd0.091681272638163, 32'sd-0.004553609467041741, 32'sd-0.05283279290738991, 32'sd-0.011245004628226139, 32'sd0.04289257872936706, 32'sd0.06637244815126694, 32'sd0.049329634533123314, 32'sd0.0402956260475176, 32'sd-0.07997469881189391, 32'sd0.03288885457730663, 32'sd-0.023483486009057, 32'sd0.004288354013012202, 32'sd-0.06198159646350014, 32'sd-0.004413356603926042, 32'sd0.03024960061275407, 32'sd0.007874954452991174, 32'sd-0.10161059754361314, 32'sd0.03512594744397867, 32'sd0.004253962101634625, 32'sd-0.12362527243987965, 32'sd0.0751386827805371, 32'sd0.07443217738462309, 32'sd0.08677417199681431, 32'sd-0.010680874070349013, 32'sd-0.011167340283900115, 32'sd0.025017447814663682, 32'sd-0.13780194373969562, 32'sd0.05864375974312838, 32'sd-0.06942759991208815, 32'sd0.050063545116647755, 32'sd0.013601443991897723, 32'sd0.07035476468389605, 32'sd0.0919467821751195, 32'sd0.004424861540091178, 32'sd0.05254136383913594, 32'sd0.028258837806811644, 32'sd0.043226677841353776, 32'sd0.07970549575761801, 32'sd-0.01776623230122242, 32'sd-0.06896790260096, 32'sd0.042743843575000696, 32'sd-0.029053680524964334, 32'sd-0.037254296479612765, 32'sd-0.03571373384501233, 32'sd0.061572155765910866, 32'sd0.002531884583445842, 32'sd-0.0030793523754732662, 32'sd0.007336972073930899, 32'sd0.028446762597243325, 32'sd-1.4581985043470176e-123, 32'sd-0.0013644187895677084, 32'sd0.012369237974631655, 32'sd-0.05369658365329343, 32'sd0.011409548544712982, 32'sd-0.08637314996613144, 32'sd-0.062113046678647, 32'sd-0.03725495701789098, 32'sd-0.16783329621210386, 32'sd-0.01083504839971032, 32'sd-0.055233709780076225, 32'sd0.07007106121373703, 32'sd0.13688901090882236, 32'sd0.09058286812803497, 32'sd0.12211179809915865, 32'sd0.05012734482922657, 32'sd0.007391246877372352, 32'sd0.012271441477953173, 32'sd-0.004088639357809922, 32'sd0.014955618734905154, 32'sd0.04709781123953205, 32'sd0.11415700201314252, 32'sd0.08436961181638836, 32'sd-0.003037350319822528, 32'sd0.06899636655045757, 32'sd0.037369241884657435, 32'sd0.047558523938046555, 32'sd-1.6345144834157188e-125, 32'sd2.1679130518559944e-124, 32'sd1.0366498564069416e-121, 32'sd0.03233119407169889, 32'sd-0.08657732358591734, 32'sd0.04574963585461075, 32'sd0.0034387060367177466, 32'sd0.027243198857982532, 32'sd-0.06351738861490076, 32'sd-0.08806022690290224, 32'sd0.03173333742471109, 32'sd-0.1974623859488681, 32'sd-0.058307947599445104, 32'sd0.05472187980582389, 32'sd0.06418916026261182, 32'sd0.07822895195559565, 32'sd-0.09467344666730193, 32'sd0.0625622995367078, 32'sd-0.0442245802009799, 32'sd0.03293142703911676, 32'sd0.05316853292987471, 32'sd0.1553169893526387, 32'sd0.0709720159340253, 32'sd-0.004214399478724939, 32'sd-0.07996496388606689, 32'sd-0.05732838292097672, 32'sd0.03983897107000034, 32'sd0.02876330060968817, 32'sd8.491399854191707e-121, 32'sd2.9447261336044833e-116, 32'sd1.5179688935247605e-116, 32'sd0.06420893778247705, 32'sd-0.10161250606112121, 32'sd0.03299584942773496, 32'sd-0.12337096729842181, 32'sd0.04010139745739486, 32'sd-0.07583599646768545, 32'sd0.06207862981459074, 32'sd0.027244237511862977, 32'sd0.07539676723618917, 32'sd-0.025243276402649374, 32'sd-0.013437933340794597, 32'sd0.09693377365504424, 32'sd0.03574070357706226, 32'sd-0.14359109053657726, 32'sd-0.05489618528808751, 32'sd-0.15393763966268922, 32'sd0.0624974236751976, 32'sd0.14807099983766867, 32'sd-0.003545713264758565, 32'sd-0.04659450428905474, 32'sd-0.04817256512027751, 32'sd-0.05744017564264101, 32'sd-0.04282258505895422, 32'sd-0.06772814195863291, 32'sd-0.0010817299747388172, 32'sd4.872085329399167e-123, 32'sd1.6395299135921879e-122, 32'sd-7.362662974243192e-117, 32'sd-4.3449762728536436e-123, 32'sd0.014372163268553702, 32'sd0.0071775935561292255, 32'sd-0.056247373067246, 32'sd-0.09479510646576758, 32'sd-0.0881846096233174, 32'sd0.14896718365351236, 32'sd0.06615779977622688, 32'sd-0.059271057482984925, 32'sd0.17602895938893226, 32'sd0.12280844087761476, 32'sd-0.13215847407381023, 32'sd-0.10723302708324167, 32'sd0.03376090206047358, 32'sd0.023790165064909528, 32'sd-0.04119161440507366, 32'sd0.07299780199710201, 32'sd0.09222672093479613, 32'sd0.07778638755373032, 32'sd0.04724656676725254, 32'sd0.13449177567958767, 32'sd-0.0865474968850267, 32'sd-0.007018647744871093, 32'sd0.0014825630315656315, 32'sd-1.5851204966200173e-120, 32'sd1.9251111413859114e-117, 32'sd8.585651499866185e-117, 32'sd3.7821856386815285e-118, 32'sd8.894731412321474e-127, 32'sd4.740838917229436e-126, 32'sd0.000726392678076127, 32'sd0.00925808166735694, 32'sd0.02472683097565239, 32'sd0.034975448821882256, 32'sd-0.014924497305759189, 32'sd0.002602703053697283, 32'sd0.036028837968252014, 32'sd-0.019806465878939403, 32'sd-0.0840204236544526, 32'sd0.10573066417240333, 32'sd-0.020586967043522093, 32'sd0.026600192939007082, 32'sd0.021840992163904165, 32'sd0.06915972089953837, 32'sd0.01985734799423081, 32'sd-0.0027386264845549895, 32'sd-0.017457613956372908, 32'sd-0.054957045619907885, 32'sd-0.11614770825836888, 32'sd0.006554034450805741, 32'sd-1.2740190650933717e-127, 32'sd-3.0316055114486778e-121, 32'sd-3.166971226549721e-121, 32'sd4.369479731304127e-123},
        '{32'sd-5.400397618577105e-118, 32'sd5.431932374293187e-126, 32'sd-4.387001136314275e-118, 32'sd8.278372773523777e-117, 32'sd1.742936514873311e-123, 32'sd-8.631192744785797e-121, 32'sd-1.8069376329350766e-123, 32'sd-6.148274038189464e-119, 32'sd2.0695181572414885e-117, 32'sd-1.802242919939413e-123, 32'sd4.7266820465790723e-126, 32'sd1.0239033724423782e-118, 32'sd-0.04941042559395878, 32'sd0.03170954270475814, 32'sd0.021911207783834687, 32'sd0.018944545489035177, 32'sd-7.122149071184838e-127, 32'sd9.852246996728982e-123, 32'sd-2.3420628565122498e-126, 32'sd-2.3421243748975947e-121, 32'sd-7.405436425002705e-128, 32'sd3.270162628798334e-125, 32'sd-2.1818074584038916e-121, 32'sd1.8185494381359664e-124, 32'sd2.132565368663857e-123, 32'sd3.170194693521869e-122, 32'sd8.164081745084701e-121, 32'sd-9.336253731131737e-119, 32'sd3.668670072613294e-123, 32'sd-1.947337881007463e-126, 32'sd-1.9427673703674813e-117, 32'sd-2.6393493495780213e-116, 32'sd-0.01357503750759087, 32'sd-0.02861618160788779, 32'sd-0.10454331319022735, 32'sd-0.007353600597215194, 32'sd0.029971456152523154, 32'sd-0.08254888493210465, 32'sd-0.018628647297795245, 32'sd-0.03732136478200415, 32'sd-0.05032419561305818, 32'sd-0.0059057483581015655, 32'sd0.08166008391913343, 32'sd0.10174532874695005, 32'sd0.014490079118658803, 32'sd-0.043728068239090305, 32'sd0.011076395939049, 32'sd0.0007815025030302697, 32'sd-0.08755857522780089, 32'sd-0.030052179481044838, 32'sd-0.013429861893672122, 32'sd-0.006570213107287839, 32'sd-1.2608362361692518e-117, 32'sd3.520421708009663e-120, 32'sd7.704174158451068e-117, 32'sd-7.643722310258198e-127, 32'sd4.826044331732849e-126, 32'sd-1.0310595330702083e-119, 32'sd-0.011851172743618526, 32'sd0.027851212407553932, 32'sd-0.04482095357640443, 32'sd0.06373751309294852, 32'sd-0.020151182656952798, 32'sd0.05103256164837318, 32'sd0.022119288255504948, 32'sd-0.017012289168276854, 32'sd0.09690112199626671, 32'sd-0.07454627795936741, 32'sd0.03252594266684899, 32'sd0.0379449839421351, 32'sd0.07116165127005955, 32'sd0.14754477591721873, 32'sd0.18808065091910825, 32'sd0.06180632962213875, 32'sd0.0974535962131722, 32'sd0.026159059636438102, 32'sd-0.028370630161286086, 32'sd0.03552689956807915, 32'sd-0.08547567161529948, 32'sd-0.01003966556573763, 32'sd-0.06093989454093107, 32'sd0.008611047344008225, 32'sd-7.83439000034306e-123, 32'sd2.5502138757147625e-124, 32'sd1.820641536199014e-126, 32'sd3.4440816858771335e-130, 32'sd0.05089371776001621, 32'sd-0.020873286755720963, 32'sd-0.023286139525637746, 32'sd-0.0242471584865605, 32'sd0.09545629919399828, 32'sd-0.043430414880270454, 32'sd-0.048968847792293185, 32'sd-0.007599682298931, 32'sd0.06638457873783862, 32'sd-0.009144588089111646, 32'sd0.11896634613733129, 32'sd0.0680598710656004, 32'sd0.10578046386021388, 32'sd-0.0020190874981089037, 32'sd-0.016493729545787705, 32'sd0.11678659396686727, 32'sd0.06272830530575887, 32'sd0.15696140583607587, 32'sd-0.025311866143462636, 32'sd-0.055986406892861496, 32'sd0.000854506722617175, 32'sd-0.11096185714694298, 32'sd0.020851289176499938, 32'sd-0.056613112047446026, 32'sd0.027590251666372235, 32'sd2.644848233762154e-119, 32'sd-6.076543272656405e-119, 32'sd0.06783783279174845, 32'sd0.06604371789129031, 32'sd-0.017476217988397085, 32'sd-0.06424416053690812, 32'sd0.04526320152190584, 32'sd0.049276854453289096, 32'sd-0.05530902053684857, 32'sd-0.07190264905279756, 32'sd-0.06638971748444293, 32'sd-0.12098545699379754, 32'sd0.017864626132792927, 32'sd-0.11797207276250896, 32'sd-0.003367291530544819, 32'sd-0.005667801681712683, 32'sd-0.022919144847943693, 32'sd-0.014897136371878955, 32'sd-0.07312866963520201, 32'sd0.01877200000803109, 32'sd-0.003464330982653013, 32'sd0.046325889341604164, 32'sd0.04144618421091012, 32'sd0.02128253128617711, 32'sd0.003916699151459433, 32'sd-0.03843561419353048, 32'sd-0.10297801395022216, 32'sd-0.07805831575597673, 32'sd0.02167697453351316, 32'sd1.9399817163666727e-125, 32'sd0.018891801460780164, 32'sd0.01847552123578798, 32'sd0.007022987665548019, 32'sd-0.03872815288352418, 32'sd-0.13402926766884246, 32'sd-0.1590020884961671, 32'sd-0.0080182491179213, 32'sd-0.1406367976914034, 32'sd-0.08309954483643432, 32'sd-0.17500620773703815, 32'sd-0.25945853885752246, 32'sd-0.11206074599547808, 32'sd-0.13697235775493302, 32'sd0.02612258776570009, 32'sd-0.022340856953397957, 32'sd0.06334263013697403, 32'sd-0.008135045806306127, 32'sd0.050509925147468, 32'sd0.058394518294339254, 32'sd0.022072395435074048, 32'sd0.07864891330355922, 32'sd0.14059760652082606, 32'sd0.1765145372037312, 32'sd-0.009912946332433552, 32'sd-0.14558269456909764, 32'sd-0.11043880063850495, 32'sd-0.05602290522921825, 32'sd2.697837316412401e-124, 32'sd-0.04734774345903202, 32'sd-0.0029461763833523473, 32'sd-0.009054479115271925, 32'sd0.01777386604055484, 32'sd-0.1930879802241207, 32'sd0.024494007414523778, 32'sd0.05093210262356053, 32'sd-0.126554386959729, 32'sd0.08460224411853709, 32'sd0.11857200982984355, 32'sd-0.0461705347416824, 32'sd-0.024893753609434986, 32'sd0.00038251118840348426, 32'sd0.0569852437483041, 32'sd0.1250997294055096, 32'sd0.08332060259020474, 32'sd0.04499060342684388, 32'sd0.009758279121779968, 32'sd0.06505583703706735, 32'sd-0.06797537882468487, 32'sd-0.04555517733323435, 32'sd-0.0752515048031956, 32'sd-0.014749143593854921, 32'sd-0.04998810628870198, 32'sd-0.09043023780889907, 32'sd-0.08735765070315024, 32'sd0.034651263483944976, 32'sd0.013095915706164092, 32'sd0.050032857777229434, 32'sd0.06319065387525462, 32'sd0.063308026825648, 32'sd0.015392482953843096, 32'sd-0.10235206966937359, 32'sd-0.029982474062051873, 32'sd0.0060301508821701015, 32'sd-0.07139282942042861, 32'sd-0.011366726687589762, 32'sd0.0460371646707829, 32'sd0.10284824934407492, 32'sd0.08572874534557799, 32'sd0.08054394845058077, 32'sd0.197567965022274, 32'sd0.146295016291878, 32'sd0.0652674153081006, 32'sd0.09240801231982536, 32'sd-0.06931834680512054, 32'sd0.021167895180223058, 32'sd-0.054818715895010875, 32'sd0.06398577851877262, 32'sd0.05186678850308776, 32'sd-0.018452449976482568, 32'sd-0.0543639423978031, 32'sd-0.1444510299827007, 32'sd-0.040568890984429284, 32'sd0.02428933219791067, 32'sd0.012566436623071702, 32'sd-0.11238003035248853, 32'sd0.06353553738783321, 32'sd0.002025617468471511, 32'sd-0.012481525400231074, 32'sd-0.06016001061696413, 32'sd-0.10277131345700348, 32'sd0.07513219265923764, 32'sd0.0965137708719334, 32'sd0.028297185772878458, 32'sd0.13579144966523418, 32'sd0.21523405986818694, 32'sd0.15947266954427927, 32'sd0.13824063555305993, 32'sd0.13882714729664225, 32'sd0.10574942337490505, 32'sd0.09536217826586572, 32'sd0.07217879809183315, 32'sd0.10095274759151263, 32'sd0.1021686018659821, 32'sd0.037949709233000166, 32'sd0.09236933344320754, 32'sd0.027807650136773086, 32'sd-0.026224430954411654, 32'sd-0.19660717287054427, 32'sd-0.07612410525107924, 32'sd-0.020571373870761456, 32'sd-0.05031112247622053, 32'sd-0.017353447634835283, 32'sd0.07926122291521552, 32'sd-0.0454941002400839, 32'sd-0.07005752262267761, 32'sd-0.07336200619936531, 32'sd-0.023559326584196336, 32'sd0.19600511756285524, 32'sd0.07034271293599131, 32'sd0.18033646201261075, 32'sd0.15076003922787165, 32'sd0.17636614913233065, 32'sd0.01966330967476042, 32'sd0.0810390117833252, 32'sd-0.03771854473563508, 32'sd-0.08615870290012277, 32'sd-0.018103598862496226, 32'sd0.0832742962172786, 32'sd0.01633346361298197, 32'sd0.08379131211389818, 32'sd0.12957558846394945, 32'sd0.005918902285291222, 32'sd-0.03191592120973215, 32'sd0.03511539401107626, 32'sd0.010893668117207812, 32'sd-0.05308251429991282, 32'sd-0.06958915134691551, 32'sd-0.04978597329768033, 32'sd-0.03263670152439872, 32'sd-0.005086789237702749, 32'sd-0.03106560140021123, 32'sd-0.02039400943276936, 32'sd0.09500846924879959, 32'sd0.003040435868227141, 32'sd0.003953063607767373, 32'sd0.16364574955081215, 32'sd0.10819200327229414, 32'sd0.1506430051853041, 32'sd-0.014848817610327383, 32'sd-0.07934088749792441, 32'sd-0.07256932937019381, 32'sd-0.08308955364491455, 32'sd-0.1663261583803159, 32'sd-0.3696478941870368, 32'sd-0.09427664269010025, 32'sd0.03108499364970245, 32'sd0.05922507516072512, 32'sd0.14016809094717916, 32'sd0.12781026191830128, 32'sd0.021514809041485408, 32'sd0.07863685058408128, 32'sd0.00997596866117685, 32'sd-0.05802255586247231, 32'sd-0.0971227953780945, 32'sd-0.0015004147793050632, 32'sd0.013258113640646212, 32'sd-0.025830771970901528, 32'sd-0.01979272666882322, 32'sd-0.023683130394775955, 32'sd0.05791044099163495, 32'sd0.09039534555071956, 32'sd0.04283270169141579, 32'sd-0.022897565206339142, 32'sd0.06778229781036088, 32'sd-0.028318922884215916, 32'sd-0.14350794357411198, 32'sd-0.049678795309001426, 32'sd-0.17300856465832332, 32'sd-0.25611427760075195, 32'sd-0.3330805328282242, 32'sd-0.2991708851917284, 32'sd-0.24485246169429387, 32'sd-0.06088506294941001, 32'sd-0.03746542385050798, 32'sd0.12626708620562171, 32'sd0.2304162437250916, 32'sd0.09102708665020942, 32'sd0.03992535089558249, 32'sd0.11510724800016915, 32'sd0.07147244224499118, 32'sd-0.16364075979428683, 32'sd-0.00024059132466862699, 32'sd0.008664097836525947, 32'sd-0.03889893274695648, 32'sd-0.06359939382449707, 32'sd0.03198853340591245, 32'sd0.032273751473150473, 32'sd-0.08472597703270088, 32'sd-0.007182219302036263, 32'sd0.08042889010992839, 32'sd-0.15215170893826566, 32'sd-0.12520620834966442, 32'sd-0.11630286243344397, 32'sd-0.14887261050147982, 32'sd-0.20013169740650075, 32'sd-0.2466882187963665, 32'sd-0.359679955593304, 32'sd-0.170078125331621, 32'sd-0.326614580146886, 32'sd0.050715673865997776, 32'sd0.20436880180823347, 32'sd0.09529309709413103, 32'sd0.11357647719855196, 32'sd0.03260271381368236, 32'sd0.07449783494314516, 32'sd-0.06977531554049077, 32'sd-0.06029917323692979, 32'sd-0.10715217475000571, 32'sd0.0056479145328892704, 32'sd-0.117125141658311, 32'sd-0.15897916261330178, 32'sd-0.03479517113399398, 32'sd0.052704043970301054, 32'sd0.014484983620827984, 32'sd-0.0779037329268685, 32'sd-0.042749965905512395, 32'sd0.0522131726931286, 32'sd-0.17640909773149455, 32'sd-0.17565582675140742, 32'sd-0.21680819767398157, 32'sd-0.0689382955365229, 32'sd-0.0222948582209971, 32'sd-0.2337636535649205, 32'sd-0.12064463129861808, 32'sd-0.09742857764501704, 32'sd-0.04627201832482409, 32'sd-0.0366449807488072, 32'sd0.06259762421774816, 32'sd0.010888859438617515, 32'sd0.061557693872694545, 32'sd0.0982497403523447, 32'sd0.038669283448400024, 32'sd0.007453920748569031, 32'sd-0.08500167318219765, 32'sd-0.07083950680962825, 32'sd-0.157204880179601, 32'sd-0.11412481944476607, 32'sd-0.09607580354234707, 32'sd-0.0830328315125516, 32'sd-0.0726742032545809, 32'sd-0.05210750229154526, 32'sd0.015824809447087255, 32'sd-0.02103671802715234, 32'sd0.01709972630083107, 32'sd0.014789837305499431, 32'sd-0.12367854636833875, 32'sd-0.14986134609505555, 32'sd-0.019812046845571692, 32'sd0.04830467153608844, 32'sd0.023478246273572537, 32'sd-0.16888766486118986, 32'sd-0.0387705874157719, 32'sd0.13125766804029995, 32'sd0.06136883204282395, 32'sd0.12282616545332824, 32'sd0.08669866918660546, 32'sd0.1819773027793238, 32'sd0.11808642683161313, 32'sd0.008449456826076234, 32'sd0.05613080965430083, 32'sd-0.05469700069937896, 32'sd0.06912081798118429, 32'sd0.021264928992564273, 32'sd-0.12849499192830122, 32'sd-0.07786329403947607, 32'sd0.027891718521566133, 32'sd-0.006816805591904247, 32'sd0.041547409573919815, 32'sd-0.021464328470741183, 32'sd-0.0485091356006452, 32'sd-0.03478797877639677, 32'sd-0.03170576089926459, 32'sd-0.03378744381294481, 32'sd-0.058791245316659684, 32'sd-0.0003929981494325085, 32'sd0.11067058808540264, 32'sd0.10105628043430445, 32'sd0.09702453560781905, 32'sd0.011763811028936932, 32'sd0.07041895748508982, 32'sd0.06767200587595512, 32'sd0.09819096374289399, 32'sd-0.006168034564264401, 32'sd0.060432672221346524, 32'sd0.037832922027869274, 32'sd0.05114716187154046, 32'sd-0.0359731497889509, 32'sd-0.022157979026228007, 32'sd0.04254107190859552, 32'sd-0.10225752944836888, 32'sd-0.09066808252257544, 32'sd-0.14582627530511164, 32'sd0.05066655181471479, 32'sd-0.10211823506562157, 32'sd-0.022589854484289178, 32'sd0.04815119027182943, 32'sd-0.061912850227173015, 32'sd0.02760608913326776, 32'sd0.09866878686666647, 32'sd0.0927016630089085, 32'sd-0.008661856530743122, 32'sd-0.02142126310519355, 32'sd-0.00983822375161978, 32'sd0.06773489013167333, 32'sd0.05051030834955662, 32'sd-0.031912486152830585, 32'sd-0.037420082036808425, 32'sd-0.015307513769824945, 32'sd-0.013499372332077009, 32'sd-0.02072201877258869, 32'sd0.002624580845041834, 32'sd0.012567176919584087, 32'sd0.10706777824352617, 32'sd-0.03470962997389955, 32'sd-0.06589234051630061, 32'sd0.0548621319897686, 32'sd-0.030015939210138138, 32'sd-0.13512912589539983, 32'sd-0.07373860243702182, 32'sd-0.15732709553334331, 32'sd-0.03878935970291099, 32'sd0.04320931228720311, 32'sd-0.02958227581010094, 32'sd-0.12204187345992855, 32'sd-0.05774532975975335, 32'sd-4.8522818140868755e-123, 32'sd0.024320013743730735, 32'sd0.07440013248367988, 32'sd-0.049049048865836, 32'sd0.06441144879340514, 32'sd0.0349650226964295, 32'sd-0.024193115967271465, 32'sd0.01156071492792956, 32'sd-0.024307992604293553, 32'sd-0.10365444481516257, 32'sd0.04455984902513621, 32'sd-0.010303969060557694, 32'sd0.05110767035763506, 32'sd0.04312539511321478, 32'sd0.2532307758000882, 32'sd0.19822165590618368, 32'sd0.02940440428216462, 32'sd-0.04949865111739283, 32'sd-0.030332265984044066, 32'sd0.09031372458613143, 32'sd-0.023228828219765525, 32'sd-0.15057751924625862, 32'sd-0.13923571335732285, 32'sd-0.01083121602810688, 32'sd0.02603369365984738, 32'sd0.03329278569600049, 32'sd-0.03665369567374479, 32'sd-0.022830609183000488, 32'sd0.01098880511798349, 32'sd0.032947881287899196, 32'sd0.08845247563571024, 32'sd0.010257975748045975, 32'sd-0.008049146327899449, 32'sd-0.025571994899728036, 32'sd-0.00023518802661616636, 32'sd-0.10645948708710568, 32'sd-0.049460130132721686, 32'sd0.05119631972209923, 32'sd0.04297093363424338, 32'sd0.08202835731568674, 32'sd0.013627481648430612, 32'sd0.03844215052427004, 32'sd0.03215930204335804, 32'sd0.037789582809459606, 32'sd0.11723630442291526, 32'sd0.08919618922374534, 32'sd0.017112815511263185, 32'sd0.08040479329076966, 32'sd-0.027876825770487064, 32'sd-0.05614105527193067, 32'sd0.011829144777014872, 32'sd-0.09304246356771241, 32'sd0.05802116176291653, 32'sd-0.07562440099330318, 32'sd-0.035580882257831764, 32'sd0.06691668862313521, 32'sd0.016639610895908253, 32'sd-0.04752732947444114, 32'sd-0.053525369271350313, 32'sd-0.0020408624426740433, 32'sd0.08923126341067689, 32'sd0.0018512309178325519, 32'sd0.12417002805530528, 32'sd0.03815594139594268, 32'sd0.04785977500212541, 32'sd-0.030301554490637074, 32'sd0.06838381322670838, 32'sd-0.0033607863776962646, 32'sd0.04259140076467268, 32'sd0.15784086305730977, 32'sd-0.03190420185041009, 32'sd0.020825472353074755, 32'sd0.08435339067648398, 32'sd0.00048154429874898284, 32'sd-0.004130580595851766, 32'sd0.10108132588252514, 32'sd-0.015196837394632765, 32'sd-0.023829958392516854, 32'sd-0.03373037938504356, 32'sd-0.06701137279680049, 32'sd0.009187411373006231, 32'sd-0.0312244571745338, 32'sd0.07720627531615704, 32'sd0.03580309802192192, 32'sd1.6071579544455723e-125, 32'sd-0.02599507673052038, 32'sd-0.0020033927276378186, 32'sd-0.056080973038429835, 32'sd0.06856669781627996, 32'sd-0.03401744923092918, 32'sd-0.013582223423572468, 32'sd0.13176155009959004, 32'sd0.08266236060991472, 32'sd0.0633919878926157, 32'sd0.1264046672844808, 32'sd0.002120962925759389, 32'sd0.07863674402799176, 32'sd-0.027647788372154175, 32'sd0.07197360605304118, 32'sd-0.013866903751423333, 32'sd-0.026628835002264126, 32'sd-0.03401135691940309, 32'sd0.10752443626574962, 32'sd0.12217626055299356, 32'sd-0.056990326285616476, 32'sd0.019988510781870646, 32'sd0.03421587555678856, 32'sd-0.009424240540744177, 32'sd-0.06687349180336705, 32'sd-0.052648487050442755, 32'sd-0.008827758138923393, 32'sd0.017609344733083197, 32'sd0.08718416020317139, 32'sd-0.03427509653763867, 32'sd-0.027817142428663472, 32'sd0.06660014542576484, 32'sd0.12980968464073225, 32'sd-0.00757812113772631, 32'sd0.003273342098382598, 32'sd-0.017392799273138453, 32'sd-0.05756203799086215, 32'sd0.008500960431675978, 32'sd0.01639087248165447, 32'sd0.01484783492628481, 32'sd0.02005444992293059, 32'sd-0.02071650236417879, 32'sd0.00310383861447507, 32'sd-0.02872186962359049, 32'sd-0.0035755333944154687, 32'sd-0.023602205163361065, 32'sd0.03147051602779823, 32'sd0.02933144024691744, 32'sd0.11176126276575984, 32'sd0.11299703741641137, 32'sd-6.990305858939723e-05, 32'sd-0.15420118612618122, 32'sd-0.025461710352279867, 32'sd-0.0665749836427244, 32'sd-0.019343230032374585, 32'sd-0.022072826299488302, 32'sd-0.003054568896226003, 32'sd-0.06542216393059673, 32'sd-0.018618131510869617, 32'sd-0.05644460418493721, 32'sd0.020116211565230288, 32'sd-0.0268396620885568, 32'sd0.00283419057514323, 32'sd0.007670283456980331, 32'sd-0.07584822550518412, 32'sd-0.08810145350001604, 32'sd-0.11886080817974767, 32'sd-0.059715384722232236, 32'sd-0.10647961440595882, 32'sd-0.1131064147674236, 32'sd-0.07228070584672386, 32'sd-0.03793726028888092, 32'sd0.11548563750083676, 32'sd0.007997272123289188, 32'sd0.053606303952140666, 32'sd0.13364333854828836, 32'sd0.02166810513815114, 32'sd0.07180407078038542, 32'sd-0.03938411530524121, 32'sd0.0005568934104314614, 32'sd-0.015321002802909362, 32'sd-0.08172911599853484, 32'sd0.003272522228438417, 32'sd0.027509083404219824, 32'sd-3.361045783435032e-114, 32'sd-0.007419672798686111, 32'sd-0.0018815223474719165, 32'sd-0.0984564303759683, 32'sd-0.0869605173608241, 32'sd0.044552349856961646, 32'sd-0.032713298412914406, 32'sd0.08078603396312156, 32'sd0.02108149636776796, 32'sd-0.02479822958641923, 32'sd0.040497510470699924, 32'sd-0.044064053366299163, 32'sd-0.12871406762320736, 32'sd0.07110375624302759, 32'sd-0.09130129762484837, 32'sd0.02469722233622725, 32'sd-0.02473754873674242, 32'sd-0.08377812524647518, 32'sd0.0017944848532989652, 32'sd0.07717926670768367, 32'sd-0.0807573302049743, 32'sd0.04343379690397063, 32'sd-0.008693941742783906, 32'sd0.028958859424956226, 32'sd0.0052964285697194345, 32'sd-0.02912577176475756, 32'sd0.050523475430946894, 32'sd1.0673999320826812e-115, 32'sd2.1112631437676714e-117, 32'sd4.039978621375058e-124, 32'sd0.006034702298768793, 32'sd0.028619493594050683, 32'sd-0.009122658877917357, 32'sd0.044138180244639925, 32'sd-0.040738819326665995, 32'sd-0.09176697826755782, 32'sd-0.05018891748905786, 32'sd-0.054057287301757226, 32'sd0.04921707453989652, 32'sd0.04592916623540397, 32'sd-0.10493424039660414, 32'sd-0.031582244762872635, 32'sd0.04330733909884565, 32'sd-0.05528154639980015, 32'sd-0.003112629978824955, 32'sd0.030143782247984984, 32'sd-0.02125717051268958, 32'sd0.034916033577716415, 32'sd0.041380136904176315, 32'sd0.016177672310924734, 32'sd-0.00508902142972719, 32'sd-0.023446042434109502, 32'sd0.037545261985376714, 32'sd-0.06148304037074163, 32'sd0.002715745616906134, 32'sd3.3977921408183965e-126, 32'sd-1.52589638915939e-126, 32'sd1.0494509012128743e-125, 32'sd-0.018297989511897414, 32'sd-0.02763889530534753, 32'sd0.04774887717000045, 32'sd0.03586684992834846, 32'sd-0.020953575038298013, 32'sd0.03685550705055481, 32'sd0.018559478997285408, 32'sd0.06242921445550505, 32'sd-0.059486225828317786, 32'sd-0.08384129507450881, 32'sd0.07134569924655247, 32'sd-0.04092416893110837, 32'sd-0.04014039932847899, 32'sd-0.06286540842905779, 32'sd-0.008273373582898681, 32'sd-0.08572716498927485, 32'sd-0.008930281025582203, 32'sd-0.024638610017141755, 32'sd0.04120565843163857, 32'sd0.041068292598861175, 32'sd-0.06467433320356733, 32'sd0.010968017279669773, 32'sd0.036842657810150545, 32'sd-0.013561219761625647, 32'sd0.01829367153407469, 32'sd-1.3258807869345736e-115, 32'sd6.917847708580934e-115, 32'sd-6.529057531403441e-117, 32'sd2.042271707292538e-127, 32'sd-0.008140378308875179, 32'sd-0.03571532801720249, 32'sd-0.028752664881580386, 32'sd-0.053586863857406256, 32'sd-0.031501489227578366, 32'sd-0.09706084930066684, 32'sd-0.02043000399208848, 32'sd0.0026499245121494454, 32'sd-0.011921892143558004, 32'sd-0.057614092293012946, 32'sd-0.0640293691633624, 32'sd-0.11423102899453011, 32'sd-0.01901290265597704, 32'sd-0.04965177624245217, 32'sd-0.06595430991985288, 32'sd-0.14644547387692583, 32'sd-0.003262163661502666, 32'sd0.04872167223474364, 32'sd0.08971005569830127, 32'sd0.049783883874400914, 32'sd-0.08033020689875632, 32'sd0.018934437720695724, 32'sd0.047812956019922415, 32'sd-2.4049294787245785e-124, 32'sd3.4985518606666513e-124, 32'sd2.959251071608447e-115, 32'sd1.7590774791035644e-123, 32'sd-6.983705763093978e-117, 32'sd2.4133302199405486e-120, 32'sd-0.005785975754721138, 32'sd0.05797392250351543, 32'sd0.07687652292101554, 32'sd0.028351335715292757, 32'sd0.027078500266017727, 32'sd-0.004741494548328616, 32'sd0.09064478743096853, 32'sd-0.000806826565491319, 32'sd-0.02108301311513144, 32'sd0.09012454265964931, 32'sd-0.04319338076503648, 32'sd0.06012115112599947, 32'sd0.09068405189181325, 32'sd-0.02615077926010013, 32'sd-0.005957030747367376, 32'sd0.020195642664739395, 32'sd0.11980027236977456, 32'sd0.006258736316596228, 32'sd0.008191656903370911, 32'sd-0.03836586429379757, 32'sd-5.0202214709876144e-126, 32'sd-3.54124001540152e-114, 32'sd-3.989442414070437e-117, 32'sd4.897604369054098e-115},
        '{32'sd2.0027088315277625e-117, 32'sd3.123567941103747e-120, 32'sd1.057519559528862e-118, 32'sd-9.300493132437136e-127, 32'sd-2.9962933820531993e-127, 32'sd-3.0948651258306706e-121, 32'sd2.6340312250816685e-123, 32'sd-2.0422114804775566e-124, 32'sd-6.84867482609618e-126, 32'sd-1.291500216768575e-119, 32'sd2.908206289697022e-126, 32'sd-5.459754626225916e-120, 32'sd0.01056036205229222, 32'sd0.050699855454458716, 32'sd0.09320622593772755, 32'sd0.05526219143532874, 32'sd1.1349132350033611e-125, 32'sd-4.3559859286977917e-126, 32'sd-4.084087079511281e-115, 32'sd3.661859427036072e-116, 32'sd8.991440393654014e-120, 32'sd-5.372058926323692e-118, 32'sd-2.2469655796523232e-120, 32'sd6.807477013404848e-126, 32'sd4.703820131921468e-123, 32'sd-1.9586232015159992e-118, 32'sd1.1565035611731549e-126, 32'sd4.376113406011664e-126, 32'sd8.094302793935578e-128, 32'sd1.673371356806822e-116, 32'sd1.7980600081754662e-121, 32'sd-1.742341110376131e-123, 32'sd-0.0037752890306875105, 32'sd0.0017831376062848205, 32'sd-0.05081737617767148, 32'sd0.03526809867808324, 32'sd-0.010825931165121937, 32'sd0.010113453829779176, 32'sd0.02251693854572923, 32'sd0.06678278843785168, 32'sd-0.08287658487331509, 32'sd0.06434069060575137, 32'sd0.1169780154781603, 32'sd0.10803445460830244, 32'sd-0.033224432299819404, 32'sd-0.03996517077924478, 32'sd0.04709842955396514, 32'sd-0.02224250685779812, 32'sd0.06776031339267614, 32'sd0.04453474595613866, 32'sd-0.015469398746228286, 32'sd0.012681153172180494, 32'sd-6.432755531642888e-117, 32'sd-3.796162721960975e-122, 32'sd-1.2565676988985642e-124, 32'sd3.534129144129361e-116, 32'sd3.85359796525277e-118, 32'sd-2.0849984048962897e-127, 32'sd0.0015775354586921165, 32'sd0.06607708089955563, 32'sd0.0003438406069445414, 32'sd-0.04678737532276284, 32'sd0.016976655762597385, 32'sd-0.09376361336922627, 32'sd0.08742822993771873, 32'sd0.05892537750094465, 32'sd0.1083906849403364, 32'sd-0.016502785490253653, 32'sd0.013963252268934788, 32'sd-0.04713023185224444, 32'sd0.015405060990242345, 32'sd0.0410163755567823, 32'sd-0.06763094038253235, 32'sd0.08380601717525832, 32'sd-0.019942578999948953, 32'sd-0.0013733089050097687, 32'sd0.07220520955749982, 32'sd0.05356835576317154, 32'sd0.01535713605593476, 32'sd0.09187877233829338, 32'sd-0.0769809753600609, 32'sd0.0306902350154249, 32'sd-3.5389525547232303e-118, 32'sd3.1389646074189595e-120, 32'sd-4.2598510758694415e-126, 32'sd4.2863322879434313e-125, 32'sd-0.010331990737269533, 32'sd-0.017891154229698093, 32'sd0.0004996199528103754, 32'sd0.11274987003586426, 32'sd0.061905679981079945, 32'sd0.062112037339222305, 32'sd0.09076436739719976, 32'sd0.042748812485107986, 32'sd-0.013192398329085309, 32'sd-0.09519925126038592, 32'sd-0.08690510509612895, 32'sd-0.038169829440938274, 32'sd-0.10845577209945204, 32'sd-0.16969610162792473, 32'sd-0.18197292629281708, 32'sd-0.12364348275495571, 32'sd0.07012885560189382, 32'sd-0.020991041281773447, 32'sd-0.07450953215123313, 32'sd-0.11712815065272342, 32'sd-0.03676891719531863, 32'sd-0.01935745454253679, 32'sd-0.0041664958913865645, 32'sd-0.09865545128616339, 32'sd-0.005129894344277181, 32'sd1.677840752006976e-125, 32'sd1.0253945716518678e-124, 32'sd0.04465315084329719, 32'sd-0.02147639232707166, 32'sd-0.003384737468025839, 32'sd-0.17649855581820006, 32'sd-0.08956924222714079, 32'sd-0.15065479311013005, 32'sd-0.0015691237897135551, 32'sd-0.12416368488141427, 32'sd-0.12563992016477246, 32'sd-0.11190914104773912, 32'sd-0.23115555529719542, 32'sd-0.16689963265652885, 32'sd-0.18424041053884635, 32'sd-0.08699703263754875, 32'sd-0.1480722767205641, 32'sd-0.024255820559492387, 32'sd0.005922362219166198, 32'sd-0.05732708498593987, 32'sd-0.04869448573476628, 32'sd-0.07290870125415437, 32'sd0.1719801048056599, 32'sd0.05674806745243005, 32'sd0.03692603124402905, 32'sd0.08365457934452547, 32'sd0.03507545361785342, 32'sd-0.009945307477673734, 32'sd0.0016840065181741397, 32'sd3.6557870358834e-116, 32'sd0.020896660295846175, 32'sd-0.026016037700032187, 32'sd-0.07984793763002158, 32'sd0.05782024865801049, 32'sd-0.08474400405015187, 32'sd-0.06067758265943557, 32'sd-0.12795694624851559, 32'sd-0.062089328693985354, 32'sd-0.1262534144106347, 32'sd-0.09670113565686093, 32'sd-0.0827408822174577, 32'sd-0.10707315444411356, 32'sd-0.22518050491241376, 32'sd-0.05571665429332444, 32'sd0.02198357897493251, 32'sd-0.061806191717282334, 32'sd-0.0652537047795635, 32'sd-0.06702871501261368, 32'sd-0.06111558556472035, 32'sd0.0033676694869803413, 32'sd0.13246497261651968, 32'sd0.012899965649297285, 32'sd0.05578583076527834, 32'sd0.041535378287904774, 32'sd-0.02155758287215628, 32'sd0.07897210520996552, 32'sd0.06569381462268231, 32'sd-5.897493840798514e-128, 32'sd0.018615960036281364, 32'sd-0.11130076634407239, 32'sd0.04100233547089204, 32'sd-0.040751913570152204, 32'sd-0.04968337126143506, 32'sd-0.13151721093373533, 32'sd-0.10739049334490423, 32'sd-0.15098311123652766, 32'sd-0.04246286792457626, 32'sd0.029085794502910024, 32'sd-0.004578547624855238, 32'sd0.06855244754161872, 32'sd0.016607743834244307, 32'sd0.08759240032668295, 32'sd0.014887342187055156, 32'sd-0.09811402194121545, 32'sd0.036459580774371246, 32'sd-0.18455733516927453, 32'sd-0.20221776171494932, 32'sd-0.11976688780239367, 32'sd-0.05339542707474754, 32'sd-0.026953299487637507, 32'sd0.04977683312830569, 32'sd0.0568004824463878, 32'sd0.12556700495107934, 32'sd0.13220591526420872, 32'sd-0.04644674540957482, 32'sd0.008619740590637482, 32'sd0.079479917235747, 32'sd0.0027044420810865355, 32'sd-0.02400014569369457, 32'sd-0.0030617385195983817, 32'sd-0.044857407524307225, 32'sd0.013795314897654022, 32'sd-0.0726905905884701, 32'sd-0.004496197991474901, 32'sd0.09763278600105041, 32'sd0.09479433194928875, 32'sd0.007872498231768353, 32'sd0.013290784426174328, 32'sd0.1280685949419897, 32'sd0.07423406686093147, 32'sd-0.0009953043136516455, 32'sd-0.008561204256312648, 32'sd-0.1002231943397679, 32'sd-0.12303015449942951, 32'sd-0.1733558441627324, 32'sd-0.18093137706208848, 32'sd-0.16861851498690603, 32'sd-0.05479758913463798, 32'sd-0.08815683719269195, 32'sd0.05295539673034191, 32'sd0.14833535763905348, 32'sd-0.001888977976718321, 32'sd-0.03912763136775761, 32'sd0.0017629205519740863, 32'sd-0.0553219159185031, 32'sd0.0927123239083247, 32'sd0.04051371638972216, 32'sd0.049889863534993466, 32'sd0.013021174296561347, 32'sd-0.011683246053475671, 32'sd0.0166138259367802, 32'sd0.07967499450815105, 32'sd0.13774537379126267, 32'sd0.2818586700738004, 32'sd0.1561985520982834, 32'sd0.15912699511621767, 32'sd0.06621646636297229, 32'sd0.05327814065593633, 32'sd0.06883544781164608, 32'sd0.030002168394858038, 32'sd0.04146131785990782, 32'sd0.07940076250949407, 32'sd0.04248528492052481, 32'sd-0.09620650268495898, 32'sd-0.09238740582146773, 32'sd-0.14667593495380193, 32'sd-0.04869755273130505, 32'sd0.05009999752552507, 32'sd-0.012105091378570224, 32'sd0.03151959326736343, 32'sd0.021378456526355272, 32'sd0.06179370956201389, 32'sd-0.06964180136816478, 32'sd-0.0067279257551121465, 32'sd0.017736471123196068, 32'sd-0.01866170902940242, 32'sd0.11154610211287996, 32'sd0.15132881656699065, 32'sd0.07620697308536113, 32'sd0.09780511233625214, 32'sd0.25387486698979567, 32'sd0.23685772816048234, 32'sd0.14245843551034987, 32'sd0.22958726337184068, 32'sd0.14049501536396058, 32'sd0.205315343255916, 32'sd0.08666237604028457, 32'sd0.1510308233161099, 32'sd0.05616871204653152, 32'sd-0.008967471458211139, 32'sd-0.03567707924109136, 32'sd0.020532856770916624, 32'sd-0.09686697655783619, 32'sd-0.042551834073790186, 32'sd0.11200713927212813, 32'sd-0.04010878820358794, 32'sd0.0614335257302941, 32'sd0.03815557543542288, 32'sd-0.04384336559862262, 32'sd0.0372631227832018, 32'sd-0.05307103360564503, 32'sd0.03835483462046816, 32'sd-0.07883262506972845, 32'sd-0.006076500741106123, 32'sd0.0136911180886642, 32'sd0.15014186769529372, 32'sd0.02202737699558469, 32'sd0.1552854233134249, 32'sd0.2357016387909781, 32'sd0.12784161655335932, 32'sd0.1676243450547216, 32'sd0.08212592732305263, 32'sd0.09272796414670144, 32'sd0.1208399536744603, 32'sd0.12751217078340127, 32'sd0.1572898371205678, 32'sd0.10944460448936724, 32'sd-0.06897822050593537, 32'sd0.04135999798077511, 32'sd0.02194570623386416, 32'sd0.043329848842107534, 32'sd-0.08938214887361404, 32'sd-0.009250839780866762, 32'sd0.035768939588497944, 32'sd0.012231011921045636, 32'sd-0.006952625696137555, 32'sd0.02801439300926244, 32'sd-0.01702070654448772, 32'sd-0.0002513979317000491, 32'sd0.03677830386007218, 32'sd0.052225680202044156, 32'sd0.02088674558661064, 32'sd0.06338911774500217, 32'sd-0.03272254679380758, 32'sd-0.014386135222920928, 32'sd-0.08516883299511151, 32'sd-0.028680533281537607, 32'sd0.049575113551871115, 32'sd-0.003240030945247525, 32'sd0.033344848076473296, 32'sd0.15690733269251314, 32'sd0.21412194368333773, 32'sd0.15658991640475353, 32'sd0.1038839679794657, 32'sd0.1288815834705366, 32'sd0.030954320573789895, 32'sd-0.12796962320702054, 32'sd-0.08477065808207983, 32'sd-0.0798477367022186, 32'sd-0.015034035288736806, 32'sd0.011283944490884065, 32'sd-0.01548153354526656, 32'sd0.07370911350193649, 32'sd-0.08307654208480193, 32'sd-0.011170572931130711, 32'sd0.05608086983123948, 32'sd0.062351963639147245, 32'sd-0.0626568212295664, 32'sd0.027550502924764186, 32'sd0.06752451779935638, 32'sd-0.061361330610431676, 32'sd-0.060763697862688516, 32'sd0.00199162819645738, 32'sd-0.10980385447121002, 32'sd-0.10753164247048506, 32'sd-0.21583724209385685, 32'sd-0.08610342148893475, 32'sd-0.05043307560087284, 32'sd0.036177657900124054, 32'sd0.0995676765190309, 32'sd0.02250634106028836, 32'sd0.03447978047471736, 32'sd-0.057683882665138506, 32'sd-0.06773527995085411, 32'sd-0.07388578064920473, 32'sd-0.04579478915705774, 32'sd-0.04513463932292243, 32'sd-0.10116665830302775, 32'sd0.026946764053643563, 32'sd-0.08522416675104534, 32'sd-0.0006238416855183554, 32'sd0.05563774881815234, 32'sd0.04270555537395343, 32'sd0.018100465663009508, 32'sd0.060275388837356496, 32'sd0.01434584442001468, 32'sd-0.04786104310691632, 32'sd0.02291104942157063, 32'sd-0.06750339964335145, 32'sd-0.04219987865646702, 32'sd-0.07706913876821227, 32'sd-0.00930969112140364, 32'sd-0.19668656915944957, 32'sd-0.11429792356965202, 32'sd0.062471079400953936, 32'sd0.0675932552748957, 32'sd0.11803497082791176, 32'sd0.11585221842131398, 32'sd0.004943567731547858, 32'sd0.04904611280368766, 32'sd-0.06533894452978202, 32'sd0.020298744170452403, 32'sd-0.1790907032822198, 32'sd-0.09121306896248309, 32'sd-0.12131576421648949, 32'sd0.016706118921339035, 32'sd-0.053299295784659584, 32'sd0.09731771480963809, 32'sd0.04193603851591298, 32'sd-0.05956226189946458, 32'sd-0.04921973811098683, 32'sd-0.0811027167126815, 32'sd-0.04253610991617456, 32'sd0.05011671429068872, 32'sd-0.05435615431749324, 32'sd0.059134792470865755, 32'sd-0.13996292255502574, 32'sd-0.07348710894721648, 32'sd-0.12477096317090242, 32'sd0.0019602592959137716, 32'sd-0.10371189492517449, 32'sd-0.044456477686392305, 32'sd-0.026844491745554217, 32'sd-0.05376007900779359, 32'sd0.018631649439237133, 32'sd-0.07542268262582112, 32'sd-0.06882786147741744, 32'sd-0.16941847243295444, 32'sd-0.06100511260733803, 32'sd-0.07089899839433635, 32'sd-0.10113705289714289, 32'sd0.023335756940274212, 32'sd-0.013852497580730792, 32'sd-0.06363799724776983, 32'sd0.12050468387829026, 32'sd0.10313438705341875, 32'sd-0.0019683048434972475, 32'sd0.05803963332242211, 32'sd0.010275195253217875, 32'sd0.030452373226660872, 32'sd-0.13160555503422508, 32'sd-0.10460457406097053, 32'sd-0.0765427787184494, 32'sd-0.03618683121414575, 32'sd-0.10102546338414949, 32'sd-0.04374484101536918, 32'sd-0.0957041019473804, 32'sd-0.03458358731312462, 32'sd-0.004029353408968606, 32'sd0.01172037121591946, 32'sd-0.028508390310059813, 32'sd-0.14740516015038757, 32'sd-0.15112223173317943, 32'sd-0.0707532730341359, 32'sd-0.12908356511738828, 32'sd-0.05483851995340911, 32'sd-0.035153093090071585, 32'sd0.03726593875400257, 32'sd0.04930160429738771, 32'sd0.051157830451050684, 32'sd0.040582332078811394, 32'sd-0.018948637311369997, 32'sd0.018495199014239853, 32'sd0.08616191508689133, 32'sd0.00975468373052423, 32'sd0.06706426765357573, 32'sd0.004940234889078474, 32'sd0.03303598898239937, 32'sd0.043882857203690034, 32'sd-0.05762972089363382, 32'sd-0.06615581595747513, 32'sd-0.06891607054570614, 32'sd0.03569927120768459, 32'sd0.09689757223982073, 32'sd-0.020022747029385116, 32'sd0.0990568100777311, 32'sd0.11733998801765222, 32'sd0.021735056657351794, 32'sd-0.0014743035613687615, 32'sd-0.00929843729179223, 32'sd-0.05555744953589241, 32'sd-0.0738625234020813, 32'sd-0.06846881291747448, 32'sd-0.0835176171586758, 32'sd-0.009996003151178443, 32'sd-0.03616940677130406, 32'sd0.042204433031866544, 32'sd0.08677328449343273, 32'sd0.08586031341392125, 32'sd0.1714781468391773, 32'sd0.07141275699586626, 32'sd0.13043312124554504, 32'sd-0.009163945755939028, 32'sd0.07806376249075059, 32'sd-0.019878059294963446, 32'sd-1.0225900570597205e-120, 32'sd-0.0058054963297701975, 32'sd-0.013432499808920922, 32'sd-0.07689362509292677, 32'sd-0.043312102126622815, 32'sd-0.07603875180745737, 32'sd0.012976708730354416, 32'sd0.0074543627893866315, 32'sd-0.02627640930073675, 32'sd-0.05168969055399283, 32'sd-0.05315202216269978, 32'sd-0.029940441114460484, 32'sd0.05755094038944836, 32'sd0.05670865441734828, 32'sd-0.057944211757873836, 32'sd-0.05807997295642133, 32'sd-0.0666864826825929, 32'sd-0.031066948126932357, 32'sd-0.04652027175347368, 32'sd0.12559104129776638, 32'sd0.03631946257422844, 32'sd0.09792061344413171, 32'sd0.13748924804023874, 32'sd0.042143223351662665, 32'sd0.023866026474497787, 32'sd0.11412375583000359, 32'sd0.10585393628521396, 32'sd-0.031111605735903415, 32'sd-0.02921979020880614, 32'sd-0.07817843291232278, 32'sd0.023926550498366783, 32'sd-0.01727852848183487, 32'sd-0.012059780448757315, 32'sd-0.07395531328869351, 32'sd-0.08949002431698139, 32'sd-0.024338147847100994, 32'sd-0.11462214594453098, 32'sd0.02981799790236883, 32'sd0.019647778279774045, 32'sd0.05161111851730446, 32'sd-0.003735691629835776, 32'sd-0.0827978040454517, 32'sd-0.1029263857115562, 32'sd-0.150268461289741, 32'sd-0.11802049842289096, 32'sd0.12593598653110266, 32'sd0.09081604197410394, 32'sd0.05896857172379481, 32'sd0.06345172850134002, 32'sd0.020012328868979967, 32'sd-0.01001777756881521, 32'sd0.011516222237321334, 32'sd-0.05214215995652155, 32'sd0.013486044932239517, 32'sd0.1042152840729329, 32'sd0.0864372346940506, 32'sd0.03650804738158695, 32'sd0.03548355349829753, 32'sd-0.008844212880254545, 32'sd-0.036837825053869636, 32'sd0.022904731740158123, 32'sd-0.008053790753080284, 32'sd-0.18338805343058734, 32'sd-0.09525530826295399, 32'sd-0.01632677734079972, 32'sd-0.07167589351951148, 32'sd-0.06798414078851907, 32'sd-0.06530363360989574, 32'sd-0.14321979751448138, 32'sd-0.21710292862598388, 32'sd-0.07630611257069939, 32'sd-0.07633013113051573, 32'sd-0.06284061761799103, 32'sd0.05811536962066196, 32'sd0.12822922371145445, 32'sd0.15400597258639606, 32'sd0.12298360082092037, 32'sd0.06397622386475277, 32'sd0.01848125380509791, 32'sd-0.09466941195215726, 32'sd-0.04742635224857519, 32'sd-0.04422162079871323, 32'sd0.005857002301530881, 32'sd0.04539282288488097, 32'sd-6.059633453074024e-127, 32'sd-0.03716485152321992, 32'sd-0.07482480887381347, 32'sd-0.0958033012705229, 32'sd0.018926578945816286, 32'sd-0.011940107629686288, 32'sd-0.131617281045919, 32'sd-0.08257119549867298, 32'sd-0.1258171739716925, 32'sd-0.21226872524087298, 32'sd-0.14927621821715834, 32'sd-0.04926418636136183, 32'sd-0.20115707951914288, 32'sd-0.22562684905458646, 32'sd-0.14424179742070187, 32'sd-0.16007615039815873, 32'sd-0.060470572185053, 32'sd0.06726486502927523, 32'sd0.02309407653236356, 32'sd0.058822962947401594, 32'sd0.04264868365105404, 32'sd0.011388742654008613, 32'sd0.05453474732271369, 32'sd0.030701556128949207, 32'sd0.06502011801012016, 32'sd0.164801174168073, 32'sd0.07159651770860892, 32'sd-0.011310520703020892, 32'sd0.008430944691372065, 32'sd0.0021619373885071636, 32'sd-0.06409409241468793, 32'sd-0.030667733110160283, 32'sd0.009917637630318695, 32'sd0.04049510272130486, 32'sd-0.05300433906914855, 32'sd-0.041615286412299474, 32'sd-0.0684465951706307, 32'sd-0.05298920056373875, 32'sd-0.022724081380293207, 32'sd-0.058924080785289656, 32'sd-0.025065144069342495, 32'sd-0.10044352961007484, 32'sd-0.17094743788106173, 32'sd-0.1438656511692497, 32'sd0.021493526427846247, 32'sd0.013665334040034012, 32'sd0.05710691034248584, 32'sd0.08490636993460571, 32'sd0.05128734044840027, 32'sd0.00741131525902104, 32'sd0.02968157691712736, 32'sd0.07119304289361439, 32'sd0.015320138553207227, 32'sd0.038611246813513564, 32'sd-0.025733068365986926, 32'sd0.0060501062140789815, 32'sd0.030220066173897393, 32'sd0.0019095557747880192, 32'sd-0.08737512564126698, 32'sd-0.05772818597359607, 32'sd-0.007791964319482026, 32'sd-0.036681278158703194, 32'sd0.025597074325967396, 32'sd-0.023405476094933316, 32'sd-0.1399943772751738, 32'sd-0.016703161738257147, 32'sd-0.10603072824721346, 32'sd-0.07248446903543757, 32'sd-0.040079705873643325, 32'sd0.06844188255222507, 32'sd0.08024700322265489, 32'sd-0.05056497195475698, 32'sd0.00891352543321739, 32'sd-0.013391670248380071, 32'sd-0.019416655362558766, 32'sd0.12753593387803336, 32'sd0.05535066214576633, 32'sd-0.023830910271959625, 32'sd0.09746294799898392, 32'sd-0.014794705393054802, 32'sd-0.015745735159602255, 32'sd0.05379568104788371, 32'sd-0.08266209440026344, 32'sd0.05637046525976251, 32'sd-9.150628451470442e-124, 32'sd0.0610471200715363, 32'sd-0.015895517821752227, 32'sd-0.030925340806388688, 32'sd-0.05978381856476225, 32'sd0.11135443956779711, 32'sd0.07348053202243504, 32'sd-0.039881835858732284, 32'sd-0.032109793447327305, 32'sd-0.052542398541747144, 32'sd-0.10027323164280413, 32'sd0.06007645675797128, 32'sd-0.12225255266785025, 32'sd0.025264947844555206, 32'sd0.04984116282641709, 32'sd0.1055776775228473, 32'sd-0.03347782792924559, 32'sd-0.06258305964383386, 32'sd0.09250756894264846, 32'sd-0.05692260311593194, 32'sd0.06237110520236969, 32'sd-0.054404176160842595, 32'sd0.07495185984309621, 32'sd0.023849238538552395, 32'sd0.06747956138822535, 32'sd0.013551990485690111, 32'sd-0.014722212793727492, 32'sd-1.6258292724299342e-115, 32'sd-1.347074688600092e-128, 32'sd-2.607175552083692e-124, 32'sd-0.008968072415464734, 32'sd-0.06641946583311746, 32'sd-0.061046768082400386, 32'sd0.07120745063907673, 32'sd-0.07726406333631877, 32'sd-0.0653432092686749, 32'sd-0.026249916245865604, 32'sd0.028657444132590734, 32'sd-0.04806447624003956, 32'sd-0.11527803110716722, 32'sd-0.19683898300385924, 32'sd0.05870980424553154, 32'sd-0.019408654290805048, 32'sd-0.0957834552598302, 32'sd-0.00018740928613198072, 32'sd-0.020771182322276534, 32'sd0.005857045405081812, 32'sd0.016112281779696484, 32'sd0.03920871147760061, 32'sd-0.08766986347162858, 32'sd0.06783707126701188, 32'sd0.029708189330978574, 32'sd-0.05672841403885281, 32'sd-0.019481966000875452, 32'sd0.010505550518442394, 32'sd1.6635198164328937e-125, 32'sd-8.719845174201025e-122, 32'sd-2.4222442437382866e-124, 32'sd0.014196262593054162, 32'sd-0.013340155581812925, 32'sd-0.0606131561740196, 32'sd0.014790975748096059, 32'sd0.09381004791647167, 32'sd0.0595180615461882, 32'sd0.1411577535643636, 32'sd-0.038876699520317984, 32'sd0.08524432043624099, 32'sd-0.05364414289476848, 32'sd0.13659212460256423, 32'sd-0.02370828270901881, 32'sd0.0586611778901981, 32'sd0.035540164963054496, 32'sd0.02977303898718843, 32'sd0.10054944652465418, 32'sd0.05483538212814064, 32'sd0.09454232184124867, 32'sd0.042565619747407024, 32'sd0.03246742332872188, 32'sd0.05512724502765343, 32'sd-0.03136889142362617, 32'sd-0.05870973947464815, 32'sd0.007541760994588208, 32'sd0.015884435787065297, 32'sd2.9919416877522526e-124, 32'sd1.1758495082178474e-118, 32'sd-3.126033319996652e-122, 32'sd1.1425937130578794e-119, 32'sd0.06818348159470138, 32'sd-0.08592758309936617, 32'sd0.09650225491674333, 32'sd0.07524731239988353, 32'sd-0.01608806786684564, 32'sd-0.005652263169492004, 32'sd0.031312066462528335, 32'sd0.09314550921855481, 32'sd0.032153591725164535, 32'sd0.15037897031165304, 32'sd0.06202437008307945, 32'sd0.05333949417539733, 32'sd0.12023243564671608, 32'sd0.08494206375138208, 32'sd0.081170427188602, 32'sd0.004197604900737957, 32'sd-0.0075516743050150145, 32'sd0.1008329844053142, 32'sd0.02087520879909137, 32'sd0.009068581738147596, 32'sd0.026933667984864802, 32'sd-0.04916868648188618, 32'sd0.01752130991629003, 32'sd7.457947442864361e-122, 32'sd1.510612028344739e-119, 32'sd2.3329743087706205e-124, 32'sd1.811814224650481e-123, 32'sd2.987369674528031e-121, 32'sd-1.0760266275953135e-118, 32'sd0.05248129419417932, 32'sd0.024422622758006433, 32'sd-0.0035055463741561427, 32'sd0.03349590146527081, 32'sd0.05918512297258716, 32'sd-0.08668497097528459, 32'sd-0.018746763991939492, 32'sd0.013155219311837442, 32'sd0.06595593607779167, 32'sd0.10023088529820731, 32'sd0.08462102601500958, 32'sd0.054914549205509006, 32'sd0.10792055412630501, 32'sd0.13788507423939902, 32'sd0.02959975486213463, 32'sd0.013739388724675401, 32'sd-0.007227755284599257, 32'sd0.08540905834583412, 32'sd-0.07414969074795644, 32'sd0.08476077245901228, 32'sd-1.1459214186767065e-126, 32'sd-5.023412987778039e-118, 32'sd2.6815259214518535e-124, 32'sd-5.157192448069864e-122},
        '{32'sd8.22828592159813e-117, 32'sd-6.604793893375367e-122, 32'sd6.31732217225114e-124, 32'sd-1.3954823288729262e-117, 32'sd2.6685365157472964e-117, 32'sd-3.6330376414606715e-122, 32'sd5.353363896417365e-123, 32'sd-1.4201829938783532e-118, 32'sd2.938976396279552e-121, 32'sd-6.100877292824609e-127, 32'sd-1.0715363107500377e-120, 32'sd1.2953871183426747e-117, 32'sd0.05350998993053539, 32'sd0.0687507652588213, 32'sd0.0452122480073532, 32'sd0.016412268288610386, 32'sd-2.1060757094160695e-117, 32'sd7.306867499867165e-124, 32'sd5.912566467125252e-115, 32'sd8.015146945809902e-119, 32'sd-3.9097871855212744e-119, 32'sd-5.907563096281192e-122, 32'sd-1.4933992210779228e-125, 32'sd2.9851420433892174e-123, 32'sd-1.536168664414421e-115, 32'sd2.303708980046002e-124, 32'sd-1.0197131110884565e-124, 32'sd3.7942404895723363e-128, 32'sd5.715277442258329e-120, 32'sd-1.835240495373716e-121, 32'sd8.609879026590098e-117, 32'sd3.9942591284056225e-115, 32'sd-0.003228627065406895, 32'sd-0.02362210372757555, 32'sd-0.011798245950096934, 32'sd-0.13074092648410973, 32'sd0.018079816550244057, 32'sd0.01323981788039662, 32'sd0.015349454994030278, 32'sd-0.004684822153800077, 32'sd0.044191471331012463, 32'sd0.06077290612336415, 32'sd-0.04035517926845138, 32'sd0.03826462050118897, 32'sd0.02055182034791932, 32'sd0.05973249648247548, 32'sd0.04542416194381097, 32'sd-0.022197017390735704, 32'sd0.008376889045945543, 32'sd0.026831894478775965, 32'sd0.0621369303755797, 32'sd0.03874945685712659, 32'sd-7.497577606240706e-124, 32'sd1.4716889927583814e-124, 32'sd7.68863716968933e-116, 32'sd-1.253868417858324e-123, 32'sd-1.752555316219484e-123, 32'sd1.7666166414845266e-117, 32'sd0.05163870640272244, 32'sd0.025854117710873342, 32'sd0.05949176695439977, 32'sd-0.0699295694864211, 32'sd-0.05882376483470701, 32'sd-0.02649772748021529, 32'sd-0.020129614563185617, 32'sd0.031757834094634674, 32'sd0.14657367636308788, 32'sd-0.04564614228876477, 32'sd0.07294585278724273, 32'sd-0.11234909655329454, 32'sd0.11421528012069625, 32'sd0.07907552990110873, 32'sd-0.05974145947760568, 32'sd0.1303002293923507, 32'sd0.0886858789870597, 32'sd-0.03843492116382617, 32'sd0.08505370947113614, 32'sd0.10613247853516797, 32'sd0.012507572592457586, 32'sd0.023882562246835812, 32'sd-0.005780146198516387, 32'sd0.04866897937293917, 32'sd1.8363042552761035e-121, 32'sd-2.774381001574941e-119, 32'sd-3.7551466321135254e-122, 32'sd2.1057773068864974e-117, 32'sd0.023101364967710262, 32'sd-0.08162079459995202, 32'sd-0.012202007420774737, 32'sd0.09533892141674288, 32'sd0.03338802438455792, 32'sd-0.04941785035287417, 32'sd0.18681911501092605, 32'sd-0.016202782318792054, 32'sd-0.03200096823106981, 32'sd0.1943662913445968, 32'sd0.04092017375754603, 32'sd0.04870125182220829, 32'sd0.18306250639094215, 32'sd0.16780894615254577, 32'sd0.026908895847062176, 32'sd-0.13735154212125666, 32'sd-0.01974509019194791, 32'sd0.0219886427940804, 32'sd0.0691790589216147, 32'sd0.04183953270351611, 32'sd-0.05212550266822303, 32'sd-0.04778650242469244, 32'sd-0.11375221546845617, 32'sd0.05045771624996778, 32'sd-0.01160337058417029, 32'sd1.0730891485385314e-119, 32'sd-4.7356061507698535e-117, 32'sd0.030294247687678126, 32'sd0.010592435882117677, 32'sd-0.004670964781628364, 32'sd-0.11318269721190574, 32'sd0.01241541356584401, 32'sd0.029183395743628354, 32'sd-0.002235264113694597, 32'sd0.09091693812923872, 32'sd0.03330475129521419, 32'sd0.19667353504831472, 32'sd0.15699192515188845, 32'sd-0.06153297133436686, 32'sd-0.019158950283468087, 32'sd0.038577204520690966, 32'sd-0.06378155117859577, 32'sd0.01051508758297989, 32'sd0.04930016361991231, 32'sd-0.06634954686821883, 32'sd-0.03441107139398005, 32'sd-0.10273950159775201, 32'sd-0.08471198846762353, 32'sd-0.10184668969663048, 32'sd0.01621051863601757, 32'sd-0.02132345786150713, 32'sd0.031876927736638805, 32'sd-0.00043220382427545685, 32'sd0.009332393133046622, 32'sd-2.0432305459581607e-121, 32'sd0.04371022966741778, 32'sd-0.024410042293208208, 32'sd-0.008514493775971068, 32'sd0.07145142753004304, 32'sd-0.0597752972570028, 32'sd0.09413931971303262, 32'sd0.05443725701649232, 32'sd0.06624133967752759, 32'sd0.11656538058776038, 32'sd-0.01991772224359242, 32'sd-0.09023677642515791, 32'sd-0.029022302735155825, 32'sd-0.05291120527354402, 32'sd-0.08679668416157671, 32'sd-0.0821406957991852, 32'sd-0.025919636989706545, 32'sd0.03532354477633989, 32'sd-0.15626502135706624, 32'sd-0.08693622533370646, 32'sd-0.08004382455151292, 32'sd-0.09222586141206227, 32'sd-0.2007257858412356, 32'sd-0.1228076818329236, 32'sd0.009088249794413252, 32'sd-0.01376753278642529, 32'sd-0.1265169327114532, 32'sd0.025579963372256324, 32'sd9.458912384628368e-121, 32'sd0.055467325459390274, 32'sd0.03663848861071297, 32'sd0.08464499516392171, 32'sd0.055278488708797396, 32'sd-0.05733019662730745, 32'sd0.05638767286507711, 32'sd-0.02484166892798963, 32'sd-0.035270378618053565, 32'sd0.09655035705399027, 32'sd-0.028668171666300927, 32'sd-0.024516451714497227, 32'sd-0.09719501586934383, 32'sd-0.12100627580206678, 32'sd-0.1517168813805901, 32'sd-0.01698031363532767, 32'sd0.07679238330103585, 32'sd-0.10867714815039074, 32'sd-0.202013721824277, 32'sd-0.15148169491066404, 32'sd-0.18863996455950188, 32'sd-0.25954721374256245, 32'sd-0.14214475324503448, 32'sd-0.19566042227761796, 32'sd-0.17085668312767055, 32'sd0.09339614619044431, 32'sd-0.07068469639369206, 32'sd0.0709818583680119, 32'sd0.060423533396723766, 32'sd-0.023189491607461653, 32'sd0.03561907935859266, 32'sd0.05534580900495827, 32'sd-0.024938460596045563, 32'sd-0.009025524205212136, 32'sd0.06259134608979791, 32'sd-0.07262253565945341, 32'sd-0.049199269501740174, 32'sd-0.11915371445284655, 32'sd-0.07010954377936807, 32'sd-0.12139034407328765, 32'sd-0.08075072266116902, 32'sd-0.05854666479451258, 32'sd-0.17629389249197294, 32'sd0.02595439805805745, 32'sd0.0030963961244455628, 32'sd-0.11612705450459826, 32'sd-0.08503968672689362, 32'sd-0.13750137811442978, 32'sd-0.146735689580709, 32'sd-0.18433329441540278, 32'sd-0.2365545722047505, 32'sd-0.2715469556974511, 32'sd-0.06656769550496502, 32'sd-0.002859861265597483, 32'sd-0.11556492371990931, 32'sd0.04912091094153917, 32'sd-0.009063921105293792, 32'sd0.05724879229801867, 32'sd-0.08582740181501627, 32'sd-0.16091155209214617, 32'sd-0.07349033366188422, 32'sd0.07510046550521567, 32'sd-0.05886010721226251, 32'sd-0.09851647277385447, 32'sd0.07367307457440528, 32'sd-0.08527231249158163, 32'sd-0.05796416107791656, 32'sd-0.13222531568658583, 32'sd0.02542723673211372, 32'sd-0.09427333326202991, 32'sd-0.09366207605611106, 32'sd0.058974115381143416, 32'sd0.1770798613720501, 32'sd-0.06336713146936328, 32'sd-0.03479259892138434, 32'sd-0.10955071897339523, 32'sd-0.033153950073294775, 32'sd-0.12557783079064969, 32'sd-0.121132852396927, 32'sd-0.19927539649065126, 32'sd-0.10654771550270228, 32'sd-0.0817065291888323, 32'sd-0.02837021207167607, 32'sd0.08373049443015934, 32'sd-0.01004052031674171, 32'sd0.03201696693929877, 32'sd-0.01368128918358866, 32'sd-0.03203390867090066, 32'sd0.041235240452672094, 32'sd-0.07514577668634956, 32'sd-0.03730237522724037, 32'sd-0.09761604937786514, 32'sd0.016136615707213524, 32'sd-0.01584956595670937, 32'sd0.01826167723749732, 32'sd0.0468811981378135, 32'sd0.046630662472510846, 32'sd-0.06660152786590631, 32'sd0.030773216511023778, 32'sd-0.01510404074220319, 32'sd0.0722742957635041, 32'sd0.021633306922332472, 32'sd-0.09631573537616421, 32'sd-0.02196775298642252, 32'sd0.07613439090806233, 32'sd-0.05533258850678814, 32'sd-0.0856265844266181, 32'sd-0.032966480623952174, 32'sd0.016380270548333523, 32'sd-0.038709074955838654, 32'sd-0.0008072533832590302, 32'sd0.024647692109047274, 32'sd0.04360415289618492, 32'sd-0.017145976003971185, 32'sd0.047969991114561766, 32'sd0.16177783286999192, 32'sd0.045220982905344015, 32'sd0.009827844115862239, 32'sd-0.024999600941791218, 32'sd-0.07490224024868271, 32'sd-0.042724361685096926, 32'sd0.004694500893306791, 32'sd0.061102663087050285, 32'sd0.037517141871261046, 32'sd-0.0013218276361310285, 32'sd-0.045558687278114726, 32'sd0.04275983544141059, 32'sd-0.20460874303700344, 32'sd-0.09199714823760302, 32'sd-0.09508924255510882, 32'sd-0.027614628829670543, 32'sd-0.029243306839347026, 32'sd-0.0038280797334887067, 32'sd-0.05443425325991365, 32'sd-0.1570322190751197, 32'sd0.0018313396697905947, 32'sd0.07267548587868689, 32'sd-0.1297212987415535, 32'sd0.04731463731124452, 32'sd-0.06274094423369973, 32'sd-0.039322122023001664, 32'sd-0.04581461473417223, 32'sd0.0312686986733083, 32'sd0.05113282784899512, 32'sd0.045169370896028724, 32'sd0.08238895727216718, 32'sd-0.06748295929303028, 32'sd-0.08536253532838388, 32'sd0.058587148567610596, 32'sd0.10703174816627803, 32'sd-0.02180973069998108, 32'sd-0.019937354857150376, 32'sd0.047067972771847585, 32'sd-0.06867356513945105, 32'sd0.009904504722230222, 32'sd-0.1336881909448939, 32'sd-0.14910490245899852, 32'sd-0.12490324038988386, 32'sd-0.10283779594949959, 32'sd0.02417546323425327, 32'sd-0.07342671894464997, 32'sd0.06181327279710185, 32'sd0.03877371769602203, 32'sd0.03811781097662211, 32'sd-0.009335039944435406, 32'sd0.06065402435135499, 32'sd-0.02891625794518135, 32'sd-0.07124429808896829, 32'sd0.048920041241744795, 32'sd-0.008320793662714574, 32'sd0.00933206377661125, 32'sd0.011646565174970026, 32'sd0.06704492822734842, 32'sd0.0039503671722769034, 32'sd-0.1518898710513728, 32'sd-0.040396754711848774, 32'sd0.08470473478612642, 32'sd0.061354166709046566, 32'sd0.19115608782375493, 32'sd0.05758259668818351, 32'sd0.033081981208846846, 32'sd-0.0019320857740554118, 32'sd-0.1117760478659594, 32'sd-0.19683128220815319, 32'sd0.11589145996782008, 32'sd-0.08628709314052885, 32'sd0.024828586179219077, 32'sd-0.12074914557751744, 32'sd0.09333006475166133, 32'sd0.10962799944668693, 32'sd0.08194736254411993, 32'sd0.08982626971656874, 32'sd-0.003975947308536387, 32'sd0.04251322609819309, 32'sd-0.0382255799095482, 32'sd0.002613088801557459, 32'sd-0.006745731306766082, 32'sd-0.006830266404289707, 32'sd0.015948019313036015, 32'sd-0.037038608592871974, 32'sd0.03916754514982628, 32'sd0.023981562474789827, 32'sd-0.09804824573495427, 32'sd0.030576530653265963, 32'sd0.1410346418749586, 32'sd0.1304304150267892, 32'sd0.11832777587787668, 32'sd0.06550119792531436, 32'sd0.03018573637754332, 32'sd0.18130319756039848, 32'sd0.05127060073181517, 32'sd-0.04037023813095771, 32'sd0.17722180068213947, 32'sd0.11334516845558883, 32'sd0.15346910523021182, 32'sd-0.030954150980706165, 32'sd-0.07324566001260009, 32'sd0.09326609580167727, 32'sd0.16641388403524088, 32'sd0.17422047580424063, 32'sd0.09633504734866552, 32'sd-0.015346712105842718, 32'sd0.025005748658594548, 32'sd0.08446055595116299, 32'sd0.020714124667514835, 32'sd-0.0066793498348313605, 32'sd-0.0027872222270212167, 32'sd-0.09873398152399372, 32'sd0.039304932843013646, 32'sd0.08729655558255071, 32'sd0.05328603235320562, 32'sd0.05995981792541116, 32'sd0.0761762960305002, 32'sd0.16460779644792325, 32'sd0.06032474312524451, 32'sd-0.047746326460922604, 32'sd0.12522412754555165, 32'sd0.11572919693656755, 32'sd0.06451380915379958, 32'sd0.06241387539581253, 32'sd0.17840059176059397, 32'sd0.027915314734257103, 32'sd0.12142241901961986, 32'sd0.04686414136787519, 32'sd0.03569512160261746, 32'sd0.030763846227814765, 32'sd0.0646126854772102, 32'sd0.11906478811248092, 32'sd0.08615356413996365, 32'sd-0.02071689229320395, 32'sd-0.027629563965134454, 32'sd0.056802023836825415, 32'sd-0.039832498627159735, 32'sd-0.05636228141613511, 32'sd-0.05446202294621481, 32'sd0.05452485869943161, 32'sd0.011873126136640605, 32'sd-0.08827449433232022, 32'sd0.10391517327531344, 32'sd0.09536314744305449, 32'sd-0.020709465800647472, 32'sd-0.056933350676544016, 32'sd-0.08727716846780463, 32'sd-0.14965040495523663, 32'sd0.0749055730628445, 32'sd0.12666576224899373, 32'sd0.06656886891664443, 32'sd0.060267092125623395, 32'sd0.19577335050690275, 32'sd0.04428855240129004, 32'sd0.1191726654869128, 32'sd0.08512514498070434, 32'sd0.06985186455380879, 32'sd-0.031594265464105264, 32'sd0.007380075448072443, 32'sd0.013102995436476767, 32'sd-0.008668668785883332, 32'sd0.03929347576155766, 32'sd-0.046140184268273716, 32'sd-0.05987904534204632, 32'sd0.008770727959568068, 32'sd0.03430169849634168, 32'sd0.043230346737749614, 32'sd0.08286892007641504, 32'sd0.011405879930876316, 32'sd0.00837479788690105, 32'sd0.11604166084103966, 32'sd-0.06781718471750868, 32'sd-0.11312533538928288, 32'sd0.013564895349197019, 32'sd0.04381529627828459, 32'sd0.049343985686476986, 32'sd0.07362254916132076, 32'sd0.03634688495911903, 32'sd0.16350960703069548, 32'sd0.14674129729229016, 32'sd0.037811319403026386, 32'sd0.09380553776040886, 32'sd0.18724881769650228, 32'sd0.11966053867289962, 32'sd0.08114417829098323, 32'sd0.0931294105839388, 32'sd0.06730999668140718, 32'sd-0.003431006551648999, 32'sd-0.014743320622099565, 32'sd0.010619615627577022, 32'sd0.007705575292952196, 32'sd0.045340417004983535, 32'sd-1.7807160367284377e-123, 32'sd-0.022567706684897954, 32'sd-0.02240033587725723, 32'sd0.045974375286995335, 32'sd-0.11690806126718203, 32'sd0.01807562502411905, 32'sd0.12822527300739395, 32'sd-0.1259359989711026, 32'sd-0.023972979476888565, 32'sd0.0018951255388688245, 32'sd-0.09917337834308025, 32'sd0.0042580413353334335, 32'sd-0.04104768766013874, 32'sd0.05819321154960036, 32'sd0.052720023436147144, 32'sd0.016455531957419722, 32'sd0.059301083589029316, 32'sd0.053888876778647246, 32'sd0.04319455658272052, 32'sd0.05304469273755365, 32'sd0.11127200988628816, 32'sd0.08336277006694252, 32'sd0.05096499292145122, 32'sd0.07319602799382181, 32'sd-0.06421037413750039, 32'sd0.0374133276093835, 32'sd-0.011836959057873218, 32'sd0.010533305122267361, 32'sd0.0026608283526064146, 32'sd-0.029220664605149688, 32'sd-0.0005767648155405278, 32'sd0.06375105622328646, 32'sd0.04156639957900568, 32'sd0.10120018392268078, 32'sd0.0851857013564164, 32'sd-0.023652489269772436, 32'sd-0.02603270529739451, 32'sd-0.01061435177766732, 32'sd-0.0006602822300982666, 32'sd-0.037426249278312375, 32'sd0.04208650702295924, 32'sd0.0013810131157286738, 32'sd-0.06119560404750626, 32'sd0.0684084861902167, 32'sd0.08529048520946104, 32'sd0.10206227468035474, 32'sd0.03252425674233437, 32'sd0.13273831151043577, 32'sd0.08150854314855109, 32'sd-0.05071929875859955, 32'sd0.09815851778051864, 32'sd0.15028090519734932, 32'sd-0.0635336024259656, 32'sd0.10197960106608621, 32'sd-0.049574045016748655, 32'sd-0.038947489913424824, 32'sd-0.005361328381822235, 32'sd0.03936510679158193, 32'sd0.023265026967892084, 32'sd-0.06671085349329708, 32'sd-0.05696567071450087, 32'sd0.07590475861935117, 32'sd0.05138706397035316, 32'sd0.017682057790980258, 32'sd0.01043869738400106, 32'sd-0.06161628699698784, 32'sd0.041711527429212955, 32'sd-0.012177916163773408, 32'sd-0.06619401845477711, 32'sd-0.09523031755029956, 32'sd0.006321718077012959, 32'sd-0.04840355014990815, 32'sd0.08014113548390964, 32'sd0.09794747008470411, 32'sd-0.05048459621883626, 32'sd0.05323815274845945, 32'sd-0.08938442013870318, 32'sd-0.016040328404483807, 32'sd0.158348895936856, 32'sd0.06317321518086734, 32'sd-0.12842930931880528, 32'sd0.06482923328063364, 32'sd-0.050092533141202704, 32'sd-0.014844093944495436, 32'sd-1.4140308202124866e-118, 32'sd-0.0854734214066791, 32'sd-0.06191687149631871, 32'sd0.09860095522853368, 32'sd-0.11191362205127785, 32'sd0.04704217103556534, 32'sd0.11950023705223968, 32'sd0.2136100340843088, 32'sd0.158047803702191, 32'sd0.03809534569168661, 32'sd0.07822466060533609, 32'sd0.025638818508497394, 32'sd-0.05447715368486031, 32'sd-0.012618614446803334, 32'sd0.022169107122482233, 32'sd-0.029991468792723873, 32'sd-0.007534839043625675, 32'sd-0.0861665248447718, 32'sd-0.05333094043204995, 32'sd-0.10702490329975596, 32'sd-0.11670266877546405, 32'sd-0.09614943719445179, 32'sd-0.09116316506059859, 32'sd-0.13387387385742083, 32'sd-0.049970193568177536, 32'sd-0.07015887940496508, 32'sd-0.015018026384006294, 32'sd-0.015705439637220483, 32'sd-0.03815742385606915, 32'sd0.00789167104701973, 32'sd0.030881772338848017, 32'sd0.14081193250446059, 32'sd-0.028291221773019615, 32'sd-0.07802962862801222, 32'sd0.0625166833255123, 32'sd0.13016524792608508, 32'sd0.05866722963936383, 32'sd0.1402254759982346, 32'sd0.09617265303778574, 32'sd-0.05109916985529311, 32'sd-0.07269322820327141, 32'sd0.15347343197349858, 32'sd0.08625044470030127, 32'sd-0.02606718789718381, 32'sd-0.037835080697383935, 32'sd0.012185159270737924, 32'sd-0.05611611632769523, 32'sd-0.11134011556741484, 32'sd-0.03792144542426387, 32'sd-0.05434305535141922, 32'sd-0.09673674520823408, 32'sd-0.01121970866475115, 32'sd-0.0930476133791323, 32'sd-0.012675103357407383, 32'sd0.044836016827848484, 32'sd-0.018278891568989358, 32'sd0.048479459580810236, 32'sd0.027994762451472293, 32'sd0.019116207346646295, 32'sd0.020665526042777417, 32'sd-0.1886098491582625, 32'sd0.06566689948569673, 32'sd-0.0811494014664244, 32'sd-0.02203899219893143, 32'sd0.09137114264239671, 32'sd0.11709417897775043, 32'sd0.11916238669330799, 32'sd-0.04016458472570479, 32'sd-0.023548632504247248, 32'sd0.06367594448316254, 32'sd-0.0542107633847787, 32'sd-0.08734803485591254, 32'sd-0.14756109834675796, 32'sd-0.1667445773091465, 32'sd-0.22794588510683542, 32'sd-0.12461771490589095, 32'sd-0.23493667526471315, 32'sd-0.06309184094011015, 32'sd-0.06830418517162035, 32'sd-0.08691048829222124, 32'sd-0.048603001139059965, 32'sd-0.046375591144739915, 32'sd-0.09031315938522361, 32'sd0.03993480763377734, 32'sd1.198095443632581e-122, 32'sd0.0040793803119737945, 32'sd0.10466880642410456, 32'sd0.08438554343547525, 32'sd-0.08710036933183492, 32'sd-0.0958038920351206, 32'sd-0.16299925897792195, 32'sd-0.16054001105519994, 32'sd-0.09344030951768204, 32'sd-0.041835768196967694, 32'sd0.038101331928982955, 32'sd0.030508774018709838, 32'sd0.011448217377985943, 32'sd-0.13830686438671422, 32'sd-0.050861616259880255, 32'sd-0.08674253613829616, 32'sd-0.22997960940157758, 32'sd-0.24974116664338303, 32'sd-0.30749417695361475, 32'sd-0.22670069419822048, 32'sd-0.09918046737773778, 32'sd-0.14667853097434966, 32'sd-0.12957460366442614, 32'sd-0.11549309664150408, 32'sd0.019694969108445145, 32'sd-0.02600418686360069, 32'sd-0.06165058002097417, 32'sd-1.4427042381675496e-124, 32'sd-1.3868465712519815e-120, 32'sd1.2066309496987264e-123, 32'sd0.050816427854068744, 32'sd0.053847211940293654, 32'sd-0.07969762226930129, 32'sd-0.10629494763310486, 32'sd-0.07860647703029613, 32'sd-0.1680241486492234, 32'sd-0.20127347345942817, 32'sd-0.018427591344157442, 32'sd0.014182698943303785, 32'sd0.02381023660465617, 32'sd-0.20021389672225787, 32'sd-0.15228993448146855, 32'sd-0.08243011946921341, 32'sd-0.17560193985869887, 32'sd-0.12158357456568866, 32'sd0.013551172541051251, 32'sd-0.15455106112670144, 32'sd-0.13432033487892814, 32'sd-0.04547238208965315, 32'sd-0.022029772915008933, 32'sd0.0031005687474371223, 32'sd-0.044275042966953025, 32'sd-0.019151250366280934, 32'sd-0.051319958564622424, 32'sd0.04994328334778428, 32'sd-2.7605661350592726e-120, 32'sd6.528611284973944e-127, 32'sd7.01663799943542e-117, 32'sd-0.04712251102787951, 32'sd0.005750764350817398, 32'sd-0.035068294212482684, 32'sd0.019891573199265298, 32'sd-0.014242730232772451, 32'sd-0.08052991451288155, 32'sd-0.17091106310902526, 32'sd-0.06729851301715536, 32'sd-0.10061951644107552, 32'sd-0.12977353397017774, 32'sd-0.11297499706822223, 32'sd-0.08794639440818139, 32'sd-0.055651773194137784, 32'sd0.013600517418775968, 32'sd-0.039054070031742306, 32'sd0.02308110104135277, 32'sd-0.08506803376989015, 32'sd0.054213171566859154, 32'sd0.04221849826090443, 32'sd-0.01128216301143938, 32'sd-0.052833901825165, 32'sd-0.11404721810462866, 32'sd-0.1039600222839051, 32'sd0.0011069932619792431, 32'sd0.013319375028793674, 32'sd1.6532149656673442e-127, 32'sd1.217460461416226e-117, 32'sd8.285202555880071e-123, 32'sd-1.0148999532190933e-120, 32'sd0.038950724374606144, 32'sd0.03674767955947893, 32'sd-0.026844957440071336, 32'sd-0.0008214871942984673, 32'sd0.0526526244310797, 32'sd-0.02173400648674629, 32'sd-0.13822681908473905, 32'sd-0.06465010394813561, 32'sd-0.06499867097428605, 32'sd-0.0076349692241646575, 32'sd-0.11528855853836421, 32'sd0.06706038560766985, 32'sd0.09085259645587615, 32'sd-0.1298358458313067, 32'sd-0.14996181925419616, 32'sd0.07516026830000205, 32'sd-0.007777556425282519, 32'sd0.024248803250752342, 32'sd-0.04153032299411742, 32'sd-0.055606397818281895, 32'sd-0.08589486392376904, 32'sd0.011969304816686958, 32'sd0.011788402051823499, 32'sd4.3099561793356744e-120, 32'sd4.911488275568927e-118, 32'sd-1.1289873003790373e-115, 32'sd2.52803167350443e-125, 32'sd-8.936941657912501e-126, 32'sd-1.5131928930865992e-115, 32'sd0.03165525227526127, 32'sd-0.011894577875125387, 32'sd0.050667287238531644, 32'sd0.013347615187605506, 32'sd-0.017534411476326114, 32'sd0.08033718088008852, 32'sd0.026638467253052363, 32'sd-0.058738847873579116, 32'sd0.1133494625631241, 32'sd-0.07628773124124559, 32'sd-0.06337695287915214, 32'sd0.03660869412484308, 32'sd0.04442193273488373, 32'sd-0.028727415510095826, 32'sd-0.0001735689122156633, 32'sd0.03035397574323279, 32'sd-0.045357825208243226, 32'sd-0.03474038015970955, 32'sd0.02722729223873418, 32'sd0.0026656432159756706, 32'sd-8.689091495581248e-116, 32'sd-2.355364290319504e-116, 32'sd-1.70655816702141e-115, 32'sd-9.870216650283846e-115},
        '{32'sd1.4412624027569554e-115, 32'sd1.09927803256746e-121, 32'sd1.8984483788088552e-122, 32'sd2.672374949462249e-124, 32'sd4.1959607021102765e-124, 32'sd-5.5683979295051445e-120, 32'sd2.008649480011873e-120, 32'sd-3.4576528745858203e-122, 32'sd2.9712067454403606e-116, 32'sd-1.751442892867451e-119, 32'sd-2.544234814539988e-124, 32'sd1.0587910486253967e-124, 32'sd0.11124254877288124, 32'sd0.12929779174036407, 32'sd0.0791153828834828, 32'sd0.062424131831286395, 32'sd4.172779833577278e-121, 32'sd3.3488354859697157e-121, 32'sd4.22949967156003e-125, 32'sd-8.057096005053537e-122, 32'sd1.37384975211794e-123, 32'sd-1.5211718034120487e-124, 32'sd8.287638907679845e-129, 32'sd-5.4049832395019245e-118, 32'sd6.888931556441369e-126, 32'sd-8.03056662832153e-116, 32'sd-3.971929665956306e-120, 32'sd-3.965751883381536e-119, 32'sd-7.364939746894961e-125, 32'sd-3.67203418377069e-123, 32'sd1.0534762963803974e-121, 32'sd1.127026098184548e-122, 32'sd0.13125169101609002, 32'sd0.07687145377105069, 32'sd0.006039320118820902, 32'sd-0.011782271352217523, 32'sd0.08964759221886656, 32'sd-0.053777700341948224, 32'sd0.07990319590619135, 32'sd-0.010791159455338201, 32'sd-0.0012676034654945311, 32'sd-0.0013991884841826078, 32'sd-0.0030707030852131973, 32'sd0.08245697261904449, 32'sd0.013030322873003628, 32'sd0.10567728953252944, 32'sd0.08119864237703088, 32'sd0.04444997990731334, 32'sd0.037851017384193844, 32'sd-0.005249057594056888, 32'sd-0.008009177229861013, 32'sd0.01681035753887628, 32'sd-3.7681738529394906e-122, 32'sd6.47880056164868e-116, 32'sd-1.2086430070900735e-118, 32'sd1.2961186975934233e-124, 32'sd-1.4738454540483557e-123, 32'sd1.0006792702553649e-120, 32'sd0.0066814953144968955, 32'sd-0.014313134709712657, 32'sd0.08187289363718879, 32'sd-0.05658326713235951, 32'sd-0.011417418265333743, 32'sd-0.0294450712815952, 32'sd0.0847029467959886, 32'sd0.07657956521202208, 32'sd0.07098159790754634, 32'sd0.040680602990803505, 32'sd-0.0363794711719017, 32'sd-0.11922282577321913, 32'sd0.10131085405710508, 32'sd0.07936879560962794, 32'sd0.02703325303291186, 32'sd-0.11943767277887035, 32'sd-0.03714424984029781, 32'sd-0.02182459441966256, 32'sd0.038692573869333, 32'sd-0.00236703315983512, 32'sd0.08085576854823727, 32'sd-0.001064041301652747, 32'sd0.03414837191725869, 32'sd0.01855513250687812, 32'sd1.6725974439954094e-116, 32'sd2.850049151739621e-118, 32'sd-1.561680391329774e-127, 32'sd-1.0802095225410632e-127, 32'sd0.029455780754793978, 32'sd0.016861287421219222, 32'sd-0.0027687361292638166, 32'sd-0.012023907702314977, 32'sd-0.1454942456694828, 32'sd-0.11680273226455769, 32'sd0.14512546005252977, 32'sd0.05098988707504584, 32'sd-0.09189504442909122, 32'sd-0.021068938184303877, 32'sd-0.03031986375013672, 32'sd-0.004264895195544624, 32'sd-0.10949483679635473, 32'sd-0.14356434486137779, 32'sd-0.07251066325261869, 32'sd-0.0804842929462814, 32'sd-0.01831404141394941, 32'sd0.05441982297086247, 32'sd-0.11166487213970004, 32'sd0.038966739267370536, 32'sd0.0727129693858424, 32'sd0.04105863286994548, 32'sd0.058252605548850096, 32'sd0.017406781918483688, 32'sd0.08995522076374354, 32'sd-8.57903601603451e-121, 32'sd-5.8806841085325475e-124, 32'sd0.03830166450193641, 32'sd0.08676398651525505, 32'sd0.04390167227630377, 32'sd-0.024802146183862322, 32'sd-0.08378360202938033, 32'sd0.052382179875423714, 32'sd0.01349854416405907, 32'sd0.08226625517495594, 32'sd0.017533313237378247, 32'sd0.12017809906086165, 32'sd-0.08144105400411317, 32'sd0.06316721112733747, 32'sd-0.09944599375570477, 32'sd-0.17602071834751465, 32'sd-0.16094489794933348, 32'sd-0.1839343731175084, 32'sd-0.20192571768501588, 32'sd-0.2099060484890046, 32'sd-0.09067686038865702, 32'sd-0.06539083419647192, 32'sd0.01212487240056999, 32'sd-0.04393966348383688, 32'sd0.00301600270929413, 32'sd0.013755911091075821, 32'sd0.03336938757032165, 32'sd0.04122667533135415, 32'sd-0.016344645241356946, 32'sd5.514725392189744e-118, 32'sd0.01156408595086212, 32'sd-0.024735245408029204, 32'sd-0.05189710220149768, 32'sd0.01521877179324665, 32'sd-0.08200419411622552, 32'sd0.07721876690311587, 32'sd0.08067420546283678, 32'sd-0.08103239360179988, 32'sd-0.04332070915282139, 32'sd-0.15829794029291647, 32'sd-0.11469245569286882, 32'sd-0.18267540856176206, 32'sd-0.11246852323541083, 32'sd-0.07324001863276959, 32'sd-0.05888794451854483, 32'sd-0.07147187058208683, 32'sd-0.14177311399520667, 32'sd0.0032915467801819267, 32'sd0.029098863371086383, 32'sd-0.13161249037429984, 32'sd-0.0833505745493432, 32'sd-0.014254194817519184, 32'sd-0.11722699049459519, 32'sd0.07650387212226975, 32'sd0.1280597931948288, 32'sd0.05016214699319651, 32'sd0.07874691944511197, 32'sd1.6994332236393667e-115, 32'sd0.10866687260086177, 32'sd0.014948763751656964, 32'sd0.06829095880914827, 32'sd-0.01765544261412703, 32'sd-0.10538195870036414, 32'sd-0.021296032328762853, 32'sd-0.004720957093145323, 32'sd-0.04092745463691774, 32'sd0.03178265799026472, 32'sd-0.002038217494717487, 32'sd-0.04645956700111619, 32'sd-0.05003668685686336, 32'sd-0.047218554032039964, 32'sd0.02106795565915083, 32'sd-0.008177783974986662, 32'sd0.03158141328565136, 32'sd-0.008300250220509793, 32'sd-0.12072575143221131, 32'sd0.06690124386130039, 32'sd-0.12030126103739062, 32'sd-0.1788672484812924, 32'sd-0.19478032181218768, 32'sd-0.038480637047454025, 32'sd-0.12754640612622165, 32'sd0.09193641284026195, 32'sd0.08652321506699204, 32'sd-0.024791759163175053, 32'sd0.04923836849026385, 32'sd0.06500231421468565, 32'sd-0.04307967967563173, 32'sd-0.04808295341889975, 32'sd-0.11123199458895996, 32'sd-0.017035491588102403, 32'sd-0.008594772358912975, 32'sd-0.05454221897033505, 32'sd-0.08297187940647521, 32'sd0.0716148877224281, 32'sd0.030690850821134427, 32'sd0.021220124545641105, 32'sd0.030007597949472907, 32'sd0.11310902869771597, 32'sd0.02540291191092135, 32'sd-0.1648043807040484, 32'sd-0.24125701747539027, 32'sd-0.168725215371703, 32'sd-0.19404452315657822, 32'sd-0.15239760132261282, 32'sd-0.05000367920429365, 32'sd0.02642504892733775, 32'sd-0.08728670691212309, 32'sd-0.09106047226335102, 32'sd-0.04659438393358678, 32'sd0.10282566898216078, 32'sd0.06883852866106271, 32'sd0.042428432653548745, 32'sd0.05019753387706269, 32'sd0.09939029373641384, 32'sd-0.02777120316236854, 32'sd-0.043838187020414095, 32'sd-0.06801546584454153, 32'sd-0.05707150803129855, 32'sd-0.04630130349358501, 32'sd-0.11263711031196139, 32'sd0.055228938015780854, 32'sd0.11268969735040663, 32'sd0.21115790735028858, 32'sd0.1437076697431075, 32'sd0.11089354637579317, 32'sd0.19240371542676224, 32'sd-0.0014738255236658032, 32'sd-0.043409979348948344, 32'sd-0.13497497506478692, 32'sd-0.16982702203275085, 32'sd-0.07678173073501601, 32'sd0.0654576087098226, 32'sd-0.03531868705149635, 32'sd0.005856339605569176, 32'sd-0.04632596320292995, 32'sd0.008410165647079061, 32'sd-0.11478721474189117, 32'sd-0.02058904738076047, 32'sd0.003737406452068268, 32'sd0.0037843892645964203, 32'sd0.12100008840240306, 32'sd0.07947618250950435, 32'sd0.1241040430616924, 32'sd0.015004411385517362, 32'sd0.02945983039290131, 32'sd-0.07351477081459067, 32'sd0.07107288603453435, 32'sd-0.030835469472883306, 32'sd0.02788749634212212, 32'sd0.017323474203110735, 32'sd0.16188203751735883, 32'sd0.025392352720703996, 32'sd0.06557852426632411, 32'sd0.07470420968308543, 32'sd0.09786976448666228, 32'sd-0.012990566798201375, 32'sd-0.12683848836527656, 32'sd-0.005468118997698141, 32'sd-0.05809741576026476, 32'sd0.13744083255217604, 32'sd0.13224295831816477, 32'sd0.17568233145744297, 32'sd0.08757586126313165, 32'sd0.016058621947078137, 32'sd0.05053382504110459, 32'sd-0.01923428893429511, 32'sd0.07701310118215851, 32'sd0.07643540126756818, 32'sd0.0017951972960572177, 32'sd-0.05786923713675997, 32'sd-0.019593530518708994, 32'sd0.033917405733285, 32'sd0.09262519047959197, 32'sd0.05315926972628068, 32'sd0.029855789859813648, 32'sd0.026683846481950456, 32'sd0.1109839408943406, 32'sd0.1698730668567955, 32'sd0.05238459085181985, 32'sd0.05643650088260882, 32'sd-0.04611272555937787, 32'sd-0.05926499591665115, 32'sd-0.13743013247869695, 32'sd-0.13076937740204617, 32'sd-0.024979972118380718, 32'sd-0.047525380045899145, 32'sd0.02523565713793209, 32'sd0.13545587363004283, 32'sd0.13177795361728623, 32'sd0.0752645121325773, 32'sd0.08309933054545585, 32'sd0.07392799476818486, 32'sd-0.05539926631955398, 32'sd-0.03360352049916576, 32'sd0.06200533831202539, 32'sd0.07677131604888732, 32'sd0.05415726388286991, 32'sd0.03533847341363439, 32'sd0.061515816887176764, 32'sd0.047881963433762754, 32'sd0.06718940048621917, 32'sd0.11524856415746239, 32'sd0.028525680987351587, 32'sd-0.013634005171496117, 32'sd0.08855644191646936, 32'sd0.07930767320416078, 32'sd-0.04101691536631977, 32'sd-0.0939126894193556, 32'sd-0.29090085615744565, 32'sd-0.19377943793080848, 32'sd-0.06221741996916156, 32'sd-0.08627975578387043, 32'sd-0.059270164422381234, 32'sd-0.04944164744008352, 32'sd-0.12458316385706449, 32'sd0.09327407603431079, 32'sd0.09860075585860381, 32'sd0.0995076592677296, 32'sd0.14428208506704088, 32'sd0.08805025241426442, 32'sd-0.09333846365652856, 32'sd0.031986303546581864, 32'sd0.09352346094509878, 32'sd0.05665852714073154, 32'sd0.003989700389724163, 32'sd0.04101423164698656, 32'sd0.00305122313197197, 32'sd0.03070173002906568, 32'sd0.09766008985255867, 32'sd0.08414335087193339, 32'sd-0.06906713031216453, 32'sd-0.011026756147713833, 32'sd0.005288205563351735, 32'sd0.001959905982072825, 32'sd-0.11377066276692493, 32'sd-0.28213586541997776, 32'sd-0.19232961669647664, 32'sd-0.12436124027744352, 32'sd-0.0031714623381323462, 32'sd0.18158270300516752, 32'sd0.17323661830195888, 32'sd-0.0323356160537685, 32'sd-0.08305356827174305, 32'sd-0.06440394565203031, 32'sd-0.05445399644354635, 32'sd0.007333620070859424, 32'sd0.13148198352134466, 32'sd0.08511270629126252, 32'sd0.0328598563607367, 32'sd0.02843603430128772, 32'sd0.022539612932085704, 32'sd0.01644387185926056, 32'sd-0.00595543615745334, 32'sd-0.0690398873982228, 32'sd-0.06303310720101112, 32'sd0.039175580838840304, 32'sd0.02854707115622282, 32'sd0.05142061689652867, 32'sd-0.080981846355598, 32'sd-0.028812671144472127, 32'sd-0.11558668095576681, 32'sd-0.2718095536466703, 32'sd-0.2567940457464846, 32'sd-0.14044802310012977, 32'sd-0.06474181397735577, 32'sd-0.008584959802865392, 32'sd-0.009650233439679823, 32'sd0.02460865030310176, 32'sd0.17195795517115892, 32'sd-0.004756255529919141, 32'sd0.06203134967757647, 32'sd0.007807460411441638, 32'sd0.03644925045018822, 32'sd0.08682501647665947, 32'sd0.04781146665370593, 32'sd0.005031509975361221, 32'sd0.1480042128842492, 32'sd0.007720713721194544, 32'sd0.004955141846038489, 32'sd0.010240574223265854, 32'sd-0.07922048169228559, 32'sd0.024156640954428103, 32'sd-0.005333920284118001, 32'sd-0.0044887317444858976, 32'sd-0.033500379954194845, 32'sd-0.005855620514062291, 32'sd0.07286674661251179, 32'sd-0.05865823390828058, 32'sd-0.0433307772917166, 32'sd-0.25439288271562926, 32'sd-0.11901507988429154, 32'sd-0.07675842525760124, 32'sd0.09997761780884697, 32'sd0.1536758728350421, 32'sd-0.02629385766201261, 32'sd0.00936437931357513, 32'sd-0.11534482074205815, 32'sd0.014249682060335684, 32'sd0.07824043212356044, 32'sd0.09568313371394022, 32'sd-0.0366852703724825, 32'sd0.049232092236240615, 32'sd-0.007440934154706071, 32'sd-0.0993279934732302, 32'sd-0.02734495880942291, 32'sd-0.04931698313808685, 32'sd0.10496745956534913, 32'sd-0.046251542076373324, 32'sd0.028504202379937914, 32'sd0.06210468363885623, 32'sd-0.07067636841953813, 32'sd0.012324397139859604, 32'sd-0.08447471360254737, 32'sd0.043138987957374544, 32'sd0.030322504600695133, 32'sd-0.10045295844650126, 32'sd-0.19211657213942301, 32'sd-0.08771982400680742, 32'sd-0.06924756129993107, 32'sd0.06670205478303987, 32'sd0.03667843650994003, 32'sd0.11635625091384048, 32'sd0.16073288782413114, 32'sd0.1274903986941495, 32'sd0.05179819018180228, 32'sd0.028321485219773502, 32'sd0.040618422390209116, 32'sd0.11389555623096843, 32'sd0.1285381621476193, 32'sd0.004970268478663556, 32'sd0.02549273693542687, 32'sd0.025048919489534454, 32'sd-0.07923072598363835, 32'sd-0.0240720561136211, 32'sd0.09130897959318496, 32'sd0.05577892250042304, 32'sd0.0067895537922785494, 32'sd-0.015577118757863386, 32'sd0.024129807292987044, 32'sd0.03212799680314701, 32'sd-0.04992985557628947, 32'sd-0.031894378541569644, 32'sd0.07304461167452118, 32'sd-0.0040112324487023504, 32'sd-0.07627672052365674, 32'sd-0.013732319277150599, 32'sd0.0029752036617177705, 32'sd-0.06265543574141615, 32'sd0.06310478135177301, 32'sd0.17714067130424194, 32'sd0.24010420742170005, 32'sd0.09578485269122938, 32'sd0.06270738477112323, 32'sd0.038526008120086636, 32'sd0.17324456535296082, 32'sd0.19346628949463074, 32'sd0.08266700569199693, 32'sd-0.02575656687878968, 32'sd-0.027901922433791707, 32'sd-0.10929298939890626, 32'sd0.005884376702858947, 32'sd0.026286046441420043, 32'sd0.08567118248003149, 32'sd-0.10269164875424161, 32'sd-4.1920145006565026e-123, 32'sd0.020369754007330487, 32'sd-0.11179560546273984, 32'sd0.07561665157700925, 32'sd0.01911112046390728, 32'sd-0.027278121776939095, 32'sd0.003063193733063037, 32'sd-0.0868027509142671, 32'sd-0.01376794523958134, 32'sd0.08313412874346048, 32'sd-0.0298795136698551, 32'sd0.03616696296735729, 32'sd0.15165173965761283, 32'sd0.16704437114919837, 32'sd0.1326026091814823, 32'sd-0.00025737649485514186, 32'sd-0.023092784996304683, 32'sd0.01007573350607279, 32'sd0.1367801422492076, 32'sd0.09493490855619596, 32'sd0.03648051923853861, 32'sd-0.12641028375780688, 32'sd-0.06231781260822832, 32'sd-0.1375799150488984, 32'sd-0.1400039334932499, 32'sd-0.10376805706123433, 32'sd-0.06640622844690706, 32'sd-0.02095786519085291, 32'sd0.0641172032757549, 32'sd-0.06342589759302099, 32'sd0.021477099130150244, 32'sd0.03989924871872728, 32'sd-0.03869390591067495, 32'sd0.013806127848273918, 32'sd0.01518563452561375, 32'sd0.20290350874920915, 32'sd0.04345879716796608, 32'sd-0.035437960692341, 32'sd0.036984922725919384, 32'sd0.08345817389608134, 32'sd-0.0372686306979598, 32'sd0.09073487309797665, 32'sd0.10961471730030202, 32'sd-0.04236270348661386, 32'sd0.018199463945899698, 32'sd0.2145731218242881, 32'sd0.10040015141037907, 32'sd0.19506899409450737, 32'sd0.004876789777660978, 32'sd-0.06275043820554646, 32'sd-0.038885751583570105, 32'sd-0.06992289444119858, 32'sd-0.05210110829671035, 32'sd-0.11030594985710594, 32'sd-0.037392108872274794, 32'sd0.08625977814276657, 32'sd0.003422164907686134, 32'sd0.05838230169086196, 32'sd-0.1354884158284024, 32'sd-0.07893723864542018, 32'sd0.18934023284724275, 32'sd0.13767748386106457, 32'sd0.050692766024000156, 32'sd0.13618292731536846, 32'sd0.13792276193903982, 32'sd-0.05378100201490741, 32'sd-0.0417263187789649, 32'sd0.046063867799064004, 32'sd-0.06266062179659289, 32'sd-0.14284746785478739, 32'sd-0.0214392492890465, 32'sd0.03480438775484425, 32'sd0.17204398329018475, 32'sd0.015101410468619753, 32'sd0.0017862325567994065, 32'sd0.06345804147975356, 32'sd-0.10390432728214877, 32'sd0.04189529712530015, 32'sd0.04189778696850992, 32'sd-0.01944750549807159, 32'sd-0.046729411457783664, 32'sd-0.23318567867873202, 32'sd0.09813340810109514, 32'sd-0.01555174400803553, 32'sd-7.208626523151216e-120, 32'sd-0.015360987779318706, 32'sd-0.05082154678715115, 32'sd0.04275075088350262, 32'sd0.18092275346004308, 32'sd0.10084744078952179, 32'sd0.022263573318771893, 32'sd0.07407180303491603, 32'sd0.06465509321717473, 32'sd-0.01348448957550151, 32'sd0.060313787714541364, 32'sd-0.1372366930210175, 32'sd-0.16402174234455766, 32'sd-0.15729974149166348, 32'sd0.005935084839788536, 32'sd0.01572014559356298, 32'sd0.05054522654247814, 32'sd-0.14759577047623518, 32'sd0.001211292544439206, 32'sd-0.02479707470796579, 32'sd-0.062243216161752414, 32'sd-0.10098816268445145, 32'sd-0.07838281704083529, 32'sd-0.059993001619531514, 32'sd-0.006236678420010834, 32'sd-0.15503274055096355, 32'sd0.09191891610233215, 32'sd0.03927066772060603, 32'sd-0.03220599024313742, 32'sd0.00398643730207187, 32'sd0.01648037774670815, 32'sd0.15968403810115855, 32'sd0.02238702533236272, 32'sd0.08674007747644635, 32'sd0.006721746454425098, 32'sd0.060086321420612696, 32'sd0.02143638409555483, 32'sd-0.12582022391906397, 32'sd0.012264835730617046, 32'sd-0.12618268893384754, 32'sd-0.09225726192168782, 32'sd-0.15170542848344828, 32'sd0.020322275217937, 32'sd-0.1329597824300031, 32'sd-0.018931220411731994, 32'sd-0.0686947632948776, 32'sd0.018715061265317173, 32'sd-0.10733744180671767, 32'sd-0.16848909263712278, 32'sd-0.09004559203605575, 32'sd-0.06375987839328602, 32'sd0.035954451933336844, 32'sd0.03341627891173017, 32'sd-0.006759600460637983, 32'sd0.05537918854534612, 32'sd0.08144210080842651, 32'sd-0.025710589112822518, 32'sd-0.004847381480853569, 32'sd0.06356765730954611, 32'sd0.01792973197365957, 32'sd0.006646534039731957, 32'sd-0.041146693686478546, 32'sd-0.1460243782313577, 32'sd-0.12255266671027334, 32'sd-0.03498006919070424, 32'sd-0.12151794568807504, 32'sd-0.05297535549047085, 32'sd-0.15514924968218385, 32'sd-0.03527373894103574, 32'sd-0.14863715832268165, 32'sd-0.1557221986406682, 32'sd0.016376988269115867, 32'sd0.03369079786000648, 32'sd0.019856325440419927, 32'sd0.03930921044103532, 32'sd0.019562340925585918, 32'sd-0.06006867577101178, 32'sd-0.10413192597861404, 32'sd-0.10687109002241973, 32'sd0.047519047533103445, 32'sd0.010654864689996314, 32'sd-0.006463293514432663, 32'sd-0.08981388880701033, 32'sd0.009778106462996669, 32'sd4.53889340245593e-127, 32'sd-0.0003312807547187147, 32'sd0.021536409279338642, 32'sd-0.026745760724703603, 32'sd-0.04222685338177324, 32'sd-0.043268849956419705, 32'sd-0.025956287950368813, 32'sd-0.1252590111028053, 32'sd-0.10357994240877663, 32'sd-0.030212028428345382, 32'sd-0.06204665698452442, 32'sd-0.003453328585224384, 32'sd-0.00984629339973886, 32'sd-0.005310231875473331, 32'sd-0.019618754855835564, 32'sd-0.01648273956113538, 32'sd0.0049509156220754235, 32'sd-0.000762459047831209, 32'sd0.05026252217700084, 32'sd-0.009066305472825303, 32'sd-0.02042050174067226, 32'sd-0.08008246076416753, 32'sd-0.054052053114586614, 32'sd0.054738906938721715, 32'sd0.10161575314584863, 32'sd-0.014960703633997588, 32'sd-0.08342395090554, 32'sd-2.7774003305335127e-123, 32'sd2.149570169271882e-116, 32'sd-1.3766281537141097e-121, 32'sd0.08489301100667596, 32'sd-0.020218923094191765, 32'sd0.0443659542291778, 32'sd-0.02386872439505464, 32'sd-0.05790404930038176, 32'sd-0.06843958714758128, 32'sd-0.0124375246342145, 32'sd0.014019292432517387, 32'sd-0.007971216244447672, 32'sd0.014393598856060863, 32'sd0.000323582876148755, 32'sd-0.07582038458424027, 32'sd-0.0009734834133604273, 32'sd-0.06115234541964925, 32'sd-0.07848076659966875, 32'sd0.0456105712039072, 32'sd-0.07098651394399395, 32'sd-0.02291748500478083, 32'sd0.11943203511626514, 32'sd0.06604910466187454, 32'sd-0.03591651872028462, 32'sd-0.05249420315032571, 32'sd0.07476016409143088, 32'sd-0.0550849723421265, 32'sd0.05455743655281146, 32'sd-5.9392228776166175e-121, 32'sd-1.6032917234068218e-119, 32'sd2.2164841026401412e-125, 32'sd-0.040395579802966076, 32'sd0.017706472194147272, 32'sd-0.053789634270582025, 32'sd-0.012892826016733498, 32'sd-0.12392874445271253, 32'sd-0.01649272111459904, 32'sd-0.04502706774012576, 32'sd0.11819847574368343, 32'sd-0.008863188034527042, 32'sd-0.12357420581647689, 32'sd0.016516155732954365, 32'sd-0.046704919266012376, 32'sd-0.07817106792908, 32'sd-0.10924641229055301, 32'sd0.08961308016787045, 32'sd-0.02457542089573971, 32'sd-0.040307203849545656, 32'sd0.09226747891502692, 32'sd0.02008241930357953, 32'sd-0.03166922494489422, 32'sd-0.022117077659318557, 32'sd-0.014302382292633453, 32'sd-0.05044129767010629, 32'sd-0.043114062563387255, 32'sd0.04546113449540948, 32'sd-3.086982664165136e-126, 32'sd1.4362346087616438e-118, 32'sd2.5852763143026956e-126, 32'sd4.869145858149673e-124, 32'sd0.00037365445933859473, 32'sd-0.07744620882941922, 32'sd-0.012134653486340451, 32'sd0.017175217249440426, 32'sd0.06714974443105903, 32'sd0.04134717389577401, 32'sd0.03596429289271581, 32'sd-0.0477696536299145, 32'sd-0.011318780160969738, 32'sd0.017945258602807254, 32'sd0.002382980882635842, 32'sd0.03926261728442205, 32'sd-0.09582816639799, 32'sd0.020843910129892305, 32'sd-0.012456308488415741, 32'sd-0.04664287331372956, 32'sd0.05382960238369878, 32'sd0.09223160913106765, 32'sd0.06750775708695345, 32'sd0.0027171713198147268, 32'sd-0.05872491198197224, 32'sd-0.00876188446893101, 32'sd-0.002043964971224788, 32'sd8.611664381415907e-117, 32'sd-1.4694425680398913e-121, 32'sd-3.7542252239171136e-119, 32'sd8.572097180340232e-117, 32'sd3.357631292260597e-124, 32'sd-1.8669976633219757e-127, 32'sd0.018334722911660432, 32'sd-0.014144090745849394, 32'sd-0.0005374422133851637, 32'sd0.12233533218344977, 32'sd0.006907736081502278, 32'sd0.05055622899102391, 32'sd0.029088592143827814, 32'sd0.04996096511201763, 32'sd0.051661882325722, 32'sd-0.00893480324142705, 32'sd0.11203763555054737, 32'sd0.026297552194751005, 32'sd0.07336185221564023, 32'sd-0.006077452077546535, 32'sd0.0215485599682858, 32'sd0.1324932706401678, 32'sd0.020830162437451404, 32'sd0.03524250909155845, 32'sd-0.06039437577848424, 32'sd0.021398919459417035, 32'sd-1.2744965820689879e-125, 32'sd-1.6626976593283286e-121, 32'sd-2.420278418129188e-125, 32'sd1.0110257645291184e-128},
        '{32'sd1.8526740373928363e-119, 32'sd1.5147030966176966e-120, 32'sd-6.686489879403961e-122, 32'sd-2.4864295890228243e-120, 32'sd9.136133319543934e-128, 32'sd7.850837955208712e-119, 32'sd-1.282334365432715e-122, 32'sd-2.8554184941821223e-127, 32'sd-3.7385160491599015e-123, 32'sd-4.218568365326489e-124, 32'sd-7.542472051998174e-126, 32'sd-1.3324363394139711e-126, 32'sd0.0540879886946106, 32'sd0.027807676983603542, 32'sd0.08163245432737194, 32'sd0.13011112673683028, 32'sd-5.385438174436746e-119, 32'sd-3.457718117982125e-114, 32'sd1.05064993282542e-124, 32'sd6.799202232722328e-126, 32'sd2.7293490068655044e-114, 32'sd3.1882804613875793e-128, 32'sd1.8476890491687628e-117, 32'sd-4.854978625143705e-115, 32'sd-9.637253545995231e-121, 32'sd4.328372799443397e-125, 32'sd-5.432035388543894e-125, 32'sd9.846329943470504e-128, 32'sd-1.0812019112591353e-125, 32'sd5.090114182675354e-124, 32'sd3.362310816794531e-119, 32'sd-1.3453396286898521e-123, 32'sd-0.037915233193697294, 32'sd0.037516498573270184, 32'sd-0.0039533243828873185, 32'sd0.0666682684225456, 32'sd-0.09144288805372773, 32'sd0.013942953116409584, 32'sd0.05312528747494357, 32'sd0.024724365554485202, 32'sd0.009685589624591002, 32'sd-0.03524071455811132, 32'sd0.06703458220207768, 32'sd0.06897146091513753, 32'sd-0.013689985219314941, 32'sd0.02000719516342895, 32'sd0.0035037916684212255, 32'sd-0.042570145700799235, 32'sd0.03482177736674562, 32'sd0.031504417114490244, 32'sd0.049486302996972945, 32'sd0.07191047484251256, 32'sd1.0883328792620212e-122, 32'sd1.5420247635958536e-120, 32'sd2.5972647578866078e-126, 32'sd3.9597447245141644e-116, 32'sd-4.069198690544048e-116, 32'sd-4.013950637302691e-127, 32'sd0.07422492461077536, 32'sd0.011256954803596507, 32'sd-0.02538530837901131, 32'sd-0.00855353152901124, 32'sd-0.010986156411801036, 32'sd-0.05301910702953396, 32'sd-0.06518360094265409, 32'sd-0.0577815854222036, 32'sd-0.09746654089551623, 32'sd0.04908023564134113, 32'sd0.02569194847694219, 32'sd0.16587409792811028, 32'sd0.02402825827530934, 32'sd0.12680721916325058, 32'sd0.059518994283701686, 32'sd0.04387267431985554, 32'sd0.0682061271139961, 32'sd0.11927286035204009, 32'sd0.097015120551198, 32'sd0.036162043310623844, 32'sd-0.021230171197137434, 32'sd0.024068272094594837, 32'sd0.07947180289419153, 32'sd0.09790618847761304, 32'sd-6.798496323786102e-115, 32'sd2.8622663111979595e-116, 32'sd1.4067321435652983e-115, 32'sd-1.2622644734115958e-121, 32'sd0.09429062935984016, 32'sd-0.025488200895253586, 32'sd0.055810542396565015, 32'sd0.10158284852118524, 32'sd0.004542181732424388, 32'sd0.021615546158705073, 32'sd0.10113186011970243, 32'sd0.11332091498821176, 32'sd0.14268218626870152, 32'sd0.0025250837623650314, 32'sd-0.03257267953964833, 32'sd0.030009596164413642, 32'sd0.041458531960480695, 32'sd-0.038864777256324416, 32'sd0.1500969944699515, 32'sd0.006288127618427274, 32'sd0.0882475763322953, 32'sd-0.07137557734561278, 32'sd0.018235019961122857, 32'sd0.05031755568152641, 32'sd-0.024365507946062494, 32'sd-0.05401622366953932, 32'sd0.06164055070269669, 32'sd-0.0003278943109075362, 32'sd-0.018142288016945222, 32'sd-4.328115446941737e-124, 32'sd1.4194859836312153e-115, 32'sd0.045237513816537324, 32'sd0.05915529030555599, 32'sd0.09467090433653905, 32'sd0.015710671355078493, 32'sd0.0355609038935355, 32'sd0.10598804892365407, 32'sd0.10516826396729737, 32'sd-0.008457842167063533, 32'sd0.11925138477006887, 32'sd0.0011754250595300132, 32'sd0.10003550335317461, 32'sd0.1384997778412615, 32'sd0.057985428830457555, 32'sd-0.015822625745433607, 32'sd-0.004665273908349452, 32'sd-0.011549306008199244, 32'sd-0.08949019476717178, 32'sd0.0030356974692286372, 32'sd-0.055117231974532666, 32'sd-0.07034124640662362, 32'sd-0.03867320773062922, 32'sd0.08462964909321333, 32'sd0.12367557926450197, 32'sd0.082305020114643, 32'sd-0.030987710856704237, 32'sd0.06463458145248124, 32'sd0.07992766302279217, 32'sd6.780369267303927e-126, 32'sd0.11015665913664052, 32'sd0.015474594222923854, 32'sd0.09441728055667627, 32'sd-0.09930767901617042, 32'sd0.01883028274731723, 32'sd-0.07812437093423188, 32'sd0.07775439011046158, 32'sd-0.062058555333238494, 32'sd-0.06969531553043674, 32'sd0.025058050689102048, 32'sd-0.0321279808522128, 32'sd0.05861395972898421, 32'sd-0.11914488111805642, 32'sd-0.03820351850491495, 32'sd-0.029122763378837478, 32'sd-0.0343856488924614, 32'sd-0.10525475928695262, 32'sd0.10686452019164695, 32'sd-0.008746728656718215, 32'sd-0.11056900588255111, 32'sd0.028901042767283884, 32'sd-0.034207678602781344, 32'sd-0.006810839357795086, 32'sd-0.009213220979232174, 32'sd0.002047060136064564, 32'sd0.07782961217747254, 32'sd-0.018539415770651282, 32'sd-8.539978267957986e-122, 32'sd0.0648948246690627, 32'sd0.0038205817808266603, 32'sd0.008277718939156208, 32'sd-0.05983539388603312, 32'sd-0.011203963776873271, 32'sd-0.10876789126851649, 32'sd-0.11136977162367367, 32'sd-0.0036210407783827587, 32'sd-0.04245261043455501, 32'sd-0.056780504596656886, 32'sd-0.006763235914615919, 32'sd0.05735692850573861, 32'sd-0.055158370920648916, 32'sd-0.005543769321589245, 32'sd0.045983652051370255, 32'sd-0.046975546674432676, 32'sd0.0268541823298198, 32'sd-0.04095444361870235, 32'sd-0.05730512537604417, 32'sd-0.12772916010415966, 32'sd0.024297003598404802, 32'sd-0.06485920904564244, 32'sd-0.09002000262690348, 32'sd0.05138547567049649, 32'sd-0.007163224759880296, 32'sd0.05560267266738116, 32'sd-0.02059131484496797, 32'sd0.08533986453638102, 32'sd-0.05846109398157603, 32'sd-0.023698443277037764, 32'sd0.024323638736600785, 32'sd-0.05109723691674497, 32'sd-0.0798957363818374, 32'sd0.01588383597967224, 32'sd-0.003698651551489781, 32'sd-0.03332967401710521, 32'sd-0.018869671307729888, 32'sd0.02004650249778596, 32'sd0.03661018177931028, 32'sd0.0037212979289899897, 32'sd0.18124006710244667, 32'sd0.07391770168708275, 32'sd0.12419892639268221, 32'sd0.05196340050825809, 32'sd-0.011019202632633101, 32'sd0.041833329967058644, 32'sd-0.044074046776060964, 32'sd-0.04031484487972549, 32'sd-0.14774912450069685, 32'sd-0.16035686972432367, 32'sd0.003726970412685375, 32'sd0.006488605568792283, 32'sd-0.09937573158304831, 32'sd0.035199798336209585, 32'sd-0.0011546023516068693, 32'sd0.08116279374593811, 32'sd0.01223389535229449, 32'sd-0.03063889231729722, 32'sd0.01819076761426476, 32'sd-0.10749529865658118, 32'sd-0.07898101207604612, 32'sd-0.042017057580287856, 32'sd-0.005456829609009149, 32'sd0.03655548717709179, 32'sd0.003052930233801135, 32'sd-0.007658567421602499, 32'sd0.021082879911923664, 32'sd0.13605944971526934, 32'sd0.15786061998129985, 32'sd0.14438004579807331, 32'sd0.15527464936796762, 32'sd0.01849115200481172, 32'sd0.12290260718967704, 32'sd0.11696069827513512, 32'sd0.12125397790432813, 32'sd-0.007098924774495875, 32'sd-0.017252437858872677, 32'sd0.01203600004567819, 32'sd-0.009277003893082785, 32'sd-0.038268278044180086, 32'sd0.0253868625002123, 32'sd-0.07574143103689024, 32'sd0.04912733333650719, 32'sd0.0027412051644006255, 32'sd0.06798958595354085, 32'sd0.057087990951981714, 32'sd-0.035270606789376775, 32'sd-0.12078344603775677, 32'sd-0.11789687261654597, 32'sd0.08347114894395052, 32'sd0.008120590574519328, 32'sd-0.02958337087256503, 32'sd0.03394470593683377, 32'sd0.006610170916363265, 32'sd0.020138615190414908, 32'sd0.062322218286822044, 32'sd0.11228830652386569, 32'sd0.08981351947027351, 32'sd0.0801833268791084, 32'sd0.06705167701493892, 32'sd0.10791860604226272, 32'sd0.12471492231193648, 32'sd0.11125576302465205, 32'sd0.08093243076212822, 32'sd-0.17947395667946806, 32'sd-0.09989816904380609, 32'sd-0.0567399061244624, 32'sd0.03187344370964232, 32'sd0.05131720897174949, 32'sd0.04206971091932099, 32'sd0.006097935543495953, 32'sd0.0794395837408052, 32'sd-0.028452651654477665, 32'sd0.02000481949838031, 32'sd-0.06712632328839196, 32'sd-0.1375829323744797, 32'sd-0.022580029361366244, 32'sd0.033075881245797585, 32'sd0.0461986969868291, 32'sd0.09495981405531922, 32'sd0.05678109470564885, 32'sd0.02885171902549805, 32'sd-0.00037668887161986436, 32'sd-0.012040454975767213, 32'sd0.1374421683486329, 32'sd0.1515911620378185, 32'sd0.29062793738229414, 32'sd0.14881723879107722, 32'sd0.1300700098974638, 32'sd0.046417316334766125, 32'sd0.12174104825190166, 32'sd0.16973608300087115, 32'sd-0.12017155078629257, 32'sd0.0953947819472236, 32'sd0.07774578358673605, 32'sd-0.08736997301444328, 32'sd0.07594176603592447, 32'sd-0.10072682749809729, 32'sd0.03623484318875502, 32'sd0.08108986205658861, 32'sd0.11870035117992286, 32'sd0.020578657347150003, 32'sd0.16004592758784755, 32'sd0.031233919849305992, 32'sd-0.04865358386286774, 32'sd0.10965066966633467, 32'sd0.03884893089926904, 32'sd0.047918161206432025, 32'sd0.02658389242245989, 32'sd0.022188336741713433, 32'sd0.01786014254528557, 32'sd0.03348037627600994, 32'sd-0.06308865706002265, 32'sd0.04812326251246821, 32'sd0.14564778774806098, 32'sd-0.030663619872345633, 32'sd0.06587800274885675, 32'sd0.19321265979871216, 32'sd0.026738411698322615, 32'sd0.21744091703624763, 32'sd0.03531200376712413, 32'sd0.08093593590929862, 32'sd-0.020432273568327053, 32'sd-0.0805482818220243, 32'sd0.09094206215021712, 32'sd0.04321255595853869, 32'sd0.02374325407734529, 32'sd0.03999239237755803, 32'sd0.00787076048169065, 32'sd0.03046063124111726, 32'sd0.07516972439849733, 32'sd0.05490134316575234, 32'sd0.006712924485353382, 32'sd0.010664361724605172, 32'sd-0.07759050305990298, 32'sd-0.057861439007999574, 32'sd0.04280271359023615, 32'sd-0.10357741494864427, 32'sd-0.11530240232527716, 32'sd-0.11628905957192559, 32'sd-0.09964642514503151, 32'sd0.02225643691811595, 32'sd0.013418066072868363, 32'sd0.12138548849644726, 32'sd0.016523395845153076, 32'sd0.17876488026334691, 32'sd0.10563294241773383, 32'sd0.15803500630932713, 32'sd0.004233675530387992, 32'sd-0.0516114691888391, 32'sd-0.04483325641530896, 32'sd0.0066599682341417325, 32'sd-0.009741950381319359, 32'sd-0.017460623631994833, 32'sd-0.047504302536158255, 32'sd0.052209083327771896, 32'sd-0.043225968258353, 32'sd0.010394452086729584, 32'sd0.055818475783178854, 32'sd0.05653282101369332, 32'sd-0.09392277479833874, 32'sd0.05628655162704425, 32'sd-0.08024146346550466, 32'sd0.04020145143866484, 32'sd-0.04217835113410892, 32'sd-0.17508140965542976, 32'sd-0.10220274892611601, 32'sd-0.12140161753200737, 32'sd-0.12879004432961094, 32'sd-0.004610426502367219, 32'sd0.039795924527148065, 32'sd0.011410883958022467, 32'sd0.05721916489522269, 32'sd0.09837224666930378, 32'sd0.11271782128393446, 32'sd0.14575829218320155, 32'sd0.05839085040560672, 32'sd-0.0638825370028747, 32'sd-0.14451951064206675, 32'sd-0.09986777356579392, 32'sd-0.043873825942796325, 32'sd-0.000702187003376776, 32'sd-0.003345261159021883, 32'sd0.030746736395413737, 32'sd0.08986770677193655, 32'sd0.06697522212283981, 32'sd-0.0063133713032563965, 32'sd-0.036248100564877685, 32'sd0.00039889479744146145, 32'sd0.0734106749964536, 32'sd-0.06062776113302864, 32'sd0.030112240253978077, 32'sd-0.025141638989496163, 32'sd-0.08697514006948083, 32'sd-0.1270383434169321, 32'sd-0.148549020762797, 32'sd-0.20097682843947323, 32'sd-0.09739786075746901, 32'sd-0.031925360085496596, 32'sd0.048017911332778114, 32'sd-0.013825730669307335, 32'sd0.126386650101842, 32'sd-0.001480581632594998, 32'sd0.12105762389874825, 32'sd0.03829266437099831, 32'sd-0.048390618077537334, 32'sd-0.010430912211038318, 32'sd-0.04124598732434613, 32'sd0.028648599218986277, 32'sd0.06595779505046698, 32'sd-0.05545662796789823, 32'sd0.023732828417220343, 32'sd-0.0013621091020820126, 32'sd-0.10439297090785703, 32'sd-0.09525804364518725, 32'sd0.03394657774220856, 32'sd-0.026321267981709674, 32'sd-0.030173089189670335, 32'sd-0.10866237080729492, 32'sd-0.05574093564909284, 32'sd-0.04657637115125194, 32'sd-0.1460454904590412, 32'sd-0.14665130280366248, 32'sd-0.1351360682929434, 32'sd-0.04426764383037089, 32'sd-0.08861235826581114, 32'sd-0.08099784899127013, 32'sd-0.07159465918425975, 32'sd-0.018836697792437032, 32'sd-0.029942737078403173, 32'sd0.028209969213828345, 32'sd0.10235734210438972, 32'sd0.1036570814604399, 32'sd0.0036636100048067738, 32'sd0.117654626439796, 32'sd0.05339960763901103, 32'sd0.021224525187750164, 32'sd-0.05195549641039057, 32'sd0.04868652530010303, 32'sd0.05225057739210593, 32'sd0.03739184132513487, 32'sd-0.10282319925439412, 32'sd0.020733628867580973, 32'sd0.07120675715404179, 32'sd0.09682718777187228, 32'sd-0.05208048488815793, 32'sd-0.040874794595471296, 32'sd-0.05064060486404911, 32'sd-0.05607530267642168, 32'sd-0.0703799686674996, 32'sd-0.0672080426688315, 32'sd0.005803584429409557, 32'sd-0.11967978264473537, 32'sd-0.03669111154759277, 32'sd-0.07227978901192723, 32'sd0.028343118530507135, 32'sd0.04600167068186802, 32'sd-0.012716357657338357, 32'sd-0.08003810378030093, 32'sd-0.024900820415572164, 32'sd-0.014360338864605375, 32'sd-0.0857403745465095, 32'sd-0.014145157096088448, 32'sd0.11980418956079808, 32'sd-0.05213930268549733, 32'sd-0.0677761752514394, 32'sd0.02036249736106397, 32'sd-5.435265887074544e-121, 32'sd-0.03505280716909276, 32'sd-0.02515522937711314, 32'sd0.044490745519692836, 32'sd0.06678387095879978, 32'sd0.014310535147712584, 32'sd-0.020341748011485968, 32'sd-0.050539881233251614, 32'sd-0.04295884285708299, 32'sd-0.03950453888419938, 32'sd0.011931840551728853, 32'sd-0.0538433601207243, 32'sd-0.006605774393511771, 32'sd-0.028098949022667238, 32'sd-0.06403363534160633, 32'sd-0.10626832138189278, 32'sd-0.10471015278803007, 32'sd0.024526693181349812, 32'sd0.12283423348921332, 32'sd0.06494283728529747, 32'sd0.005493002349817773, 32'sd0.057302873624756306, 32'sd0.021548536370298275, 32'sd-0.10164767551105976, 32'sd0.029016827903183034, 32'sd0.021777680106298568, 32'sd-0.018119742065426502, 32'sd0.0169339192701915, 32'sd-0.010790833920506414, 32'sd0.021515782009841417, 32'sd0.0036101637852514698, 32'sd0.0538423685389017, 32'sd-0.005829635030454457, 32'sd-0.008601992344451567, 32'sd0.05411198268007164, 32'sd-0.0571865764254152, 32'sd-0.06974716443011993, 32'sd-0.1270099650621268, 32'sd0.05262200881252087, 32'sd-0.02091767268749629, 32'sd-0.016206241393395365, 32'sd-0.04467588567286131, 32'sd-0.10552750278073755, 32'sd-0.11967557661248304, 32'sd-0.09754749580743083, 32'sd0.1250629003915233, 32'sd0.0754840460729991, 32'sd0.03174595358177266, 32'sd0.053625170563460875, 32'sd0.049170577966332875, 32'sd0.07684581627247353, 32'sd-0.11339175262650238, 32'sd-0.056158826639449315, 32'sd0.008046473174380626, 32'sd-0.056418019836644004, 32'sd0.09113156757909358, 32'sd0.051246974465694164, 32'sd-0.07119439197435476, 32'sd-0.0203171704769923, 32'sd-0.007284179420041008, 32'sd0.02208225786982837, 32'sd0.02486697679233438, 32'sd-0.11747573339451632, 32'sd-0.01204273300556915, 32'sd-0.09024451620043272, 32'sd-0.03635782423026993, 32'sd-0.028972413168111916, 32'sd-0.05715457740201362, 32'sd0.01691918250367088, 32'sd-0.12810411201442135, 32'sd-0.028217603518424356, 32'sd0.0026645278436611317, 32'sd-0.052726508569717695, 32'sd0.03805999891502212, 32'sd0.12044043387636003, 32'sd0.17160518518094559, 32'sd0.14383433495667136, 32'sd0.006509855219363551, 32'sd-0.01899721080474056, 32'sd-0.2238865512582177, 32'sd0.016033168512440823, 32'sd0.009543194536428516, 32'sd-0.0776959900685935, 32'sd0.04552704421371408, 32'sd1.9483958290807104e-124, 32'sd0.045033164982876565, 32'sd0.005619644576208963, 32'sd-0.11159442422017679, 32'sd0.0056900983802477875, 32'sd-0.0032318641697841213, 32'sd-0.07542768488934423, 32'sd-0.06231132407311891, 32'sd-0.006200186604860375, 32'sd-0.07404635694454037, 32'sd-0.113060560390763, 32'sd-0.011795790475361547, 32'sd-0.09479754712265749, 32'sd-0.024809553332687827, 32'sd0.014321983385714776, 32'sd0.022992437251608776, 32'sd0.061717349128127444, 32'sd0.11955381141392314, 32'sd0.014072799874863791, 32'sd0.041139935839731766, 32'sd-0.019290279515626573, 32'sd-0.12600839060593366, 32'sd-0.08069662463124222, 32'sd-0.08035870341834199, 32'sd-0.11424650076503905, 32'sd0.07649024769871966, 32'sd0.0859521350742955, 32'sd0.059495858097002745, 32'sd0.08446660719579416, 32'sd0.020140529141173532, 32'sd-0.01810859781307061, 32'sd0.0159554394354579, 32'sd-0.04824647116890148, 32'sd0.021619755495781955, 32'sd-0.04170424665679968, 32'sd0.04335351650188495, 32'sd-0.10201419593222114, 32'sd0.024000614949137425, 32'sd-0.0711124231096787, 32'sd-0.03249846153845699, 32'sd0.017406301755559593, 32'sd0.053694516567194074, 32'sd-0.025034366823471068, 32'sd-0.004131315822772959, 32'sd0.07401799467457967, 32'sd0.021264147101184582, 32'sd0.03701816062320936, 32'sd-0.041943833264663166, 32'sd0.03963335925143487, 32'sd-0.08711387014886075, 32'sd-0.05648499819008497, 32'sd-0.01856222026173276, 32'sd-0.07110850697444922, 32'sd0.09629278996041084, 32'sd0.02656053360862159, 32'sd0.0832718497190776, 32'sd0.11715972038440646, 32'sd-0.019893566926535038, 32'sd0.0850504806293918, 32'sd0.01455624995655277, 32'sd0.08198727450895539, 32'sd0.09535100509606866, 32'sd0.04791040297957374, 32'sd0.0016071837361361343, 32'sd-0.014893564354640744, 32'sd0.02594147240550132, 32'sd-0.017425762513301236, 32'sd0.14509681070708083, 32'sd0.0921348305651186, 32'sd0.08786281170019036, 32'sd0.12392511063208655, 32'sd-0.01502385050887004, 32'sd-0.011559947512305352, 32'sd0.010531247355147778, 32'sd-0.03312325551525147, 32'sd0.08805082951570213, 32'sd-0.0819000494270249, 32'sd-0.10886785021227476, 32'sd-0.08417513754372104, 32'sd-0.038503069381845, 32'sd-0.01583762317437552, 32'sd0.02656072839895851, 32'sd-0.011691306970938616, 32'sd0.030493583486868005, 32'sd-1.0877342575891748e-121, 32'sd0.07481360919313951, 32'sd-0.00871153656475951, 32'sd-0.028827320056028692, 32'sd-0.05891693213979427, 32'sd0.009497448229722318, 32'sd0.10141086528409529, 32'sd0.015191745557191858, 32'sd-0.018037740101668562, 32'sd-0.10324378163359842, 32'sd-0.02628746958139436, 32'sd0.0653750613772202, 32'sd-0.0005968134597848968, 32'sd0.020325429140901585, 32'sd0.07658865882160054, 32'sd0.11486696645607299, 32'sd0.02969715876752637, 32'sd0.0318451836788829, 32'sd0.06715223576756811, 32'sd0.053487516623215776, 32'sd-0.02671183267622579, 32'sd-0.03676412818772088, 32'sd-0.06254737723543215, 32'sd0.07435598043672802, 32'sd0.03847758042700465, 32'sd-0.016587262042302948, 32'sd0.06659221570812385, 32'sd-1.0403742864285135e-124, 32'sd1.0797909434350675e-117, 32'sd-2.0234663434394803e-117, 32'sd-0.03015173518863594, 32'sd0.0928599438152217, 32'sd-0.021036062914152658, 32'sd-0.025834967770887222, 32'sd0.03344457513274559, 32'sd0.010676847482237923, 32'sd0.04463861368514704, 32'sd0.12991794901130113, 32'sd0.049367186778104706, 32'sd0.009845609887148657, 32'sd0.019781790391328224, 32'sd0.0067174504588862856, 32'sd0.03626974189610072, 32'sd-0.06738559630646451, 32'sd-0.05211496610958331, 32'sd-0.02588101186169631, 32'sd0.019928607024007693, 32'sd-0.07870206560373323, 32'sd-0.0862028235170561, 32'sd-0.005002585974681786, 32'sd0.07471907989610299, 32'sd0.09824274671324058, 32'sd0.00037161828752456383, 32'sd0.029105536576351124, 32'sd-0.01845285788867982, 32'sd-1.3403821940052077e-122, 32'sd2.4588980229007546e-124, 32'sd-5.3747659658396606e-118, 32'sd0.07990290403758701, 32'sd0.10033816644928166, 32'sd0.04613522753545893, 32'sd0.019039302582194495, 32'sd-0.0178293866693576, 32'sd0.06819006529033557, 32'sd0.14886719376538599, 32'sd0.1165667034157124, 32'sd0.023465030978160176, 32'sd0.08299492201719193, 32'sd0.07026343677949211, 32'sd-0.06144050484886521, 32'sd0.17682906643901752, 32'sd-0.054547754270812245, 32'sd0.006086383633062838, 32'sd-0.017074373512090592, 32'sd0.05005926234504361, 32'sd-0.029379148488982473, 32'sd-0.07068099491213203, 32'sd-0.026320048858022624, 32'sd0.09321774917660128, 32'sd-0.05383729264758136, 32'sd0.08028922305602477, 32'sd0.032592225849902096, 32'sd-0.005464220822123941, 32'sd-3.7989905305262444e-122, 32'sd-9.851260970355385e-119, 32'sd3.395815559841424e-120, 32'sd-1.1478361354397767e-115, 32'sd0.11615944492032841, 32'sd0.05420584541186538, 32'sd-0.08505125524852258, 32'sd-0.09021176935978603, 32'sd0.020669326383147935, 32'sd-0.004071032047474949, 32'sd0.12591716499278066, 32'sd0.17947444409452207, 32'sd0.04873276013883843, 32'sd0.023450698672928125, 32'sd0.03631568733481002, 32'sd0.04722402868488121, 32'sd0.08866997430502734, 32'sd0.09831643399783763, 32'sd0.037861164462463695, 32'sd0.10047457099087083, 32'sd0.12463247203514251, 32'sd-0.037110597650961925, 32'sd-0.07762739110378623, 32'sd0.0659519918525369, 32'sd-0.02662933785927428, 32'sd0.02691742998293101, 32'sd0.059116281740704955, 32'sd-8.077115397437658e-119, 32'sd1.1078178094070049e-119, 32'sd-1.4902726143183727e-121, 32'sd4.0730824395934146e-125, 32'sd1.725376878200103e-117, 32'sd-1.8124335790804554e-126, 32'sd0.13938673489995157, 32'sd0.06789680599623789, 32'sd0.058095152707780144, 32'sd0.07340990135654292, 32'sd0.05497599632411944, 32'sd-0.0474085005898253, 32'sd0.12357058166136273, 32'sd0.025374953841892773, 32'sd0.06161872147494604, 32'sd-0.0070863902618241645, 32'sd0.07139672158986171, 32'sd0.11345118925873526, 32'sd0.04761980034343487, 32'sd0.042033240211834015, 32'sd-0.030236681363115102, 32'sd0.0697970751985652, 32'sd0.0829022401667917, 32'sd0.01160062200455461, 32'sd0.03380531966701835, 32'sd0.08007954177634194, 32'sd-2.6908748344047567e-129, 32'sd-3.5652748081855837e-122, 32'sd3.8911446042068827e-119, 32'sd1.48167033360453e-125},
        '{32'sd-5.217516573875417e-118, 32'sd-1.720827083883539e-125, 32'sd1.3551198870914572e-118, 32'sd1.7673359143798615e-123, 32'sd-1.663731856332069e-122, 32'sd-7.482513958099271e-115, 32'sd-2.1291834933807432e-126, 32'sd1.9533706916553868e-126, 32'sd-3.4328520670371285e-116, 32'sd-1.702826253220544e-125, 32'sd-4.840628746382608e-123, 32'sd-2.011443597738564e-117, 32'sd-0.10035012128335367, 32'sd0.0224178556269391, 32'sd-0.024723374290084553, 32'sd0.009372787018047814, 32'sd8.21687393331524e-126, 32'sd2.5155986668290515e-121, 32'sd-1.1932935712912242e-118, 32'sd-6.323597455982651e-125, 32'sd1.1849911232517884e-115, 32'sd4.086686287727158e-123, 32'sd-1.0062586572052853e-119, 32'sd9.390705324815846e-121, 32'sd8.339153460235514e-123, 32'sd9.761903838351692e-115, 32'sd2.1615708360559667e-120, 32'sd6.5876088517804475e-121, 32'sd-6.35904411199256e-120, 32'sd-1.5107155501185323e-115, 32'sd-3.0143782682486044e-118, 32'sd-6.439525570460676e-117, 32'sd-0.013105237905677504, 32'sd0.014919781950549962, 32'sd-0.05219092996734193, 32'sd0.021459166598534595, 32'sd-0.05704612470015093, 32'sd-0.043388194134339836, 32'sd-0.009756033132931432, 32'sd-0.0016521095989318797, 32'sd0.08042121037647489, 32'sd-0.11775253237340988, 32'sd-0.12375579685993049, 32'sd-0.11085494876847503, 32'sd-0.08459339709684212, 32'sd-0.10133837421302713, 32'sd0.015351629733035268, 32'sd-0.09188539266563216, 32'sd-0.0008349160604236398, 32'sd-0.0897737773580864, 32'sd-0.06994263546367012, 32'sd-0.060417432310082717, 32'sd-8.835881683660219e-127, 32'sd4.454168527489533e-118, 32'sd5.7531230799239505e-115, 32'sd9.805726659881516e-124, 32'sd7.457568415352501e-126, 32'sd-1.438628300874775e-115, 32'sd-0.058959374004163595, 32'sd-0.06704322799337342, 32'sd-0.09706176328557133, 32'sd-0.09485185959614009, 32'sd0.04226064034779094, 32'sd-0.05472529935460548, 32'sd0.05535552521180799, 32'sd0.019909802332113737, 32'sd0.08409639235130846, 32'sd-0.04748245154175441, 32'sd0.06960797809536236, 32'sd0.1166609660617135, 32'sd0.04779812105410053, 32'sd0.013177314570987378, 32'sd0.0347175855595036, 32'sd-0.07625938765808479, 32'sd-0.10147229354388941, 32'sd-0.019989363399139662, 32'sd-0.059112482397034954, 32'sd-0.033998950264227015, 32'sd0.023330716591385185, 32'sd-0.05935185057366491, 32'sd-0.02739047605824393, 32'sd0.023189102456743924, 32'sd1.3240959402379678e-127, 32'sd-3.5614998750663253e-118, 32'sd8.12974385888e-129, 32'sd1.0143741882573225e-121, 32'sd-0.05184535772589459, 32'sd0.027657870636260885, 32'sd-0.07138139794571056, 32'sd-0.13678906760697004, 32'sd0.032673825723440846, 32'sd-0.03951926330277931, 32'sd0.055722459949183505, 32'sd-0.03578496466533036, 32'sd0.11475623989325404, 32'sd0.022627486692165993, 32'sd0.03645904054801158, 32'sd0.1129264529239917, 32'sd-0.051228064010223444, 32'sd0.12821278728262087, 32'sd0.1714691503868212, 32'sd0.11509294301001285, 32'sd-0.0036968485344875974, 32'sd0.042117502926416216, 32'sd-0.000738139050385035, 32'sd0.041128444255587156, 32'sd-0.09846076259330132, 32'sd-0.01885592537987762, 32'sd-0.07857206812307954, 32'sd-0.10560336928128645, 32'sd-0.07892666292212715, 32'sd1.4350730354441245e-118, 32'sd-4.307438210192347e-115, 32'sd0.02574113371527086, 32'sd-0.07188120763263545, 32'sd-0.08854782915166584, 32'sd-0.07896216789454334, 32'sd0.02419085764445825, 32'sd0.10290362902945685, 32'sd0.01413917244804481, 32'sd0.05813725463585441, 32'sd0.16698391128205226, 32'sd-0.01791192621751713, 32'sd0.04818110457176955, 32'sd0.15505574038317635, 32'sd-0.0302011158498056, 32'sd0.05408518759575842, 32'sd-0.020205834347088867, 32'sd0.14530316273520957, 32'sd0.16168448942175612, 32'sd0.08801844755474653, 32'sd-0.019546123702589343, 32'sd0.0285654672486301, 32'sd-0.007190195223185081, 32'sd0.020575831137116238, 32'sd-0.03241232428857485, 32'sd-0.031643476441910914, 32'sd0.0215216897852485, 32'sd-0.017111797004146764, 32'sd0.048986190722811976, 32'sd-7.877007887606444e-121, 32'sd0.025830245010157, 32'sd-0.07800705448278507, 32'sd-0.05411559871774845, 32'sd-0.04638523707735565, 32'sd0.09752077362798342, 32'sd-0.032059918043400845, 32'sd0.13751993952521027, 32'sd-0.04509079430402277, 32'sd0.07063095687702557, 32'sd-0.041708130040534065, 32'sd0.08877375677979736, 32'sd0.14164891536434113, 32'sd0.13022257797237588, 32'sd0.10950925172352023, 32'sd0.025903395649398947, 32'sd0.023445002950978844, 32'sd0.05523039641565156, 32'sd-0.015591906372976933, 32'sd-0.04157260264005796, 32'sd0.06065395745885185, 32'sd0.17742213797977383, 32'sd-0.045788357722733555, 32'sd-0.046495747994879856, 32'sd-0.18918280009311686, 32'sd-0.03137885689761946, 32'sd0.010407276300989173, 32'sd0.06360510366602727, 32'sd-2.8829069644596513e-120, 32'sd-0.04889157096279657, 32'sd-0.033871275488267245, 32'sd-0.028896585117285392, 32'sd0.044245580675206155, 32'sd0.07810274289115521, 32'sd0.05049348633549886, 32'sd0.11340730213919531, 32'sd0.058551668902134715, 32'sd0.0056692755356736926, 32'sd0.026577007498133524, 32'sd0.04115639536238384, 32'sd0.10833857858558224, 32'sd0.01579216230048886, 32'sd0.09969573079818797, 32'sd-0.027586667274690838, 32'sd0.07489805260916484, 32'sd-0.02114399803780013, 32'sd0.06521191316767473, 32'sd0.059132587694436696, 32'sd0.0823484257891971, 32'sd0.15014110858669166, 32'sd0.05203345931515707, 32'sd-0.005460516061552802, 32'sd0.03422578718831798, 32'sd-0.023088367951381878, 32'sd-0.03775052712749392, 32'sd0.026569660225990062, 32'sd-0.0024646642477604407, 32'sd-0.07719610820354708, 32'sd0.009642896535429036, 32'sd-0.04378083004786384, 32'sd-0.012652268328867133, 32'sd-0.07792165419718174, 32'sd0.03109080615243958, 32'sd-0.056097384178082056, 32'sd7.114096246021454e-05, 32'sd0.10163025061587416, 32'sd0.06694523738288961, 32'sd0.13078980405383728, 32'sd0.12185373557117085, 32'sd0.1098335313017073, 32'sd0.11162448283785206, 32'sd0.037953107885825586, 32'sd-0.09633115311927737, 32'sd-0.02964097522589985, 32'sd0.07376289500743993, 32'sd0.1472415520779583, 32'sd0.025391044273495745, 32'sd-0.005261829681356871, 32'sd0.0982163790171785, 32'sd0.05962859009337217, 32'sd0.0211554842217721, 32'sd0.04767210369272934, 32'sd-0.08331084672567754, 32'sd-0.06004548684906634, 32'sd-0.030804840609074898, 32'sd0.04945063220707643, 32'sd0.041835832628725964, 32'sd-0.03927040895396485, 32'sd-0.05360741952430613, 32'sd-0.04177157163315142, 32'sd0.06420895974510164, 32'sd0.060807098783299394, 32'sd-0.03288817709859235, 32'sd0.04134875432050084, 32'sd0.11723180003421124, 32'sd0.20561725532560352, 32'sd0.15896492015574465, 32'sd0.10845793582979808, 32'sd-0.03529210586560569, 32'sd-0.047981161949218844, 32'sd-0.062278030137380085, 32'sd0.027978436309331528, 32'sd0.037506883575160015, 32'sd0.012344642629505395, 32'sd-0.05183180375797881, 32'sd-0.04366622807148547, 32'sd0.09561997677198084, 32'sd0.13998249061564735, 32'sd0.05784006620840217, 32'sd0.013407429539040968, 32'sd0.051835801214688705, 32'sd-0.04005182308946193, 32'sd0.09593708975095941, 32'sd0.11198493478675911, 32'sd-0.040833033201169745, 32'sd-0.13236518748447515, 32'sd-0.04470236313597636, 32'sd-0.09714388596355224, 32'sd-0.04763112404976776, 32'sd-0.11148773794226902, 32'sd-0.06673787376230457, 32'sd-0.032262844417701046, 32'sd0.08767369591863285, 32'sd0.14647903953479544, 32'sd0.16969506903411916, 32'sd0.1432922444800589, 32'sd0.09540012582480167, 32'sd0.07060385934187262, 32'sd-0.1315128614769193, 32'sd0.04272773481421892, 32'sd0.04077245941790182, 32'sd0.05946819088179685, 32'sd-0.03947210442975529, 32'sd0.00237238323112861, 32'sd-0.03551572891897485, 32'sd0.03841014705274221, 32'sd-0.015492339734431449, 32'sd0.03309200026180842, 32'sd0.004845603647319343, 32'sd-0.06787771870718122, 32'sd-0.008458621570064868, 32'sd0.053910873605769634, 32'sd-0.012340604769856234, 32'sd-0.07234581971723623, 32'sd-0.06748228977292595, 32'sd-0.07555806214137101, 32'sd-0.17302740451502227, 32'sd-0.11012183421359463, 32'sd-0.18731625544310446, 32'sd-0.14544598285842159, 32'sd-0.022463368520436497, 32'sd0.04987512027843106, 32'sd0.16262901203873012, 32'sd0.16492011736279252, 32'sd0.07481588331850349, 32'sd0.040187239444281195, 32'sd-0.051663392363234376, 32'sd0.040416031849801734, 32'sd0.11590472658091899, 32'sd-0.07503033940154705, 32'sd-0.03790109963124265, 32'sd-0.1331580474740333, 32'sd-0.16738117960853735, 32'sd-0.02745179194783069, 32'sd-0.1302497475539536, 32'sd-0.06821104386770112, 32'sd0.052779165616227725, 32'sd-0.015258137145773402, 32'sd0.025183011112976, 32'sd0.08960407834493324, 32'sd0.09867702714657191, 32'sd0.03390245650588362, 32'sd0.04637310652960781, 32'sd-0.08820081040542006, 32'sd-0.10246265499157292, 32'sd-0.21892766124041874, 32'sd-0.16300130696633036, 32'sd-0.18692884257206666, 32'sd-0.11825684860211516, 32'sd-0.028090421973778402, 32'sd0.16466566733247637, 32'sd0.029782693538436204, 32'sd0.09166007093307808, 32'sd0.2128679232503067, 32'sd0.08228918078477945, 32'sd0.09564756634451745, 32'sd-0.02569944075500629, 32'sd-0.07098019150627659, 32'sd-0.10201129056837006, 32'sd-0.1271518935058912, 32'sd-0.05682889703836682, 32'sd-0.03976657752213501, 32'sd-0.12281932570050032, 32'sd-0.0025929484119289288, 32'sd0.011429729476399655, 32'sd-0.08856105545584697, 32'sd-0.03210139734901925, 32'sd0.05238085480084795, 32'sd0.01107667487268884, 32'sd0.06743045061361053, 32'sd-0.1151743398173729, 32'sd-0.038469774481866406, 32'sd-0.04573582704617217, 32'sd-0.14647864871901287, 32'sd-0.11269602564197116, 32'sd-0.29154429015900696, 32'sd-0.365485493978742, 32'sd-0.20924901071993865, 32'sd-0.05131750076859505, 32'sd0.02411794636500116, 32'sd0.16279952129549913, 32'sd0.115059596902617, 32'sd0.13938208564790383, 32'sd0.09284019692408713, 32'sd-0.09036939647817083, 32'sd-0.07852887588383126, 32'sd-0.14912199531053463, 32'sd0.005443389922765204, 32'sd0.03902351972558687, 32'sd0.05970035087176051, 32'sd-0.06655508738211106, 32'sd-0.08851559828296382, 32'sd-0.023705444239269072, 32'sd-0.03652385780190987, 32'sd-0.038481590665641, 32'sd0.1259795575852663, 32'sd0.09406385840429644, 32'sd-0.10178994762110878, 32'sd-0.01669633520638237, 32'sd-0.0009492164676600547, 32'sd-0.10080234183751141, 32'sd-0.12270285571959744, 32'sd-0.13504780702412286, 32'sd-0.24867934018842397, 32'sd-0.352306078854389, 32'sd-0.23861513693254155, 32'sd-0.12252071134021875, 32'sd-0.06638354108760923, 32'sd0.15248447976761226, 32'sd0.1699483505218169, 32'sd-0.02440306624605403, 32'sd-0.015522982754338683, 32'sd-0.06540305399423943, 32'sd-0.11298574066303915, 32'sd-0.0372090201572634, 32'sd-0.07684223805833319, 32'sd-0.06850271917573723, 32'sd0.024560253026220436, 32'sd-0.18210954252567538, 32'sd-0.08975636935804418, 32'sd-0.03486294526996259, 32'sd-0.08326477636095629, 32'sd-0.0608792958004271, 32'sd-0.019740368018165852, 32'sd0.015018111969797306, 32'sd-0.0110262225350306, 32'sd0.03894575127395036, 32'sd-0.043678932463333944, 32'sd-0.10150796464378092, 32'sd-0.21459699682939146, 32'sd-0.23996998271389383, 32'sd-0.1073447541671114, 32'sd-0.18472103734938744, 32'sd-0.05455230117021041, 32'sd-0.05623892710936174, 32'sd0.029920342668527444, 32'sd0.11318108485945619, 32'sd0.23288829595264404, 32'sd0.019444476408253683, 32'sd0.006643649759516924, 32'sd-0.021047119275721553, 32'sd-0.035917060182063865, 32'sd-0.16985336462430542, 32'sd-0.08689177510831655, 32'sd-0.034351717678045963, 32'sd0.09503146851659011, 32'sd-0.12674366604526596, 32'sd0.06287763785305885, 32'sd0.15293563455048625, 32'sd0.009327361507909297, 32'sd-0.02553324008845156, 32'sd0.018815684215588668, 32'sd0.0886885206442852, 32'sd0.007140092128482244, 32'sd0.12971073231688005, 32'sd-0.0296122517988915, 32'sd-0.055313165373754795, 32'sd-0.10731801546255382, 32'sd-0.06547649730491581, 32'sd0.053414559509530384, 32'sd-0.06399965250554737, 32'sd-0.0358721382997837, 32'sd-0.0668696107287531, 32'sd-0.030264828012012635, 32'sd0.029718753386901744, 32'sd-0.007657320392481173, 32'sd0.04361966248641368, 32'sd0.049033352315881774, 32'sd0.054751587902495805, 32'sd0.026984773399583637, 32'sd0.013776142821744448, 32'sd-0.01473460435406983, 32'sd-0.021437393522373345, 32'sd-0.06460228340202323, 32'sd-0.0883116226808909, 32'sd-0.06058250950237958, 32'sd0.0537565064388389, 32'sd-0.08841405350248482, 32'sd-0.025037657837801482, 32'sd0.019617503758337335, 32'sd-0.010221610586106385, 32'sd-0.01007914782646839, 32'sd0.08897881174047417, 32'sd0.03597275252370799, 32'sd0.04268478411576054, 32'sd-0.10298265940701384, 32'sd0.018006766862707572, 32'sd0.09147963015755266, 32'sd0.0960152043537889, 32'sd-0.012202579381428064, 32'sd-0.08706057170829602, 32'sd-0.004469418414483634, 32'sd0.0498899749005901, 32'sd0.06889813737665544, 32'sd0.022379176343277615, 32'sd0.10660274968867413, 32'sd-0.020221239390575352, 32'sd0.19475014019664294, 32'sd0.12353767713849956, 32'sd0.012736624852023417, 32'sd-0.016316757522973305, 32'sd0.08891339974902966, 32'sd-0.040278934947016974, 32'sd-0.017504611420027173, 32'sd0.05516787293428029, 32'sd-0.03636899116624806, 32'sd3.4108290461104333e-121, 32'sd-0.025857325997446515, 32'sd0.014692037240577818, 32'sd-0.01695111075106547, 32'sd-0.04216712826115556, 32'sd-0.05022036034696663, 32'sd0.03780796037068375, 32'sd0.13030264943103192, 32'sd0.04132208894578416, 32'sd0.154587024922841, 32'sd0.0025111057545662858, 32'sd0.05354360542141768, 32'sd-0.1500802016365176, 32'sd-0.12287382475276268, 32'sd-0.02013347806662678, 32'sd0.18965888105186765, 32'sd0.11017662533759158, 32'sd0.03692491265815072, 32'sd0.12263607547533303, 32'sd0.06352309464127844, 32'sd0.07626690103862467, 32'sd0.0432599804816619, 32'sd0.026838816018680017, 32'sd0.08449878875890028, 32'sd-0.059598626644643694, 32'sd0.08151039607588341, 32'sd-0.00563703850186334, 32'sd-0.0498912018546461, 32'sd0.00572246437175367, 32'sd0.04238393038714195, 32'sd0.0032509706037484737, 32'sd0.001963961955527861, 32'sd0.008236785279373432, 32'sd0.05023276745564428, 32'sd0.016034906481400848, 32'sd0.08258287612727831, 32'sd0.05269591087870212, 32'sd0.11795890815686073, 32'sd0.025377820949181493, 32'sd-0.05080397648799004, 32'sd-0.10455696439748384, 32'sd-0.06842944516315991, 32'sd0.09800890584294217, 32'sd0.0870429653168808, 32'sd0.06098433113227523, 32'sd0.08933793992769093, 32'sd-0.0022950037787412506, 32'sd0.11755911248909048, 32'sd0.24359438131491462, 32'sd0.05683573183368099, 32'sd-0.0740856206251413, 32'sd-0.047794513085752624, 32'sd0.1132625806105232, 32'sd-0.020952038820655147, 32'sd0.12629835329776226, 32'sd0.10565349657384741, 32'sd-0.047339833208869905, 32'sd0.03783892870043726, 32'sd0.018418672086451655, 32'sd0.07899064157717421, 32'sd0.14652478981990763, 32'sd0.03937928334828717, 32'sd0.0351055377519604, 32'sd0.14818726661421222, 32'sd0.1490240544648161, 32'sd0.05870067846302836, 32'sd0.004518083286281845, 32'sd-0.04050006650652371, 32'sd-0.10141573907986529, 32'sd-0.08430673723110442, 32'sd-0.019790015546122752, 32'sd-0.03807027135467371, 32'sd0.0223410755041067, 32'sd-0.0008509043279464284, 32'sd0.06889807230621275, 32'sd0.10455375313818804, 32'sd0.12000959108916535, 32'sd0.0192904572960417, 32'sd-0.05893015068957091, 32'sd-0.004114949934851619, 32'sd0.10582798359243996, 32'sd0.06147722889593652, 32'sd0.0364975837238546, 32'sd0.06742120727144754, 32'sd2.3344931348560682e-119, 32'sd-0.01668280194154934, 32'sd-0.02766057594963831, 32'sd-0.02011783116052197, 32'sd0.014428499710411304, 32'sd-0.029479426569699582, 32'sd-0.009746468374346355, 32'sd0.09071594672968943, 32'sd0.04310415906654139, 32'sd-0.0977846528510442, 32'sd-0.07652370960148153, 32'sd-0.2203200300173867, 32'sd-0.12200493711720964, 32'sd-0.01155430629549641, 32'sd-0.18086699419276137, 32'sd-0.002822229443763186, 32'sd0.03635126006612924, 32'sd0.02204498098323377, 32'sd-0.0343302568972634, 32'sd0.1437336759463961, 32'sd0.03360718502518908, 32'sd-0.10226691569156252, 32'sd-0.044558291194614644, 32'sd-0.15279253532574202, 32'sd0.038381367950220194, 32'sd0.06763094054627292, 32'sd0.08448806694881138, 32'sd-0.014387740012328573, 32'sd0.0928929091801529, 32'sd-0.03440478973178981, 32'sd-0.0038105338759837964, 32'sd-0.0008656968142661305, 32'sd0.07732205718480747, 32'sd-0.05486327954280781, 32'sd0.0553951397539606, 32'sd-0.003845963220225555, 32'sd0.02957471215193618, 32'sd-0.00505073230756599, 32'sd-0.09545957567433651, 32'sd-0.17710766275197803, 32'sd-0.04626979675579047, 32'sd-0.020502365509922765, 32'sd-0.0011455359811261409, 32'sd-0.11106902694206512, 32'sd-0.06887411960483632, 32'sd0.003158490360786521, 32'sd-0.04762456221103726, 32'sd-0.008403520053832386, 32'sd-0.01353800078392695, 32'sd-0.05172526105832822, 32'sd-0.13513881105373285, 32'sd-0.09073777059284222, 32'sd0.052341078837747385, 32'sd-0.011124918030674962, 32'sd0.015160340815896664, 32'sd0.011273151016481582, 32'sd0.04714906065865652, 32'sd0.04929947778627882, 32'sd-0.09758517041717493, 32'sd-0.043929179617244525, 32'sd0.08331691767365582, 32'sd0.02750133075468667, 32'sd-0.05366170106832905, 32'sd0.06369795581461, 32'sd-0.05185526596454613, 32'sd-0.11893410526414955, 32'sd-0.05730635411980482, 32'sd0.03850206358872466, 32'sd-0.1328241090399891, 32'sd-0.016653278458198237, 32'sd0.013922466011048658, 32'sd0.004203929835331389, 32'sd-0.0983813189146898, 32'sd0.09548068760560001, 32'sd0.01692874389917468, 32'sd-0.0983772909382891, 32'sd-0.17775991337432112, 32'sd0.05330419670201452, 32'sd-0.1249990729263383, 32'sd-0.11668662758512512, 32'sd-0.08201602593404408, 32'sd-0.009609933914090964, 32'sd0.002281204078094215, 32'sd-0.057124353294376644, 32'sd4.6701882583820285e-115, 32'sd0.014154279075442174, 32'sd-0.0589910357117718, 32'sd-0.0429806673281354, 32'sd0.02956468888438727, 32'sd0.024377020019898, 32'sd0.010836686191213606, 32'sd-0.015417256202879273, 32'sd0.05850441202567661, 32'sd-0.05151484414797487, 32'sd0.046254128916775626, 32'sd-0.06558633446871333, 32'sd-0.07919748014483416, 32'sd-0.08352826090043204, 32'sd0.001861835136650946, 32'sd0.058696153311430105, 32'sd0.1123710300315338, 32'sd0.14302223694349583, 32'sd-0.14327470935434378, 32'sd-0.1166588432998086, 32'sd-0.010688791108129638, 32'sd-0.0786638423037147, 32'sd-0.08963436692678615, 32'sd0.002701000672872956, 32'sd-0.10631241754133504, 32'sd0.017367573428121248, 32'sd-0.0579233805730459, 32'sd3.423503292323921e-121, 32'sd3.858292251712735e-124, 32'sd-1.6976156258226562e-125, 32'sd-0.05507578018794877, 32'sd0.032944856166854955, 32'sd-0.067160471828741, 32'sd-0.09429720635536455, 32'sd0.009443538604994268, 32'sd-0.13360742448554244, 32'sd0.028070134257686064, 32'sd0.013265900693058552, 32'sd0.04719116668517357, 32'sd0.03338723404693825, 32'sd0.11501936382271868, 32'sd0.08535398878903802, 32'sd-0.12506340549837913, 32'sd-0.02566534890174773, 32'sd0.09524154243867414, 32'sd-0.07929371875807097, 32'sd-0.07212629346212772, 32'sd-0.19320625327299987, 32'sd-0.039472305414276376, 32'sd0.017593699455482725, 32'sd0.02543801995622524, 32'sd0.014310166080970637, 32'sd-0.08291529669736972, 32'sd0.013307771402379577, 32'sd-0.044646055196354215, 32'sd-2.0924676455683773e-117, 32'sd-3.1717021288913943e-119, 32'sd1.808602561445324e-120, 32'sd-0.03406921513939342, 32'sd0.05832763483296514, 32'sd-0.02824449246219885, 32'sd0.046728427786856354, 32'sd0.08432349850984061, 32'sd0.02634925844715965, 32'sd0.03935691118635717, 32'sd0.03193954387948851, 32'sd0.05743857893276685, 32'sd0.04635206439475307, 32'sd0.1325793818661197, 32'sd0.03505397080849173, 32'sd0.09352073788622631, 32'sd0.06330993755188674, 32'sd-0.11009780929483091, 32'sd-0.0768101996642267, 32'sd-0.12409042528777904, 32'sd-0.017793660815122056, 32'sd0.034394906714843416, 32'sd0.019351581373222154, 32'sd0.023767525345525058, 32'sd-0.0408546028982228, 32'sd-0.03719738370588163, 32'sd0.0711736132273202, 32'sd0.03044794340007506, 32'sd2.170581012745817e-120, 32'sd-7.39757382070095e-127, 32'sd1.8521604824485967e-126, 32'sd1.0865467251411313e-114, 32'sd-0.019501217603278543, 32'sd0.007977209838842243, 32'sd-0.06001711105723928, 32'sd-0.006678661692795629, 32'sd0.018518824855252608, 32'sd-0.05987592990270299, 32'sd0.0009203764569799906, 32'sd0.06501399284898497, 32'sd-0.03490987367833055, 32'sd-0.13891488934323543, 32'sd-0.020440141227004726, 32'sd0.03714121794337245, 32'sd-0.1488974504662024, 32'sd-0.10537561663968963, 32'sd-0.16683063461718722, 32'sd-0.04242771962959809, 32'sd0.02919395888517019, 32'sd-0.03131950466416751, 32'sd-0.0013747650811349972, 32'sd-0.0010740335702805076, 32'sd0.010355699857648617, 32'sd0.04712215051084584, 32'sd0.02058180204986883, 32'sd8.522460846307603e-121, 32'sd-3.3277540869677338e-121, 32'sd-7.475205357791852e-115, 32'sd2.2326472218903784e-118, 32'sd-4.4891151568624955e-126, 32'sd-1.0957864286208996e-120, 32'sd-0.029164914168355746, 32'sd0.08975937118612166, 32'sd-0.05642586496912379, 32'sd-0.030796248694643185, 32'sd0.07046706062966754, 32'sd-0.032836286069188335, 32'sd-0.07122698578042691, 32'sd-0.04589803667002691, 32'sd0.02744376556174146, 32'sd-0.06069498398554357, 32'sd-0.09995538798952609, 32'sd-0.07496907006031532, 32'sd-0.02286605339444179, 32'sd0.053211719299775556, 32'sd-0.04204668088428484, 32'sd-0.02580796503806224, 32'sd-0.06682897586778894, 32'sd0.005736255304126562, 32'sd0.020610902052744455, 32'sd0.027279781352065567, 32'sd2.4919825942312996e-126, 32'sd1.1392525594244812e-119, 32'sd8.880381634438733e-119, 32'sd-8.393973130885976e-121},
        '{32'sd-1.184017291828846e-117, 32'sd2.577698742866111e-115, 32'sd7.69133463476756e-127, 32'sd-1.9961779045957894e-121, 32'sd-8.789580347647744e-127, 32'sd1.168073012083287e-118, 32'sd1.9601153990070945e-127, 32'sd3.424524426123196e-118, 32'sd-3.2079500315094644e-118, 32'sd3.3941283057569395e-120, 32'sd-3.4898085435206704e-125, 32'sd-6.09826803682351e-121, 32'sd0.07202597281289617, 32'sd-0.0006511324968407956, 32'sd0.1286890222805566, 32'sd-0.004760553133347568, 32'sd2.994398219826887e-122, 32'sd2.971010348662665e-116, 32'sd1.884108581155819e-123, 32'sd-2.5908839532219805e-126, 32'sd7.36911442264558e-122, 32'sd-2.4162851146933874e-126, 32'sd6.605338961281076e-116, 32'sd-3.6140126138231234e-126, 32'sd-1.5859815081838258e-115, 32'sd1.5806801047286227e-125, 32'sd-3.974387843864905e-123, 32'sd-4.3285163484949106e-125, 32'sd-3.71418653111858e-125, 32'sd-5.098627258569533e-118, 32'sd1.0740257600776952e-127, 32'sd-1.5770507171037578e-125, 32'sd-0.02750966720359166, 32'sd0.09234687638366566, 32'sd0.03609838785819513, 32'sd-0.030183969111329405, 32'sd0.03534347440675384, 32'sd0.06761074387756649, 32'sd0.01942078974104011, 32'sd-0.028653720880619914, 32'sd0.009435118490879588, 32'sd-0.004014270881792701, 32'sd0.04848648962984463, 32'sd0.07055419133257966, 32'sd0.02389323391945106, 32'sd0.026624372933859317, 32'sd-0.012720176408540902, 32'sd0.03578919999072194, 32'sd0.021150757829635148, 32'sd-0.05460438697083906, 32'sd0.0150350561894272, 32'sd-0.0003959452221167596, 32'sd3.5586493315568264e-117, 32'sd-2.2578331593216943e-121, 32'sd-2.581937454228662e-119, 32'sd-3.345416807473062e-122, 32'sd-8.886374525857307e-127, 32'sd-1.3951335714249584e-117, 32'sd0.06971367512695173, 32'sd0.018001473526008095, 32'sd-0.06452397472158174, 32'sd0.042097428924987634, 32'sd0.05883231392824625, 32'sd-0.07121397112130441, 32'sd-0.027093324757502417, 32'sd-0.03328177125028859, 32'sd0.1394496356915691, 32'sd-0.04786249204566954, 32'sd0.10829577600307586, 32'sd0.14931213728407552, 32'sd0.12782133365160042, 32'sd0.08497350185665303, 32'sd0.17379803834916507, 32'sd0.10586844296842522, 32'sd0.03774702772291062, 32'sd-0.024390905414622053, 32'sd0.01672983483263711, 32'sd-0.0035728886675745444, 32'sd0.012942561554573654, 32'sd0.03897554260626025, 32'sd0.021585902254904973, 32'sd0.02555826523918573, 32'sd8.888997129434636e-127, 32'sd1.7718091269644236e-116, 32'sd-3.888321198926996e-123, 32'sd3.50612162781735e-114, 32'sd0.08257960927924729, 32'sd0.011393241341344793, 32'sd0.048114610356522085, 32'sd-0.13498249298082807, 32'sd-0.00789062556396481, 32'sd-0.08651017881850219, 32'sd0.022226091293663718, 32'sd0.005683616868845687, 32'sd0.01816291533279012, 32'sd-0.030539899636996003, 32'sd0.03199974713496503, 32'sd0.06903523519437159, 32'sd-0.04117766565621112, 32'sd0.18103837357878746, 32'sd0.11823228792720349, 32'sd0.11113156081676537, 32'sd-0.0528071310758725, 32'sd0.04834472849712641, 32'sd0.013718005978175142, 32'sd-0.005892859353774727, 32'sd-0.015014950233536406, 32'sd0.05852436559735753, 32'sd-0.014141103939029473, 32'sd-0.020409688546766253, 32'sd0.027753020318111877, 32'sd3.5127726283479693e-122, 32'sd3.7507095454574116e-124, 32'sd0.05281868687486315, 32'sd-0.05223322506646338, 32'sd0.04841329158936365, 32'sd-0.040156024453470655, 32'sd-0.05017779003119199, 32'sd-0.061727035388072365, 32'sd-0.04628903002339079, 32'sd-0.14084225405318723, 32'sd-0.17586067330030097, 32'sd-0.09158407763378512, 32'sd0.0697342579877645, 32'sd0.08985398269924567, 32'sd-0.0028874232241990175, 32'sd0.16528708894985, 32'sd0.09930563355011024, 32'sd0.17344998192575464, 32'sd0.012595003367611818, 32'sd0.05781175851584399, 32'sd0.09538618868940786, 32'sd-0.040898299545732125, 32'sd-0.11403899064592422, 32'sd0.00151409447621855, 32'sd-0.06036023186186301, 32'sd-0.15371149350875807, 32'sd-0.0727002084349101, 32'sd-0.00871749540145453, 32'sd0.0008325444535981029, 32'sd-2.605523586098045e-126, 32'sd0.07591814672068319, 32'sd0.01581916179868874, 32'sd0.024817304708083195, 32'sd0.0378247818470676, 32'sd-0.050720777033076654, 32'sd-0.06181620080662472, 32'sd-0.10266674614903414, 32'sd-0.06346817655500037, 32'sd-0.11073729140834347, 32'sd-0.12639378755833558, 32'sd-0.08186894026121773, 32'sd0.02101124960552676, 32'sd0.025538151001607893, 32'sd0.12126019067388624, 32'sd0.10886168337566564, 32'sd0.15686214554602393, 32'sd-0.01810917066523328, 32'sd0.12708632144117876, 32'sd0.1092989814839137, 32'sd0.0027939870352492813, 32'sd-0.04526718481698299, 32'sd0.11183340883952148, 32'sd0.009133623152255636, 32'sd-0.10286770035883759, 32'sd0.04148769114237525, 32'sd-0.07949803611872763, 32'sd-0.01004853138065785, 32'sd5.435578875853387e-118, 32'sd-0.0035377900789180863, 32'sd0.04700827739173858, 32'sd-0.004422773479359136, 32'sd0.01522441851456784, 32'sd-0.07926655708762465, 32'sd-0.08442369743428575, 32'sd0.025841636233284684, 32'sd-0.07372015951947095, 32'sd-0.06769793052502303, 32'sd-0.04440191653052002, 32'sd-0.14378017605030868, 32'sd-0.0819674595920474, 32'sd-0.08673083095137075, 32'sd-0.08785788513281272, 32'sd0.16755334577215214, 32'sd0.05957732012506413, 32'sd-0.04798969719706257, 32'sd0.1502704971796528, 32'sd0.02928842924555354, 32'sd0.03570594529278539, 32'sd0.041259055799866544, 32'sd-0.07120579170062413, 32'sd-0.01139125364899405, 32'sd0.006153305321075589, 32'sd0.06725311362061667, 32'sd-0.12527239583750463, 32'sd0.04258144863546623, 32'sd0.011391436350483985, 32'sd-0.016234478605569303, 32'sd0.04448342648427198, 32'sd0.08728674594136625, 32'sd-0.02540586574631028, 32'sd-0.040432223662381556, 32'sd-0.07869227978819715, 32'sd-0.029772656684161458, 32'sd-0.10633703295155253, 32'sd0.05150048658699286, 32'sd-0.12983754676743406, 32'sd-0.1949817634801045, 32'sd-0.2713982277807973, 32'sd-0.16421517718532785, 32'sd-0.03917756396003109, 32'sd0.092254024573669, 32'sd0.11730960272883421, 32'sd0.09264398439161851, 32'sd0.10468319465067649, 32'sd0.1880181538669916, 32'sd0.04121558228175455, 32'sd-0.004042742540032863, 32'sd0.06984854841725721, 32'sd-0.06501899619759724, 32'sd-0.13167426386351314, 32'sd0.04202189338658855, 32'sd-0.03959740280559134, 32'sd-0.02837604011014565, 32'sd0.03601713823698482, 32'sd0.12747759271434025, 32'sd-0.008475452442205694, 32'sd-0.02276575337301295, 32'sd-0.06023594949066857, 32'sd0.06440878882888053, 32'sd0.06651344925816183, 32'sd-0.06648871165198962, 32'sd-0.1222702445575647, 32'sd-0.00796267416812989, 32'sd-0.14950335468318196, 32'sd-0.3119323718824189, 32'sd-0.3330193314997902, 32'sd-0.22680077826884915, 32'sd-0.04738970557901986, 32'sd0.02637000401674348, 32'sd0.07748939086198349, 32'sd0.15412274120916328, 32'sd-0.0035221826767384717, 32'sd0.05210098566985833, 32'sd-0.009522846978229462, 32'sd-0.06553548302915856, 32'sd-0.08120998038054653, 32'sd0.02019360065597361, 32'sd-0.07066174898828947, 32'sd-0.008768062600267013, 32'sd-0.022838062731627338, 32'sd0.049613954564747334, 32'sd-0.059488444906852955, 32'sd0.08628267469934023, 32'sd-0.028254682845394032, 32'sd0.10367225512864675, 32'sd0.07100385464465978, 32'sd0.021215106491232386, 32'sd-0.06241062783756557, 32'sd-0.0762253419862993, 32'sd0.060976469533347004, 32'sd0.12325116076888339, 32'sd-0.05649207637888124, 32'sd-0.2205327480233945, 32'sd-0.23237197221134678, 32'sd-0.09346567242584357, 32'sd0.11456134498470523, 32'sd0.1343742206667579, 32'sd0.07245490528191617, 32'sd0.06617184170029959, 32'sd0.2018170613743867, 32'sd0.07096015355121983, 32'sd-0.028944294172790003, 32'sd-0.10123730920239216, 32'sd-0.06337953799957041, 32'sd-0.02572794497757034, 32'sd-0.055136636385983345, 32'sd-0.05011222686614901, 32'sd-0.07268756010286519, 32'sd0.0024125962919592328, 32'sd0.03324439384628936, 32'sd0.01795877023364843, 32'sd0.05270538729702871, 32'sd-0.07652534753736095, 32'sd0.015887737312735756, 32'sd-0.06458809877696484, 32'sd0.0787662338488984, 32'sd-0.053705893600035526, 32'sd0.01726395339663185, 32'sd0.06857384538848542, 32'sd-0.013067711611963743, 32'sd-0.014160612644756428, 32'sd-0.10263652464190563, 32'sd-0.055830318428567796, 32'sd0.020285435744270112, 32'sd0.15681481774650824, 32'sd0.13934011853050632, 32'sd0.1729037905498279, 32'sd0.010279120613455938, 32'sd-0.06382269121289141, 32'sd-0.05945823526974745, 32'sd0.0060956581339288085, 32'sd-0.16345775957011882, 32'sd0.049456336546893805, 32'sd-0.07985575652815559, 32'sd0.009042939834246748, 32'sd-0.021501771136119386, 32'sd0.03181878730889948, 32'sd0.007517995956793906, 32'sd0.0818131205875013, 32'sd0.07789367117988195, 32'sd0.11962275864346228, 32'sd-0.055616371872374115, 32'sd0.07551872156562728, 32'sd0.08259502751552752, 32'sd0.0907262651894331, 32'sd0.10269502994040813, 32'sd0.14039786872374613, 32'sd0.028027563751078188, 32'sd-0.12366729198798557, 32'sd-0.1336210797912801, 32'sd-0.09184717450488086, 32'sd0.11006757959686059, 32'sd0.07288178008824149, 32'sd0.11617980886529503, 32'sd0.12771000591136833, 32'sd-0.03600719310372792, 32'sd0.05541790838653757, 32'sd0.06308312926222646, 32'sd-0.04979437513244874, 32'sd-0.07233433582719445, 32'sd0.012721745875990304, 32'sd-0.21047069500832563, 32'sd0.012270451428248851, 32'sd-0.03632013507019358, 32'sd0.019306410729678012, 32'sd0.019660890709574195, 32'sd0.015906112340670474, 32'sd0.03836460941450104, 32'sd0.05792935963970606, 32'sd0.04959600553005579, 32'sd0.09282276460768417, 32'sd0.04069879691088121, 32'sd0.09276084019641012, 32'sd0.03594135905317336, 32'sd0.19042089154176206, 32'sd-0.00255139942791836, 32'sd-0.0502965582525509, 32'sd-0.03702140725747572, 32'sd-0.026425766821468813, 32'sd0.06362205030214736, 32'sd0.04484014062743161, 32'sd0.17341898293140698, 32'sd0.009533545690116517, 32'sd0.02103323246249606, 32'sd0.04203987995540217, 32'sd0.004185125317965329, 32'sd0.020271084323868628, 32'sd-0.12742990450802558, 32'sd0.0043456807923335835, 32'sd-0.09538144677314234, 32'sd-0.03458552597734807, 32'sd0.024796305940862524, 32'sd0.007959373955085652, 32'sd0.049941545437162754, 32'sd-0.07627836918101821, 32'sd-0.030818637047734684, 32'sd0.06319355819473423, 32'sd0.08923216321217559, 32'sd-0.0011141427746955126, 32'sd0.087006588598552, 32'sd-0.012848301385221661, 32'sd-0.06606355450227444, 32'sd0.16396597042518912, 32'sd0.03360817873933285, 32'sd-0.035899453014421795, 32'sd-0.12975017443892348, 32'sd-0.13017842481884695, 32'sd0.05492677685416373, 32'sd0.0022873811471021267, 32'sd0.01637077981728306, 32'sd0.0891444236256848, 32'sd0.10058950187788458, 32'sd-0.10141243028940652, 32'sd-0.03566872465885779, 32'sd-0.032533484806887954, 32'sd-0.15109609144550548, 32'sd-0.14055052138581228, 32'sd-0.015284042179764116, 32'sd-0.051521393337858164, 32'sd-0.05484345053283325, 32'sd-0.0008010787423341695, 32'sd0.0664564081170666, 32'sd0.002953168833408156, 32'sd-0.03273936628779219, 32'sd0.019075272548905415, 32'sd0.06771795490096477, 32'sd0.1436595562890745, 32'sd0.009377028340918164, 32'sd-0.00033114709758163326, 32'sd0.04559982660982097, 32'sd0.03711964491554891, 32'sd-0.06912081496153658, 32'sd-0.11626106096966986, 32'sd-0.045261697142247585, 32'sd-0.047216439347311775, 32'sd0.20288521285305766, 32'sd0.08676318225918628, 32'sd0.23103322433195048, 32'sd-0.03332105223111897, 32'sd0.014198848798623898, 32'sd-0.0056770875411144015, 32'sd-0.13789721699049753, 32'sd-0.08315857257452264, 32'sd-0.1126009077024517, 32'sd-0.18084486326751925, 32'sd0.01745890844069477, 32'sd0.06908323191568799, 32'sd0.0714913904540535, 32'sd0.07258288272231984, 32'sd-0.0415106286199496, 32'sd0.06389669147760119, 32'sd-0.025203085196603008, 32'sd0.0646261442894172, 32'sd0.04642653510067268, 32'sd-0.0285008285549071, 32'sd0.05514660515847872, 32'sd-0.022617030619135243, 32'sd-0.046659084691555296, 32'sd-0.1699006715326982, 32'sd-0.22799481805509242, 32'sd0.06935824735527364, 32'sd0.02082036231096631, 32'sd0.0026014566802379777, 32'sd0.1331377249845182, 32'sd0.10703539703309603, 32'sd0.06409786580839724, 32'sd-0.10244029809080456, 32'sd-0.0961882241621397, 32'sd0.01935846083620079, 32'sd-0.029847940762195026, 32'sd-0.06485824082248659, 32'sd-0.17961565233661422, 32'sd-0.12682702380852257, 32'sd-0.056812653776590734, 32'sd-0.07020599891611827, 32'sd-0.05589932103965555, 32'sd0.05682068400904251, 32'sd0.037095874612556846, 32'sd0.033582235677267425, 32'sd0.05624896648264327, 32'sd0.0010394836965913572, 32'sd-0.030145020698053013, 32'sd-0.11181831261262504, 32'sd0.03323751793473522, 32'sd-0.0815371799124784, 32'sd-0.15097392285226827, 32'sd-0.19608961164950914, 32'sd-0.14762788494364038, 32'sd0.009738097592230708, 32'sd-0.11627441798985012, 32'sd0.07948780430372027, 32'sd-0.01597213902691132, 32'sd-0.0034986259149566196, 32'sd-0.11661790507446818, 32'sd-0.16701673165021927, 32'sd-0.00018821494149329676, 32'sd0.007404955871264765, 32'sd-0.04022157862628408, 32'sd0.027164353081407865, 32'sd-0.13392311617663877, 32'sd-0.06402028528234285, 32'sd0.12202159967921875, 32'sd-0.07777757942556209, 32'sd0.04794260091639657, 32'sd-0.048357923661668266, 32'sd1.9618671230941818e-126, 32'sd0.05122470354428352, 32'sd0.09790026294205285, 32'sd0.021137582679718422, 32'sd0.09398158031346193, 32'sd0.06717815009900241, 32'sd-0.042359895765331626, 32'sd-0.05277090719347564, 32'sd-0.14329465325240126, 32'sd-0.09830985277142998, 32'sd-0.02508013230292063, 32'sd0.031033752138945072, 32'sd0.02354875339705503, 32'sd-0.025808703023942416, 32'sd-0.011528447383797283, 32'sd0.05763405708909856, 32'sd-0.06537104814659306, 32'sd-0.07499962084435924, 32'sd0.007905921126469744, 32'sd0.01576812378731142, 32'sd-0.017467710156613345, 32'sd0.05719416800802737, 32'sd-0.008842109647860237, 32'sd0.044982082983284315, 32'sd0.18393482350933188, 32'sd0.13528364067679544, 32'sd-0.01698179277336296, 32'sd-0.04655313420524079, 32'sd0.026209725751587528, 32'sd-0.029169054205740532, 32'sd0.09220372835410828, 32'sd0.0273885886203507, 32'sd0.007269765673341756, 32'sd-0.028042660211996775, 32'sd-0.027231362277468443, 32'sd0.046714824709861096, 32'sd0.0313361048894585, 32'sd0.027391841349824537, 32'sd0.026745150924263883, 32'sd-0.052106040637579905, 32'sd0.028199856120753694, 32'sd0.08524251838434636, 32'sd0.01843789145601104, 32'sd0.01090928884071783, 32'sd-0.031870108306205465, 32'sd-0.09468927440655237, 32'sd-0.052281778842499425, 32'sd0.018672111581892612, 32'sd0.06561178594153617, 32'sd0.05132091038825742, 32'sd0.005328231485500562, 32'sd0.06502856036545912, 32'sd0.14181418952978506, 32'sd0.17065608721284395, 32'sd0.020381063948007535, 32'sd0.052151687692513625, 32'sd0.09920398662987698, 32'sd-0.0337463142756171, 32'sd-0.003798875430431112, 32'sd-0.05379370618295135, 32'sd0.020834160298597408, 32'sd-0.07540274844843915, 32'sd-0.009336590355816271, 32'sd0.03176645198239871, 32'sd-0.024681150536313128, 32'sd0.15084670961673227, 32'sd0.042131407846066844, 32'sd0.021034552927689826, 32'sd-0.08162147126447777, 32'sd0.11285784084758456, 32'sd-0.006124806090396438, 32'sd-0.03372045530538149, 32'sd0.02570039941339107, 32'sd-0.007951721294059449, 32'sd-0.03130544162767549, 32'sd-0.009749806989716198, 32'sd0.11212610587303917, 32'sd0.06743980945254847, 32'sd-0.008594292257335021, 32'sd0.0608864256534014, 32'sd0.06522589068897298, 32'sd0.07859201984538625, 32'sd-0.06150724614794159, 32'sd0.050855053984815886, 32'sd1.3480511857356447e-126, 32'sd-0.003960695152686589, 32'sd-0.03788334852639284, 32'sd0.11041224943621283, 32'sd0.12043262614245007, 32'sd-0.06479421862436766, 32'sd0.15022167922317683, 32'sd0.1037018615079422, 32'sd0.07110815514547637, 32'sd0.01645290479474264, 32'sd0.07739231492828517, 32'sd0.003885055342662163, 32'sd0.010269038787015433, 32'sd-0.01353517121808871, 32'sd-0.12676728622255304, 32'sd-0.09413959587777022, 32'sd0.14080281191735583, 32'sd0.10680125176690276, 32'sd0.18363010427867646, 32'sd-0.051182927193846345, 32'sd0.02461447174119991, 32'sd-0.022885329482021165, 32'sd0.04171446554263033, 32'sd0.010864215914459298, 32'sd0.13941033401916972, 32'sd0.01765988020196314, 32'sd-0.009756420587708942, 32'sd-0.004963293302459143, 32'sd0.058029298994972084, 32'sd0.056335756456269856, 32'sd0.04653537846659759, 32'sd0.07600587648902714, 32'sd-0.02550698655075962, 32'sd-0.0757409881557405, 32'sd0.07046049387041095, 32'sd0.0957504341220779, 32'sd0.09768772453935684, 32'sd-0.026148694778231694, 32'sd-0.012637164825028701, 32'sd-0.03707736458919216, 32'sd-0.06755773267884517, 32'sd-0.02045815220174299, 32'sd0.012594675959114805, 32'sd-0.013126498560157187, 32'sd-0.061809642103871555, 32'sd-0.021695783805196017, 32'sd-0.020670457220037436, 32'sd-0.02350127112277674, 32'sd-0.029101674134729947, 32'sd-0.05588019132986577, 32'sd-0.006796443156923945, 32'sd-0.0936644201369172, 32'sd0.06428566619006265, 32'sd0.04463777587074719, 32'sd0.06165997349448882, 32'sd0.0005854206537808762, 32'sd0.1231983320037175, 32'sd0.06311295122705564, 32'sd0.0870962211928927, 32'sd-0.04804433866125754, 32'sd0.03224611838267441, 32'sd0.13913873178359276, 32'sd0.06433187169583403, 32'sd0.06130239553137713, 32'sd0.039174548867655035, 32'sd0.019910321176401034, 32'sd-0.07155034995122757, 32'sd0.08183125332801383, 32'sd-0.012214454014276203, 32'sd-0.07851016186390396, 32'sd0.08947375850549885, 32'sd-0.032696993628881656, 32'sd0.037679970019194396, 32'sd0.035256133137158294, 32'sd0.043475493259186225, 32'sd-0.08030718868840432, 32'sd-0.055012865381120664, 32'sd0.062122667070484465, 32'sd-0.02013723749324471, 32'sd-0.03384126423606635, 32'sd-0.09255280846729622, 32'sd-0.010549068941220673, 32'sd-0.0061124111346751745, 32'sd0.004612959918491091, 32'sd-4.652928455476229e-127, 32'sd-0.05477329285133306, 32'sd-0.0161641679342772, 32'sd0.07419911266893832, 32'sd0.08711192213046816, 32'sd0.049582545175296935, 32'sd0.050097045062667496, 32'sd-0.09776307653785664, 32'sd-0.053401349217341326, 32'sd0.060671061801663054, 32'sd0.04301311404275736, 32'sd-0.008544830536821655, 32'sd0.03060455727186871, 32'sd0.1453560569658883, 32'sd0.16484717283636147, 32'sd0.12112524093449574, 32'sd0.06389029347501908, 32'sd0.007973278435755937, 32'sd0.003568070733815119, 32'sd-0.0012778190136136813, 32'sd0.03246039632068915, 32'sd-0.016838035546662796, 32'sd-0.050170572858298845, 32'sd-0.05923855602608089, 32'sd-0.08441936756348765, 32'sd0.025240762188239816, 32'sd0.07743753606168971, 32'sd-9.946605236383831e-124, 32'sd1.0147849492832761e-118, 32'sd3.4112053213398297e-116, 32'sd-0.05692236704208976, 32'sd-0.0006501929611323373, 32'sd0.07816159597396052, 32'sd0.05445714973284295, 32'sd-0.054567374962034065, 32'sd-0.078113903173023, 32'sd-0.08791171129568101, 32'sd-0.08783628317443039, 32'sd-0.0925060186944842, 32'sd0.019149406142781843, 32'sd-0.04300310407887802, 32'sd0.041279060713788805, 32'sd0.16433200068170312, 32'sd0.09485826338802214, 32'sd-0.03532600671894952, 32'sd-0.10218417570119952, 32'sd0.0946705142514664, 32'sd0.10936168402116087, 32'sd0.059524489522294895, 32'sd-0.038023180388557176, 32'sd-0.09677017480162495, 32'sd-0.0728562276860518, 32'sd-0.06408708613033146, 32'sd0.04163408979719745, 32'sd0.07285909537196858, 32'sd-2.8580612233380113e-120, 32'sd-1.4096200940209915e-116, 32'sd-2.0964330550821136e-120, 32'sd-0.011245936383292741, 32'sd0.026504160246429924, 32'sd0.03298329016396879, 32'sd0.010153342510901197, 32'sd-0.02431048072582224, 32'sd-0.10389547973709899, 32'sd0.07937073752886058, 32'sd0.08300309877848451, 32'sd-0.17928151137349568, 32'sd-0.13945994745595688, 32'sd0.013256048063780225, 32'sd-0.07086990017336012, 32'sd-0.05307481495295947, 32'sd-0.11462386654249673, 32'sd-0.11966750736003692, 32'sd0.15305174004675384, 32'sd0.14100085417646058, 32'sd0.04733698044993856, 32'sd-0.1095512551543993, 32'sd-0.05584136378702819, 32'sd-0.02513129522333509, 32'sd-0.07845084049157999, 32'sd-0.064858176921422, 32'sd0.06279476263672823, 32'sd-0.03048254019424967, 32'sd-1.845680918809125e-119, 32'sd-2.925144700350392e-125, 32'sd5.397052487916108e-123, 32'sd1.6890264346675015e-115, 32'sd0.011573064011248153, 32'sd0.018599861513560436, 32'sd-0.052969388580101015, 32'sd0.016437419778045848, 32'sd0.05174053233673788, 32'sd0.012945025597699207, 32'sd-0.08974867640073107, 32'sd0.042119912318977965, 32'sd0.06159139556347788, 32'sd0.05493039969183566, 32'sd-0.00821792522156399, 32'sd-0.03982132081244372, 32'sd-0.0542164164425599, 32'sd0.08469486270700827, 32'sd-0.1189561895360322, 32'sd-0.09251113375544695, 32'sd-0.12303372749628642, 32'sd-0.10943203242237232, 32'sd-0.06873622200773187, 32'sd-0.020569070120439053, 32'sd0.032231488751520605, 32'sd0.04635689018956607, 32'sd0.09972197502926271, 32'sd-1.759299884514858e-117, 32'sd5.470154737327435e-121, 32'sd-3.8961013833355417e-119, 32'sd3.222853041301528e-121, 32'sd1.315270913424157e-116, 32'sd1.343147365934102e-121, 32'sd0.0648763339710035, 32'sd0.02369409513223988, 32'sd0.0624045996186837, 32'sd0.029982826877926565, 32'sd-0.030057640923113776, 32'sd-0.04514157867921821, 32'sd0.0003508058863995215, 32'sd-0.08646436677397917, 32'sd-0.037284221458896816, 32'sd-0.04983295316389626, 32'sd0.005000240537905654, 32'sd0.01201893155857965, 32'sd0.10405021366084935, 32'sd0.09449349908807732, 32'sd0.06795921862893509, 32'sd0.004136848630719862, 32'sd-0.0384503789377217, 32'sd0.05179113589163804, 32'sd-0.061668162582981065, 32'sd-0.01810072132884596, 32'sd5.360004583704505e-118, 32'sd5.6484230320744394e-126, 32'sd7.727402235598269e-125, 32'sd2.142962924471766e-127},
        '{32'sd1.4556435244054126e-125, 32'sd2.618735902223262e-119, 32'sd-2.8361062264850867e-120, 32'sd3.594583209290056e-124, 32'sd1.6937606274842974e-126, 32'sd3.711621273947366e-126, 32'sd1.3864893961382553e-118, 32'sd7.616010330845094e-127, 32'sd9.020348475461748e-123, 32'sd8.731921012668725e-127, 32'sd-1.50986152740288e-119, 32'sd3.503516722227921e-115, 32'sd0.06472934122760746, 32'sd0.07413228579995634, 32'sd-0.04568766677769035, 32'sd0.022641869344348968, 32'sd-5.232971908938411e-123, 32'sd-9.293106354110307e-121, 32'sd-1.2052845176967141e-117, 32'sd5.221417436097839e-125, 32'sd3.291300692161165e-122, 32'sd-2.7977295585239133e-123, 32'sd-1.0088317386375274e-115, 32'sd-1.3616109167578807e-118, 32'sd3.352737207037307e-121, 32'sd-7.273677947894303e-115, 32'sd8.523466310167957e-127, 32'sd3.5827398156182556e-123, 32'sd2.1527934243004145e-127, 32'sd-1.0588978563087515e-121, 32'sd6.296799032389282e-127, 32'sd1.8718139927883018e-122, 32'sd0.02490688251932774, 32'sd0.06014685545671809, 32'sd-0.0330975275585531, 32'sd0.07688270940448819, 32'sd0.07767305599639959, 32'sd0.08097090340656543, 32'sd0.06267882485505824, 32'sd0.09196942241439456, 32'sd0.09592889871493691, 32'sd-0.01769652824122983, 32'sd-0.041911084716140315, 32'sd0.060028245574604545, 32'sd0.07666264817469495, 32'sd-0.025589205265184777, 32'sd0.03473678127617539, 32'sd-0.035648754516938774, 32'sd-0.07655283547663153, 32'sd-0.05816945848977028, 32'sd-0.0431923889639513, 32'sd0.04683393468197938, 32'sd1.149803530765262e-117, 32'sd-1.0998626979162599e-119, 32'sd-1.2118090380854528e-116, 32'sd1.781401123844547e-118, 32'sd-3.069795209342973e-116, 32'sd3.563923165641434e-123, 32'sd0.027724792073684078, 32'sd-0.04477459293998596, 32'sd-0.02201224640135945, 32'sd0.10760786067880303, 32'sd-0.007876849587808533, 32'sd-0.0485650813171738, 32'sd0.061568261455316485, 32'sd0.08441926087225102, 32'sd-0.03007563526240952, 32'sd0.11256292489983112, 32'sd0.044925382204474534, 32'sd0.13515294024605226, 32'sd0.09597948962419486, 32'sd0.0452123265728047, 32'sd0.027513649825271724, 32'sd-0.07698820098659843, 32'sd-0.12440541845376908, 32'sd0.04379615599937986, 32'sd0.07697000105066978, 32'sd-0.05329820524631736, 32'sd-0.0005315047829796381, 32'sd0.02916190784030741, 32'sd0.06441766260404713, 32'sd0.02564399222557369, 32'sd-3.204098286923655e-116, 32'sd1.7580926593718192e-119, 32'sd1.6095382637377528e-127, 32'sd6.27036731224231e-123, 32'sd-0.02079015917575372, 32'sd0.0028335224216553684, 32'sd-0.04059515117668935, 32'sd0.0313299886360299, 32'sd0.08540157017913953, 32'sd-0.022999919994403296, 32'sd0.0891090204848307, 32'sd0.18603223849963782, 32'sd0.09724466488647993, 32'sd-0.08515151930491895, 32'sd-0.023934820538991007, 32'sd0.043363893906623305, 32'sd0.09451402025796168, 32'sd-0.005194230901313202, 32'sd-0.06843268623842101, 32'sd-0.0360253457891619, 32'sd-0.0030261239008488464, 32'sd0.0012469078536987163, 32'sd-0.0867789854801941, 32'sd-0.06792411849013369, 32'sd0.009585936780479181, 32'sd-0.07748871447714267, 32'sd0.016577401302890215, 32'sd0.05919278439950081, 32'sd-0.02369618004024634, 32'sd-2.65174683827102e-122, 32'sd2.8376218793699764e-116, 32'sd-0.015252206872901432, 32'sd0.007566658135557386, 32'sd0.02191126497806276, 32'sd-0.10178692658862411, 32'sd0.025284742842791554, 32'sd0.11162585263363506, 32'sd0.07755835146893832, 32'sd0.02355223476618438, 32'sd-0.08617673407212138, 32'sd-0.02037198585480117, 32'sd-0.03142614026924548, 32'sd0.10019188884473385, 32'sd0.0142730401502847, 32'sd0.06777393708818454, 32'sd-0.0059673004909366134, 32'sd-0.13771619680283778, 32'sd-0.08315156981043473, 32'sd-0.15264524851386493, 32'sd-0.15811551094945459, 32'sd-0.11612952925382426, 32'sd-0.10192172823147243, 32'sd-0.1337633749927867, 32'sd-0.12399319419117552, 32'sd0.021609520400479202, 32'sd-0.0013173352640868997, 32'sd-0.08968819141271386, 32'sd-0.041949649217853206, 32'sd2.947876926521105e-128, 32'sd0.036165697212675645, 32'sd-0.030530044145650075, 32'sd-0.05709909419714112, 32'sd0.0003902668215072101, 32'sd0.008103861375938928, 32'sd0.08801494015670396, 32'sd-0.11137180949975567, 32'sd-0.097030464595615, 32'sd-0.014743028179830656, 32'sd-0.0025702564207046217, 32'sd0.03937603375882871, 32'sd0.16228821435188642, 32'sd0.13975375814583366, 32'sd-0.03408608024426571, 32'sd0.009245544509039192, 32'sd-0.014213342772391044, 32'sd-0.0733436294132197, 32'sd-0.048239109983612576, 32'sd-0.12188737224540469, 32'sd-0.02804407478721784, 32'sd-0.09897165275001928, 32'sd-0.11435951055911879, 32'sd0.0238183233005877, 32'sd0.03921050860140394, 32'sd0.00810105819936833, 32'sd-0.051175438243784246, 32'sd-0.014430152814535713, 32'sd-1.0659143544361087e-124, 32'sd-0.046257919818630255, 32'sd0.003888833575149309, 32'sd0.024944167243492885, 32'sd-0.023663728510534377, 32'sd-0.04642598973245567, 32'sd-0.09045547513419509, 32'sd-0.07723972726422805, 32'sd-0.04927460672341383, 32'sd0.0842385688729025, 32'sd-0.015278495231017776, 32'sd-0.02483672133021306, 32'sd0.1341762937649597, 32'sd0.07105468360883964, 32'sd0.07705954767696002, 32'sd-0.02624065244859618, 32'sd-0.039104025842485936, 32'sd0.004975044333834802, 32'sd0.007516348905619601, 32'sd-0.08300842513010544, 32'sd-0.08496045994966865, 32'sd0.04656858205085492, 32'sd-0.09640448612100776, 32'sd-0.02484638171247415, 32'sd-0.1282340736332448, 32'sd-0.11760341612178674, 32'sd0.09953595929437548, 32'sd-0.040145633077620084, 32'sd-0.017155174699923597, 32'sd0.09167140283747666, 32'sd-0.06573074549204902, 32'sd0.06253297241544789, 32'sd0.05485554211391231, 32'sd-0.08244147848069121, 32'sd-0.11018277140844059, 32'sd-0.09981285813662301, 32'sd0.11558252756560419, 32'sd0.09248503660254905, 32'sd-0.02751300475331839, 32'sd-0.02692694242431848, 32'sd0.0021221188757787586, 32'sd0.009895180783908782, 32'sd-0.02758528635789206, 32'sd-0.03727889203475059, 32'sd-0.02952891809462605, 32'sd-0.007952010272088472, 32'sd0.12147227015321312, 32'sd0.00870721514971122, 32'sd-0.06474005290658208, 32'sd-0.018167988820603182, 32'sd-0.06532392863903085, 32'sd-0.09269884682624467, 32'sd-0.06634451090796437, 32'sd-0.05595985876213811, 32'sd-0.04310363660227444, 32'sd0.025602114673550135, 32'sd-0.045186740886137285, 32'sd-0.03255554573390036, 32'sd0.012674276461122928, 32'sd-0.008260365359687662, 32'sd-0.005382894001991813, 32'sd0.03102013987041978, 32'sd-0.08565005188973011, 32'sd0.018164335546590592, 32'sd0.1814751237613116, 32'sd-0.015577412626655235, 32'sd-0.03171476803271773, 32'sd-0.18839686836381012, 32'sd-0.11913247458950703, 32'sd-0.15265767571814354, 32'sd0.024618123548894092, 32'sd0.03301458844367794, 32'sd-0.03965400645919476, 32'sd0.055731395854517474, 32'sd-0.0039591225600854795, 32'sd-0.0871690238445533, 32'sd-0.08652244274528767, 32'sd-0.05680147694452637, 32'sd-0.04596155808874128, 32'sd-0.03368039377818446, 32'sd-0.03517895429088795, 32'sd-0.055064890580988485, 32'sd-0.1061619242591221, 32'sd-0.052718264299564874, 32'sd0.09377402765040597, 32'sd0.016534204606121396, 32'sd-0.2107843510616385, 32'sd-0.016143925784243552, 32'sd-0.005930616583614652, 32'sd0.0955438111961438, 32'sd0.12521772839760145, 32'sd-0.029613735980582357, 32'sd0.20957920167894825, 32'sd-0.0004233254622893255, 32'sd-0.09079672126633945, 32'sd-0.11984588944348173, 32'sd-0.2135118048470314, 32'sd-0.08504161905180467, 32'sd0.12958806740523798, 32'sd0.07948397481011715, 32'sd0.07194277003258091, 32'sd0.12272760419109706, 32'sd0.05382273113860921, 32'sd-0.06821176928930969, 32'sd-0.0674804148411691, 32'sd0.025297265235225713, 32'sd-0.052294622707003004, 32'sd0.030542165727362285, 32'sd-0.041801132877809774, 32'sd-0.005690316545636119, 32'sd-0.12256732629135392, 32'sd-0.009360882004979035, 32'sd0.02994556118103205, 32'sd0.012590886163716708, 32'sd-0.08738191042599257, 32'sd-0.19408014866805712, 32'sd0.03284246488351011, 32'sd0.13447965860319525, 32'sd0.06238212235055917, 32'sd0.15726214045951956, 32'sd0.1848481194447359, 32'sd0.09961378408415249, 32'sd-0.03259423176599222, 32'sd-0.06680540964689669, 32'sd-0.18018607542926052, 32'sd-0.0674462768151522, 32'sd0.04894567311217062, 32'sd-0.004876032989644317, 32'sd0.0881326362835792, 32'sd-0.08636131330295194, 32'sd0.09420085788276994, 32'sd0.13553952663614863, 32'sd0.0942789285183247, 32'sd-0.052604330025761106, 32'sd0.08605640121115284, 32'sd-0.019111974240773988, 32'sd0.07446361413369404, 32'sd-0.030756332386025584, 32'sd-0.08101830916866047, 32'sd-0.029627506547462584, 32'sd0.008198206117004255, 32'sd-0.08446155813461784, 32'sd-0.02169914682691266, 32'sd-0.07144406925956373, 32'sd-0.022338407525512402, 32'sd0.010650386271844229, 32'sd0.13019474281329613, 32'sd0.05813451918646359, 32'sd0.02131164164424324, 32'sd-4.4795200561454726e-05, 32'sd0.06753834079890011, 32'sd0.06821338763924242, 32'sd0.0515214021596737, 32'sd0.0017087536898290794, 32'sd-0.045270941040227344, 32'sd0.007535715567719803, 32'sd0.06552551572741494, 32'sd0.10672172576924402, 32'sd0.1297799579670564, 32'sd0.13126009653888185, 32'sd0.19557987962799903, 32'sd0.017128382584619153, 32'sd0.09558863235097952, 32'sd0.06721632126471964, 32'sd-0.13895584387266302, 32'sd0.00715660357502558, 32'sd0.025441311161423893, 32'sd-0.028941672246629416, 32'sd0.038424563970570286, 32'sd-0.032866129438305816, 32'sd0.0027577296267104453, 32'sd0.026471484444128824, 32'sd-0.11248189169649976, 32'sd0.054757637712210476, 32'sd-0.06745599566276529, 32'sd0.041007297915060865, 32'sd0.07668108175897465, 32'sd0.033320556872456976, 32'sd0.11029149168132486, 32'sd0.08849337223905814, 32'sd0.030991018235493904, 32'sd0.002449931728219725, 32'sd-0.007660742899897489, 32'sd0.10687968424646818, 32'sd-0.012187781876110946, 32'sd0.06323089742013448, 32'sd0.1738954548165626, 32'sd0.09916043520401423, 32'sd0.03211265142753031, 32'sd-0.003688521630635407, 32'sd0.061055205393044654, 32'sd-0.0373723671842662, 32'sd0.14150174798569326, 32'sd-0.011834376773777173, 32'sd-0.05055727603777096, 32'sd-0.06277754872504697, 32'sd0.041498820595543794, 32'sd-0.08305383509670293, 32'sd0.037858241446973626, 32'sd-0.035485826226967006, 32'sd-0.1099509247662781, 32'sd-0.0067651857957923755, 32'sd-0.03207377238066825, 32'sd0.11598939626347968, 32'sd0.07636715825003998, 32'sd-0.002281498475825934, 32'sd0.11936809128427507, 32'sd-0.10175120377094793, 32'sd-0.16115456414895873, 32'sd-0.1865920257412887, 32'sd-0.06220467669661932, 32'sd-0.002607002164555132, 32'sd0.11708175384909067, 32'sd0.07245546464533088, 32'sd-0.0007573579235621884, 32'sd0.0572952948646374, 32'sd-0.10117588832150573, 32'sd-0.0139251653499204, 32'sd-0.05726354647194117, 32'sd-0.06270710069613597, 32'sd0.01635731408854236, 32'sd-0.11959094711617266, 32'sd-0.08164536883310343, 32'sd-0.03757693223834474, 32'sd-0.012273067532314408, 32'sd-0.03236646977032619, 32'sd0.09898793133098925, 32'sd-0.12776828897624407, 32'sd-0.19488887308651048, 32'sd-0.11742498640683104, 32'sd-0.017054738298794503, 32'sd0.0270090009258096, 32'sd0.041573356633747865, 32'sd-0.012275978143807365, 32'sd0.10413651414323995, 32'sd0.02691724013716569, 32'sd-0.07398387969973964, 32'sd-0.18861916998963701, 32'sd0.04811829748808845, 32'sd0.17381870958563098, 32'sd0.24377719657459893, 32'sd0.06572070500160662, 32'sd0.10685240343919905, 32'sd-0.004225735489024251, 32'sd-0.07486809521694772, 32'sd-0.03597670091548317, 32'sd0.011361080429515358, 32'sd0.10310036118079771, 32'sd-0.06400034777134772, 32'sd-0.0832615105718972, 32'sd-0.007369307906231022, 32'sd0.007061074711744101, 32'sd0.0165488788890691, 32'sd-0.04680909495166228, 32'sd-0.04509157213498814, 32'sd-0.03617475107405038, 32'sd-0.15161667563354517, 32'sd-0.0672657099119287, 32'sd0.020158037236537005, 32'sd-0.0696062013058896, 32'sd-0.06092109296166137, 32'sd-0.15416022811852723, 32'sd-0.010311630402122435, 32'sd-0.11745292912637893, 32'sd-0.19239038264620142, 32'sd-0.15415401721723848, 32'sd-0.06182289035565823, 32'sd0.025373743457958224, 32'sd0.10160499230481068, 32'sd0.114661990800824, 32'sd-0.023031694276950742, 32'sd-0.0051332691483582825, 32'sd0.07470095068996574, 32'sd-0.08787158313595489, 32'sd0.021166852506022935, 32'sd0.0804667440795554, 32'sd0.017240712269998012, 32'sd-0.07141073273815549, 32'sd0.07084109954952932, 32'sd-0.04748741532757734, 32'sd0.01595867697330968, 32'sd0.07362027299442246, 32'sd0.1034749678223385, 32'sd0.028726782459951795, 32'sd0.022746338710788273, 32'sd-0.018378892945482363, 32'sd0.002513863180344521, 32'sd-0.066851985730894, 32'sd-0.03484655139614449, 32'sd-0.09056990704814638, 32'sd-0.08006359451102435, 32'sd-0.027307810151950267, 32'sd-0.0430576337351395, 32'sd-0.11342212744321598, 32'sd-0.025573628102333445, 32'sd0.06424243593090712, 32'sd0.20048688763030362, 32'sd0.12664765985299145, 32'sd-0.0748670086988383, 32'sd-0.02122141627503786, 32'sd-0.0552007071829266, 32'sd-0.16294152291008945, 32'sd-0.03113495561719595, 32'sd0.05562590262118013, 32'sd0.06321436568372728, 32'sd0.07248098382414613, 32'sd0.004047931285687312, 32'sd0.041700810560038826, 32'sd3.5879311581023057e-116, 32'sd-0.028080815897925465, 32'sd0.014565440404333998, 32'sd-0.11417131892990262, 32'sd-0.061831446944879506, 32'sd0.043154573833927075, 32'sd-0.029254152819427833, 32'sd-0.14077919803226305, 32'sd-0.09908505458689616, 32'sd-0.18785101447885752, 32'sd-0.1283076953641772, 32'sd0.022751417821630853, 32'sd-0.07983964858398444, 32'sd-0.05754296758886614, 32'sd-0.0647748486134287, 32'sd0.08616987893442589, 32'sd0.10547822800031535, 32'sd0.07627277937387224, 32'sd0.14795866523226422, 32'sd-0.11865507095903788, 32'sd-0.11210574338128797, 32'sd-0.03088356567867198, 32'sd-0.13339546447173048, 32'sd-0.0725467050097408, 32'sd-0.012135802783712672, 32'sd0.05473014814747348, 32'sd-0.02745014415712942, 32'sd0.01531405247373159, 32'sd-0.05692421860146428, 32'sd0.053170085428857775, 32'sd-0.08096845924149183, 32'sd0.02093634267639472, 32'sd-0.1679049702489272, 32'sd-0.018972112495501174, 32'sd0.0675262650866686, 32'sd0.032862563032111027, 32'sd0.025200911519239713, 32'sd-0.13127645553791886, 32'sd-0.09561360163943335, 32'sd-0.05253292818382566, 32'sd-0.1252151966639155, 32'sd-0.09114431508326629, 32'sd-0.00723707027489077, 32'sd0.12308788864841513, 32'sd0.0673611433568421, 32'sd0.12010375722411375, 32'sd0.08892578578583105, 32'sd-0.059167410654354685, 32'sd-0.09688651276864056, 32'sd-0.03205013717142873, 32'sd-0.0776087414655894, 32'sd-0.19433747381943603, 32'sd-0.008090079000109898, 32'sd0.1099989686355251, 32'sd0.04352554528307571, 32'sd-0.04351736491373133, 32'sd-0.003973234232622506, 32'sd0.03363568339320753, 32'sd-0.05393441976521297, 32'sd0.036853448104947784, 32'sd-0.22696484220371888, 32'sd0.030368564823266365, 32'sd-0.04889328139400101, 32'sd0.05544594998579456, 32'sd-0.10375802098190154, 32'sd-0.12036077837401776, 32'sd-0.015315880603300433, 32'sd-0.0024590739623868364, 32'sd-0.06521960793380069, 32'sd0.06440228059608888, 32'sd0.07339253519261173, 32'sd-0.012500500568931623, 32'sd0.05617904813855563, 32'sd-0.017709322105452525, 32'sd0.015322977606680836, 32'sd0.011850084630502666, 32'sd-0.13556849748921979, 32'sd-0.01183032473000003, 32'sd-0.03343906500751721, 32'sd-0.03318041174557061, 32'sd-0.06142860646939086, 32'sd-0.016831381900166253, 32'sd-0.06237521282016511, 32'sd-0.005957201580190049, 32'sd1.5022506688646668e-119, 32'sd-0.01101276610929578, 32'sd0.03149369611771407, 32'sd-0.03535476518526822, 32'sd-0.19742901700415486, 32'sd-0.12263555525226308, 32'sd-0.04128538637864462, 32'sd0.053752375559090224, 32'sd-0.0767626552432176, 32'sd-0.02088166703179495, 32'sd-0.040515176559030086, 32'sd0.04209111737266801, 32'sd-0.031330111857996244, 32'sd-0.12863226914793535, 32'sd-0.08244344165887427, 32'sd0.01333904625738535, 32'sd0.01503949134888141, 32'sd-0.020390537739477098, 32'sd-0.05322179781258868, 32'sd-0.08088479918763417, 32'sd-0.003634141169661785, 32'sd-0.0625166280451232, 32'sd-0.05261633398653644, 32'sd-0.05796727116483646, 32'sd0.10198964788154391, 32'sd0.0912906870887376, 32'sd0.03606834439718506, 32'sd-0.009383572690251168, 32'sd-0.04622499790162779, 32'sd-0.012620799523128393, 32'sd-0.1111246695154466, 32'sd0.03420481949503518, 32'sd0.00370752144681512, 32'sd-0.00059526999353276, 32'sd-0.05849439951601272, 32'sd-0.0977590183361156, 32'sd0.020436842246377127, 32'sd0.07210811477768816, 32'sd0.029565012925378442, 32'sd0.09175874476710492, 32'sd0.04527933376076036, 32'sd-0.08429343676547724, 32'sd-0.019665766234205306, 32'sd-0.12942193756098905, 32'sd0.0520632148903603, 32'sd-0.018751944172977084, 32'sd-0.08616263574293574, 32'sd0.02789505781972483, 32'sd0.0008224962062359556, 32'sd-0.020318203421206556, 32'sd-0.05580883735003104, 32'sd0.03370508042016327, 32'sd0.07865937793354569, 32'sd0.029740812768287144, 32'sd-0.06575665427579998, 32'sd-0.040326277390543466, 32'sd-0.005521018710618969, 32'sd-0.009191098956716897, 32'sd-0.04414711282035139, 32'sd0.01598494416645704, 32'sd0.03358184591684551, 32'sd-0.07906442810267315, 32'sd-0.10041918244585957, 32'sd-0.019070499351447376, 32'sd-0.012600297910664374, 32'sd-0.00024272315364994064, 32'sd0.12125551318113124, 32'sd0.06811614758401562, 32'sd0.09702502441684924, 32'sd-0.054906014257091025, 32'sd0.01067924701856264, 32'sd-0.13669684386036532, 32'sd-0.0754067449925953, 32'sd-0.05196873327255178, 32'sd-0.020330915283055587, 32'sd0.010181383452637539, 32'sd-0.041455335819483755, 32'sd0.03932255657566413, 32'sd0.029268165433290635, 32'sd-0.0655956641273579, 32'sd0.04317151231997045, 32'sd-0.13993036959849364, 32'sd-0.023650775500909993, 32'sd-0.0013369443233122997, 32'sd3.735409574006463e-125, 32'sd-0.023469135932131825, 32'sd-0.05669717631531677, 32'sd-0.057487355304635904, 32'sd-0.08188910972489002, 32'sd-0.043874841345563714, 32'sd-0.023501453536181726, 32'sd-0.024282908473992944, 32'sd-0.028350874476674313, 32'sd0.03542135662891115, 32'sd0.08629402262377285, 32'sd0.08088884773606414, 32'sd-0.014742168125785302, 32'sd0.02246990366950434, 32'sd-0.0672241164097831, 32'sd0.006806325102236616, 32'sd-0.08750281457077766, 32'sd0.020853183217841922, 32'sd-0.06309798126620408, 32'sd0.044980962429079036, 32'sd0.06357970348856024, 32'sd0.07381863236636717, 32'sd0.06979089600363803, 32'sd0.03616579282441905, 32'sd0.040738642362739205, 32'sd0.02658172363615542, 32'sd-0.03436241000152323, 32'sd3.435683267134126e-123, 32'sd2.569071931427491e-114, 32'sd-4.7098700924617755e-115, 32'sd0.020506512424216, 32'sd-0.0062652794057216086, 32'sd-0.0027001381724863324, 32'sd0.02271072854855757, 32'sd-0.02119624303814444, 32'sd-0.022157198785326796, 32'sd-0.027610107087623598, 32'sd-0.01802829652546915, 32'sd0.10464519708199092, 32'sd0.0007891018122831745, 32'sd0.04976733033194774, 32'sd-0.15336337898935298, 32'sd0.015826514580891064, 32'sd0.04587369864101176, 32'sd0.004614359772512115, 32'sd-0.06621740875216293, 32'sd-0.09675898967832053, 32'sd0.09020659243669904, 32'sd0.08957991130113763, 32'sd-0.07687196728233975, 32'sd0.02510661797140661, 32'sd-0.03496807475204301, 32'sd0.0015876777940926944, 32'sd0.03730971749694086, 32'sd-0.024750893336968924, 32'sd1.0282181711194434e-121, 32'sd-1.604560646209521e-116, 32'sd1.0891985612166227e-115, 32'sd0.07457855504087026, 32'sd0.009781560126295207, 32'sd0.05584535954435637, 32'sd0.0068235593330380675, 32'sd0.01290279485300493, 32'sd-0.0840749201388867, 32'sd0.0775963964105408, 32'sd0.08512480874428885, 32'sd-0.012075232348847323, 32'sd0.07683072320371902, 32'sd0.06930407010192675, 32'sd-0.10702715626188104, 32'sd0.09229306450455549, 32'sd-0.1326797638274075, 32'sd-0.005479944628601062, 32'sd-0.06696888976803145, 32'sd0.021897079820068284, 32'sd-0.08534682832912548, 32'sd-0.012617778451602717, 32'sd-0.05000751169975308, 32'sd-0.05950335607626233, 32'sd0.022604485667423582, 32'sd-0.029085622320598716, 32'sd0.01296904668645139, 32'sd-0.02523200372861747, 32'sd-1.215382575637411e-121, 32'sd-2.5612163960484317e-126, 32'sd-1.9064221499762266e-126, 32'sd-4.5347712170156194e-122, 32'sd-0.02638872447125133, 32'sd0.06713260558884909, 32'sd-0.11171452063589278, 32'sd-0.1408979413207852, 32'sd0.009987062186099517, 32'sd0.05077174872873552, 32'sd0.09544159612844359, 32'sd0.08326713448734281, 32'sd-0.042009379763180005, 32'sd0.04996672016815451, 32'sd-0.016152727389672404, 32'sd0.03086625467887363, 32'sd-0.039374886955457926, 32'sd0.0350026531299739, 32'sd0.11364343582039863, 32'sd-0.007019585003617355, 32'sd-0.0381701017098634, 32'sd0.011435912029475323, 32'sd-0.08888385048498566, 32'sd0.020718145931726804, 32'sd0.005058454221669133, 32'sd-0.08312455969582207, 32'sd0.0447696304028282, 32'sd-1.0953596122104658e-122, 32'sd3.3844920827206937e-122, 32'sd-8.207095975497829e-115, 32'sd-3.241133063576825e-123, 32'sd-6.843264710774564e-126, 32'sd-2.232956113432609e-114, 32'sd-0.05078221960755738, 32'sd0.005225264495070136, 32'sd-0.036536817749118676, 32'sd-0.019863417303365383, 32'sd-0.03983968247938245, 32'sd-0.01130303303138162, 32'sd-0.0668277222312345, 32'sd-0.04647408850017563, 32'sd-0.04853439557676037, 32'sd0.04292327581968879, 32'sd0.051723391579177186, 32'sd-0.037923654494883115, 32'sd-0.033952765590786714, 32'sd0.021675221580485217, 32'sd0.08632408822518481, 32'sd0.11364729980038114, 32'sd-0.028179283965375397, 32'sd0.02179296636815062, 32'sd0.0760108015738733, 32'sd0.041750034828597994, 32'sd1.3487511980681717e-127, 32'sd-8.191144966851687e-125, 32'sd-3.871187816558203e-125, 32'sd1.3155015455430203e-123},
        '{32'sd-1.6305679394160379e-115, 32'sd3.262896530303248e-121, 32'sd-1.1850124239322112e-126, 32'sd1.316909026572848e-119, 32'sd-6.797007226916824e-119, 32'sd-3.7935495989641046e-125, 32'sd8.341384346685801e-118, 32'sd-8.193258874223442e-126, 32'sd1.9427157582554277e-125, 32'sd1.9833069212603385e-117, 32'sd2.4566890505148638e-126, 32'sd6.934454494314551e-123, 32'sd0.002659703255841903, 32'sd0.06081752878159667, 32'sd0.02628625140509112, 32'sd0.04295329990079857, 32'sd1.6793895181911925e-123, 32'sd-1.7085620322791775e-129, 32'sd2.4535480544184838e-123, 32'sd-1.9906257457014068e-117, 32'sd9.946192621017864e-128, 32'sd-1.0438166454481254e-120, 32'sd1.6987565483592046e-114, 32'sd4.1283811149778775e-123, 32'sd-1.8258247402850012e-117, 32'sd4.481246006309072e-123, 32'sd-6.044058877059442e-122, 32'sd7.616769234984007e-122, 32'sd-1.0091220394056267e-114, 32'sd-9.279813100242743e-121, 32'sd1.6213087810175605e-115, 32'sd-5.893999991721722e-125, 32'sd0.10391186389365871, 32'sd3.020320482727496e-05, 32'sd-0.034480619612111574, 32'sd-0.011043288331713618, 32'sd0.06536262491080848, 32'sd-0.011449629514706697, 32'sd-0.025104529391680782, 32'sd0.0056177254710433906, 32'sd0.023091438033136936, 32'sd0.025833735578599977, 32'sd-0.047928836505385104, 32'sd-0.058715724365771986, 32'sd0.13892956703067988, 32'sd0.0729406843095391, 32'sd0.10098094824168558, 32'sd0.15630693554381334, 32'sd0.10641823848165467, 32'sd0.11415103240139897, 32'sd0.14924729678497137, 32'sd0.06422505913894706, 32'sd-3.520443210252231e-119, 32'sd-3.3820988740053853e-116, 32'sd-2.341606753460946e-118, 32'sd-6.457639915700995e-126, 32'sd-1.0888660542499931e-119, 32'sd-2.1670384950717705e-120, 32'sd0.1309479642827972, 32'sd0.09486891563616953, 32'sd0.02787836727703533, 32'sd0.06655838525206835, 32'sd0.047937252279139225, 32'sd-0.09555800459783072, 32'sd0.01648124916316789, 32'sd-0.06778278912031369, 32'sd-0.10558973458175698, 32'sd0.10882759388202773, 32'sd0.040952143091513904, 32'sd-0.04386134564099231, 32'sd0.00942712470070578, 32'sd-0.07451096533742349, 32'sd-0.07639907345089952, 32'sd0.002162490347871043, 32'sd0.08746426052119755, 32'sd0.037631614968462214, 32'sd0.005270906442340591, 32'sd0.11862106542767972, 32'sd0.13962030445756207, 32'sd0.1099067265444561, 32'sd-0.02266474282915699, 32'sd0.1141615958932855, 32'sd-3.7628987813682086e-122, 32'sd-2.116734503484597e-121, 32'sd1.0804417023043984e-122, 32'sd7.77313127377808e-125, 32'sd0.11261550730162094, 32'sd-0.03368647802083401, 32'sd0.02366564523805479, 32'sd-0.017909749471373124, 32'sd-0.00808003058475922, 32'sd-0.0263966849297896, 32'sd0.04859255683554444, 32'sd-0.007211314481225366, 32'sd-0.04830352898946094, 32'sd0.053166832814781184, 32'sd0.03928288839151286, 32'sd-0.022583744838943452, 32'sd-0.05408866899192359, 32'sd-0.11872987523371992, 32'sd-0.03577169732106974, 32'sd-0.005275568311293342, 32'sd0.03336204165558193, 32'sd0.01990404502409912, 32'sd0.05563086807515505, 32'sd0.001857987428506096, 32'sd0.06034274438324897, 32'sd0.051526777277835625, 32'sd0.023091375439006617, 32'sd0.0588786121948725, 32'sd0.03922852857675593, 32'sd-1.936576779537769e-125, 32'sd-4.7335468109648e-115, 32'sd0.06084243376142057, 32'sd0.06557124194893076, 32'sd-0.010682006577805984, 32'sd0.09297990174279028, 32'sd0.06956165067011032, 32'sd-0.03599747718655961, 32'sd-0.009051822017380773, 32'sd0.04552290892392202, 32'sd-0.03395791509620998, 32'sd-0.11798810368090057, 32'sd0.1136743173064616, 32'sd-0.0026445028576723853, 32'sd0.07486799322239782, 32'sd-0.0624531316365028, 32'sd-0.08536278487566723, 32'sd0.032133948396327695, 32'sd0.018221711543641664, 32'sd0.014023552468100078, 32'sd0.07412992508497876, 32'sd0.09009888987906925, 32'sd0.08098405352083751, 32'sd-0.09489328152656731, 32'sd0.011611024125239356, 32'sd0.08013530666553348, 32'sd-0.008684087291280734, 32'sd-0.05011222912667007, 32'sd0.028581909536957006, 32'sd1.1346857667375963e-119, 32'sd0.0321526640725093, 32'sd0.015834006138608876, 32'sd-0.09297221307981875, 32'sd-0.012470446213867248, 32'sd-0.05963296086852195, 32'sd0.01040281591395652, 32'sd0.042781677076894155, 32'sd0.05371298662237774, 32'sd-0.009200093051772978, 32'sd-0.0479061027123393, 32'sd0.15708415398586648, 32'sd0.12672063737606037, 32'sd0.10583998412591358, 32'sd-0.03289274466133309, 32'sd0.019167725165985635, 32'sd0.09186488145569223, 32'sd0.1646077529679484, 32'sd0.05307778051863334, 32'sd0.10711269349369328, 32'sd-0.017393030560177287, 32'sd0.015251185949368667, 32'sd-0.016652376912200187, 32'sd-0.03414091053665946, 32'sd0.09867244999506188, 32'sd-0.06608874566709605, 32'sd0.046863813574377876, 32'sd0.07374901423309, 32'sd-1.4333667669319225e-124, 32'sd0.02553012849830847, 32'sd0.016211715356736774, 32'sd0.10452960701551067, 32'sd-0.04821870583032286, 32'sd-0.030597483827037926, 32'sd-0.04141199688677672, 32'sd-0.000370282625777004, 32'sd-0.016085901070641364, 32'sd0.049610329477101346, 32'sd-0.008062103116193074, 32'sd0.10525324859592175, 32'sd0.09131624203349774, 32'sd0.04846070819617413, 32'sd-0.036970792229755516, 32'sd0.005280964956708443, 32'sd-0.0072409971150536765, 32'sd0.06146438997552029, 32'sd0.08278070179566407, 32'sd0.12955860819011583, 32'sd0.009898242943828201, 32'sd0.021732869814149788, 32'sd2.0232618320890845e-05, 32'sd-0.006124360489938324, 32'sd0.02960059199572859, 32'sd0.0722197325831823, 32'sd0.0013005059028717014, 32'sd-0.008318339254143183, 32'sd0.10047055599511098, 32'sd0.09608380830649288, 32'sd0.0059873079990410425, 32'sd-0.07365540378312407, 32'sd0.06375851780485825, 32'sd0.07754171827911811, 32'sd0.09272393941057751, 32'sd0.04477610491856135, 32'sd0.043396144052477034, 32'sd-0.08481283894209535, 32'sd-0.06614235559684294, 32'sd-0.09949616915510698, 32'sd-0.1359088665640915, 32'sd0.014762880660823374, 32'sd0.007693144766521407, 32'sd-0.007142224839509737, 32'sd-0.0777700823335914, 32'sd0.03405223970264927, 32'sd0.11378148728430851, 32'sd0.03494846351892655, 32'sd0.04734003388026303, 32'sd0.01920125681842002, 32'sd0.09791866137712052, 32'sd0.08135578069793684, 32'sd0.11814732540362084, 32'sd0.05738450034525259, 32'sd0.11538459881838661, 32'sd0.08146253479544395, 32'sd0.06811172873003347, 32'sd0.06353092440244232, 32'sd-0.08668980058378992, 32'sd0.09585053008601951, 32'sd0.02497394097446148, 32'sd0.04233429613662946, 32'sd0.04768424643178782, 32'sd-0.029601915293064076, 32'sd-0.008507916191371999, 32'sd-0.030036562383121437, 32'sd-0.07133347315404226, 32'sd-0.12490696910176895, 32'sd-0.05985420091362193, 32'sd0.016740128146905384, 32'sd-0.05948884907562302, 32'sd0.0601868393572481, 32'sd0.014656059277370972, 32'sd0.04715553043636661, 32'sd0.041634189348792934, 32'sd0.18121108203105574, 32'sd0.10275687081200413, 32'sd0.03023186233306405, 32'sd0.18098597812148357, 32'sd0.14436103311832982, 32'sd0.16072035284532746, 32'sd0.03902343650533032, 32'sd0.02050533261976063, 32'sd-0.035182706941005615, 32'sd-0.01805716172442015, 32'sd0.05013851485339537, 32'sd0.09879703792387344, 32'sd0.12727260129421694, 32'sd-0.018060412263272988, 32'sd-0.004591256250315773, 32'sd-0.07377603330363083, 32'sd-0.09993735279227539, 32'sd-0.2060169367605705, 32'sd-0.04838037033159218, 32'sd-0.025649637273893123, 32'sd-0.0034047789198326872, 32'sd-0.12665830008591977, 32'sd-0.07550278742085632, 32'sd-0.06470989320525086, 32'sd0.03529651575038473, 32'sd-0.16585027484698203, 32'sd0.08046636199261155, 32'sd0.018024032747885405, 32'sd0.07173839829823356, 32'sd-0.03370532432272825, 32'sd0.10188827984061165, 32'sd0.06151431180809586, 32'sd0.13285581681257713, 32'sd-0.03546982699750082, 32'sd0.06583987494568438, 32'sd0.008357275045202174, 32'sd-0.009657428570056966, 32'sd0.06469118256580775, 32'sd0.011112052254729278, 32'sd0.09723006398834537, 32'sd0.11464209246271392, 32'sd-0.0467342316985979, 32'sd-0.11240734609385555, 32'sd-0.015509591794893585, 32'sd-0.09934786138257026, 32'sd-0.1893175814266687, 32'sd0.006707867658938681, 32'sd-0.06371811134234238, 32'sd-0.08265554842367151, 32'sd0.01728750161571665, 32'sd-0.1794223269561958, 32'sd-0.18935408836658263, 32'sd-0.1329786728853591, 32'sd-0.06245933066479284, 32'sd-0.12399201751553018, 32'sd-0.0994190485531444, 32'sd-0.13044317692367968, 32'sd-0.04318465999165261, 32'sd-0.17071758688936983, 32'sd-0.07385098463546093, 32'sd-0.10543056216138968, 32'sd-0.017437275818006904, 32'sd-0.006214034835176472, 32'sd0.07283807077525883, 32'sd0.07053392557528776, 32'sd0.0020375097490141422, 32'sd0.06506696717332301, 32'sd0.0930048672744536, 32'sd0.035727945004230106, 32'sd-0.1236607450339418, 32'sd-0.10107896202310945, 32'sd-0.11374838611064952, 32'sd-0.21667851457826118, 32'sd-0.13643354939433017, 32'sd-0.07821965314793036, 32'sd-0.015058381612713025, 32'sd-0.03708396391488201, 32'sd-0.05132094234344807, 32'sd-0.08306093730347103, 32'sd-0.17799972040581524, 32'sd-0.07828854320341894, 32'sd-0.2880169888824465, 32'sd-0.3203207735457024, 32'sd-0.267301465696564, 32'sd-0.2686002951238078, 32'sd-0.14920323298728758, 32'sd-0.28634392690707744, 32'sd-0.10530885428765198, 32'sd-0.1558636387708897, 32'sd-0.09270781281348774, 32'sd-0.006444004853536246, 32'sd-0.037666862127038056, 32'sd-0.059858978607335044, 32'sd0.02190796399496201, 32'sd0.0408441644341982, 32'sd0.07825053350060228, 32'sd0.03077351297746044, 32'sd-0.10500831607821448, 32'sd-0.10252934871158341, 32'sd-0.1112800684231598, 32'sd-0.04989515593892376, 32'sd-0.09389551101928774, 32'sd0.021135071741692216, 32'sd-0.03442572879833238, 32'sd0.09210879099323739, 32'sd0.013638255284330348, 32'sd-0.05073753182541072, 32'sd-0.14032300993263624, 32'sd-0.07220574460429481, 32'sd-0.1743233453670641, 32'sd-0.3095148537130891, 32'sd-0.11728824418713847, 32'sd-0.13648852472666578, 32'sd-0.2683419723112498, 32'sd-0.2437604216772687, 32'sd-0.2222978381570642, 32'sd-0.06390727831498627, 32'sd-0.048005013583799536, 32'sd-0.023792602991955767, 32'sd0.020090535978402005, 32'sd-0.002942112450087557, 32'sd0.036503088568710186, 32'sd0.032837370381893764, 32'sd0.061774382956709006, 32'sd0.015435432906878268, 32'sd-0.2041758478216724, 32'sd-0.09208507570028722, 32'sd-0.01811713274743047, 32'sd0.06957231039843528, 32'sd-0.008814706844066118, 32'sd0.02161217639496003, 32'sd0.02290197284772227, 32'sd-0.042044182423490783, 32'sd0.12360491793363847, 32'sd0.1656293607656583, 32'sd0.06400258037072065, 32'sd0.1532377748142871, 32'sd-0.016602555283529954, 32'sd-0.025764113741548744, 32'sd-0.08011741416954578, 32'sd-0.06931127422039729, 32'sd-0.14617450759169456, 32'sd-0.16137301541089438, 32'sd-0.1618722554264994, 32'sd-0.13010999259860484, 32'sd0.022068929543819678, 32'sd-0.046358566080194716, 32'sd-0.03621501117623785, 32'sd0.12558650480947342, 32'sd0.09645045183130734, 32'sd-0.018844007864107643, 32'sd0.08288441112497585, 32'sd-0.04787276700010799, 32'sd0.07835606815472428, 32'sd-0.0073926219885740024, 32'sd0.06255299058012036, 32'sd0.05131576526779732, 32'sd0.04950913648775022, 32'sd-0.03336735706232988, 32'sd0.07353584400127583, 32'sd-0.059849376891362535, 32'sd-0.03937641235091845, 32'sd0.06367686633213086, 32'sd0.01745971756825342, 32'sd0.2007968512631392, 32'sd0.0474132677165288, 32'sd0.06680347051730373, 32'sd0.027942898446222688, 32'sd-0.09979361010548367, 32'sd0.019796816821430325, 32'sd-0.07772424260569417, 32'sd-0.09305958594824733, 32'sd-0.14444430610117548, 32'sd-0.030855551181586463, 32'sd0.12191006776920023, 32'sd0.025161000440517715, 32'sd0.11295478177068986, 32'sd0.06411616194556526, 32'sd0.07585130257922286, 32'sd-0.026718624325030457, 32'sd0.04236770717466091, 32'sd0.17885311206979643, 32'sd0.185522438736797, 32'sd0.02919706420491772, 32'sd0.05353215520501845, 32'sd0.08059336916389237, 32'sd-0.03703020351869323, 32'sd-0.09437067558865642, 32'sd-0.0792629869715884, 32'sd-0.028383251409908317, 32'sd0.016086702531543758, 32'sd0.10397375682742534, 32'sd0.014320619289327883, 32'sd0.16063450741059196, 32'sd0.10903147527054527, 32'sd0.1242967517177029, 32'sd-0.0678967028210022, 32'sd-0.03710560538222235, 32'sd0.012877215940352611, 32'sd-0.13258176418368273, 32'sd-0.025068906764183958, 32'sd-0.009818549494066095, 32'sd0.05038445703290595, 32'sd0.09173580920987351, 32'sd0.04428514523380058, 32'sd0.06592028660524343, 32'sd-0.05032199279847595, 32'sd-0.05921381178021754, 32'sd-0.0013037855021706595, 32'sd0.1689482769398362, 32'sd0.08193376576770765, 32'sd-0.004535752458646781, 32'sd0.13607932148833252, 32'sd-0.09670039240634924, 32'sd-0.08095448257557018, 32'sd0.015174140288499015, 32'sd-0.044396464192807204, 32'sd0.17330427681530486, 32'sd0.019658969765603787, 32'sd0.037338355511358584, 32'sd0.01627725269960848, 32'sd-0.007827674428297675, 32'sd0.05462815316325499, 32'sd0.010472733743662187, 32'sd0.036052566965539684, 32'sd0.009904920914813709, 32'sd0.061703509543934255, 32'sd0.10100255507197202, 32'sd0.014696073361590897, 32'sd0.0540028937319327, 32'sd0.012515336463435318, 32'sd-0.08505855745454922, 32'sd-0.007410558976240772, 32'sd-2.676545971227088e-124, 32'sd0.03274248841249448, 32'sd-0.18042825648417152, 32'sd0.05070521044545684, 32'sd0.1580453405470052, 32'sd0.08140023666101805, 32'sd0.05029882954386691, 32'sd0.09757200485441742, 32'sd-0.012119189630326644, 32'sd0.023318771623848617, 32'sd-0.06912346267435243, 32'sd-0.037127711439930974, 32'sd0.041851830468942926, 32'sd-0.009438842315755562, 32'sd-0.1633552889941056, 32'sd-0.058543107446053295, 32'sd-0.0074616449429980684, 32'sd0.08153578703690473, 32'sd0.08560719742473256, 32'sd0.0795510712453848, 32'sd0.09710694761090093, 32'sd0.1192430219790896, 32'sd0.06838361111328455, 32'sd-0.060566588492729515, 32'sd-0.0780712805303755, 32'sd-0.18961005224149674, 32'sd-0.001661937009881949, 32'sd0.05841140636217389, 32'sd-0.012760368422138195, 32'sd0.07688055891980963, 32'sd-0.024611322793960826, 32'sd0.0751214748410229, 32'sd-0.056028322480303705, 32'sd0.07946320596540042, 32'sd0.12421248319106191, 32'sd0.04889587886163417, 32'sd0.03398846392579274, 32'sd-0.031043279425424026, 32'sd-0.06888691171599895, 32'sd-0.03711794252995126, 32'sd0.05348018061770138, 32'sd-0.20016868563228252, 32'sd-0.10533892321830504, 32'sd0.02301754393095732, 32'sd0.04324888477489255, 32'sd0.04044304478896472, 32'sd0.06857671705856663, 32'sd0.14275515079917847, 32'sd0.16772856461693553, 32'sd0.14066364192921085, 32'sd-0.05767159560127233, 32'sd-0.06802039322513567, 32'sd-0.06194627323864617, 32'sd-0.03999578103062972, 32'sd0.052392580828951485, 32'sd0.08460777070901561, 32'sd0.01604819002878796, 32'sd-0.06705045022540396, 32'sd-0.054021905163972095, 32'sd0.02559369917028386, 32'sd-0.0026595126461199325, 32'sd-0.15745992447275042, 32'sd-0.01777352316508441, 32'sd-0.03503692971146642, 32'sd-0.01266863552881179, 32'sd-0.04106920100398325, 32'sd-0.0314425842169792, 32'sd0.03198121954750074, 32'sd0.006633441103645495, 32'sd-0.041457919511650704, 32'sd0.012675195408063139, 32'sd0.012157261546957331, 32'sd0.00858306776489477, 32'sd0.14505178402964453, 32'sd0.16980770942407666, 32'sd0.11006998698231048, 32'sd0.08722719614905218, 32'sd0.04752941825081611, 32'sd0.01907256529591989, 32'sd0.11200057535849217, 32'sd0.018583716759762163, 32'sd0.054446113430889585, 32'sd0.11451514696360629, 32'sd0.02697597576239449, 32'sd6.259380426377918e-124, 32'sd-0.04274938739075668, 32'sd0.06906135900652735, 32'sd0.017152445693371567, 32'sd0.03239288515431765, 32'sd-0.11749163009675546, 32'sd-0.06401695128321906, 32'sd-0.04341644012907782, 32'sd-0.02994807637694468, 32'sd-0.037833789672368855, 32'sd0.08220441528836454, 32'sd0.03133264074702722, 32'sd-0.08984839559802876, 32'sd0.1195348658179755, 32'sd-0.062175253221990634, 32'sd-0.035190102225875965, 32'sd-0.05561416190020448, 32'sd0.16409794614256276, 32'sd-0.036497948826200936, 32'sd0.06320859598796959, 32'sd-0.0009885568790147972, 32'sd0.005558228797137223, 32'sd0.06793492521109734, 32'sd-0.17271005085331909, 32'sd-0.037383478495139705, 32'sd-0.10362424170878957, 32'sd0.04914442781617605, 32'sd0.019699220338508846, 32'sd0.011328426771113122, 32'sd-0.009936969503706573, 32'sd0.0695064506969163, 32'sd0.07682431635640438, 32'sd0.004682273513827543, 32'sd-0.026575411843124175, 32'sd1.6831569484445656e-05, 32'sd-0.05260407717035796, 32'sd-0.029630661718912175, 32'sd-0.022398760747894007, 32'sd0.15258283362023514, 32'sd0.04308721301811584, 32'sd-0.04268117415130759, 32'sd0.04037684003098112, 32'sd0.022792858956274527, 32'sd-0.001148164924871062, 32'sd0.11387738092375471, 32'sd0.17656329916765173, 32'sd0.05946684041231447, 32'sd-0.06385785186470602, 32'sd-0.0263730515473063, 32'sd-0.018893292433496564, 32'sd-0.15625455744747802, 32'sd-0.22366059571146066, 32'sd-0.043836761111633225, 32'sd-0.058562319695057215, 32'sd0.06912383979139931, 32'sd0.04763145504934969, 32'sd-0.03206075467507787, 32'sd-0.10029073059092485, 32'sd-0.007768017187627891, 32'sd-0.01424058238182652, 32'sd0.06864437861303059, 32'sd0.0028405047042495556, 32'sd-0.0667118915504095, 32'sd-0.027702628265882785, 32'sd0.011975086129597527, 32'sd0.05575915763259183, 32'sd0.07519252754146735, 32'sd0.11209352031127784, 32'sd0.09908537525620603, 32'sd0.12685700516233625, 32'sd0.11221136064188555, 32'sd0.19007093700661473, 32'sd0.10251772743890403, 32'sd0.12123258161669132, 32'sd-0.19404592302821735, 32'sd0.032818676738992504, 32'sd-0.09692671087568674, 32'sd0.020775589287251362, 32'sd-0.14232210428412603, 32'sd-0.08443517661024906, 32'sd-0.10221366501875791, 32'sd-0.09209679008630152, 32'sd-0.07155752101524386, 32'sd0.06804868261592782, 32'sd-2.544463451323094e-125, 32'sd0.043631846999407635, 32'sd-0.05317029642515282, 32'sd0.008340145992933206, 32'sd0.08703439024896704, 32'sd0.03676601622338374, 32'sd-0.04839517141495123, 32'sd-0.053495742842655236, 32'sd0.06452419346097428, 32'sd0.004814484331916046, 32'sd0.04400208770550696, 32'sd0.027014945732569472, 32'sd0.08836177422062341, 32'sd0.05503039275465477, 32'sd0.17102310702455542, 32'sd0.13145707837573653, 32'sd-0.03866877383606115, 32'sd-0.1003168643391728, 32'sd-0.02181295288389321, 32'sd-0.04984578217782041, 32'sd-0.05639847105398855, 32'sd-0.11366238468423981, 32'sd-0.037841791906480654, 32'sd0.008625165570988873, 32'sd-0.03368898830176158, 32'sd-0.04035565621004621, 32'sd0.022230076736951945, 32'sd2.732840196164927e-120, 32'sd-2.3126364056152705e-124, 32'sd-6.688444238084539e-124, 32'sd-0.09390543796590593, 32'sd0.10516830949748321, 32'sd0.05886109961194147, 32'sd-0.062242080454955925, 32'sd-0.04624000362176439, 32'sd0.02532408603167985, 32'sd-0.007964200695160364, 32'sd-0.024832194318218037, 32'sd0.012816564028794627, 32'sd0.07426003140186527, 32'sd-0.038695376376417095, 32'sd-0.02784827187315716, 32'sd0.01656087731145468, 32'sd-0.023312362599373568, 32'sd-0.20938412764675038, 32'sd-0.08828413384170444, 32'sd-0.17846784667442095, 32'sd-0.06118947336852826, 32'sd-0.03516731887265249, 32'sd0.0313980622874887, 32'sd-0.06160134086257856, 32'sd0.0907398588925649, 32'sd0.04152194422561691, 32'sd0.032720848999166094, 32'sd-0.041087469638379254, 32'sd-5.076276939689512e-115, 32'sd2.601798692358289e-126, 32'sd1.3571513772297438e-122, 32'sd0.011312961767343022, 32'sd0.0323388735074885, 32'sd-0.06108829402888972, 32'sd0.033369949937547425, 32'sd-0.06090833423915551, 32'sd-0.0035548285304217012, 32'sd-0.04716182779388154, 32'sd0.08768823428521089, 32'sd-0.12480298447262177, 32'sd-0.1587996735859645, 32'sd-0.05474750024992493, 32'sd-0.10796723871792487, 32'sd0.03501231855947515, 32'sd0.037053732347450595, 32'sd-0.13343245616939095, 32'sd-0.11548099942434491, 32'sd-0.05050160576902309, 32'sd0.08865223527569442, 32'sd0.005763766659367664, 32'sd-0.04577848735741416, 32'sd0.06996737314799639, 32'sd0.04343640190110834, 32'sd0.001769173272674298, 32'sd-0.012527549826065354, 32'sd0.017260189872458004, 32'sd6.232697421074581e-116, 32'sd2.5034815123178444e-122, 32'sd1.7315060875196545e-125, 32'sd-2.556360015150558e-126, 32'sd0.09105507955644207, 32'sd-0.04446770799705949, 32'sd0.019911099751072844, 32'sd0.02118734781054412, 32'sd-0.019007896333811343, 32'sd-0.05349011455590326, 32'sd0.029974901609360245, 32'sd0.06916621320182437, 32'sd-0.023902879973642627, 32'sd0.023766748048723713, 32'sd0.08263145023553611, 32'sd0.010523467329699542, 32'sd-0.04577051704485288, 32'sd-0.07411815457098367, 32'sd0.0398997625016468, 32'sd0.02162808065407712, 32'sd-0.032470657241012, 32'sd0.030340592258225052, 32'sd0.08346561854222974, 32'sd-0.013138738074123064, 32'sd-0.028598687426229168, 32'sd0.07266507300507069, 32'sd0.0645515937921543, 32'sd4.044586172627258e-118, 32'sd6.453515195096087e-124, 32'sd1.7554769120122877e-121, 32'sd1.8061750563568228e-123, 32'sd-4.692119109984145e-118, 32'sd-1.611247198616541e-119, 32'sd0.09897279228563842, 32'sd0.04178358202521092, 32'sd-0.03547554146888764, 32'sd0.05701192717851152, 32'sd0.09703712692168713, 32'sd0.01384049167651123, 32'sd0.09883363075842572, 32'sd0.006447357663898453, 32'sd0.008738723089072854, 32'sd0.1326195962998386, 32'sd0.19621387011890498, 32'sd0.03923652009015045, 32'sd0.04057593247667155, 32'sd-0.0018084068107459836, 32'sd-0.0003377426413080327, 32'sd-0.017777713614429997, 32'sd0.005817642568338566, 32'sd-0.002401513596154494, 32'sd-0.0019761067430745837, 32'sd0.01849254393684938, 32'sd-5.624503643982012e-122, 32'sd2.2436614841485176e-123, 32'sd8.008641516168802e-125, 32'sd-1.2529198424003644e-125},
        '{32'sd7.628660531308377e-127, 32'sd4.960680105658839e-128, 32'sd1.4210343638778798e-122, 32'sd-1.1966218819229915e-126, 32'sd5.662219930830524e-115, 32'sd-2.991685471774893e-121, 32'sd-1.0378593640878501e-119, 32'sd7.693413343965837e-123, 32'sd5.388180402679606e-123, 32'sd7.10346551880371e-124, 32'sd-1.2595188706377725e-123, 32'sd-2.4561080758535718e-117, 32'sd0.04907619402156039, 32'sd0.08446049366181635, 32'sd-0.07149742220244212, 32'sd0.015031818027502863, 32'sd-1.3750463464553677e-127, 32'sd9.601164520143873e-120, 32'sd-1.8209398705073459e-121, 32'sd4.7324164072774536e-123, 32'sd-1.6570961811937485e-120, 32'sd2.159878587658593e-127, 32'sd-2.5156632413720758e-126, 32'sd-2.599226450763323e-124, 32'sd-1.067218231890792e-119, 32'sd1.0733540891415377e-127, 32'sd3.5546664182060784e-114, 32'sd1.728216931604816e-125, 32'sd8.796017316727051e-123, 32'sd-7.800257484651349e-119, 32'sd-9.223758305721756e-125, 32'sd-6.766224577819895e-124, 32'sd0.01838465934456793, 32'sd0.0523010410873226, 32'sd-0.028767985311728538, 32'sd-0.0911894218701913, 32'sd-0.0633432752151562, 32'sd0.04600313241084234, 32'sd-0.041253667663337566, 32'sd0.014682365864109282, 32'sd0.10447404730446326, 32'sd0.00882602078216173, 32'sd0.061594355475714145, 32'sd-0.0508260253269527, 32'sd-0.05435871673897809, 32'sd0.08048689991946448, 32'sd-0.009454519520576745, 32'sd0.06573945421432108, 32'sd0.05740711586575098, 32'sd0.06001312837196392, 32'sd-0.05087299382768952, 32'sd0.04580273228409086, 32'sd-5.217519631789195e-126, 32'sd3.9672403598254674e-119, 32'sd1.2275719910427e-122, 32'sd-1.290371441184573e-117, 32'sd1.7315229582209985e-123, 32'sd-3.4639670894351926e-122, 32'sd0.08364298188264019, 32'sd0.07018891578191014, 32'sd0.04515676706022089, 32'sd-0.015262649841365676, 32'sd-0.020110302032892848, 32'sd-0.11438607289880708, 32'sd0.02381882339458226, 32'sd-0.037140005517785665, 32'sd-0.037013880753824446, 32'sd-0.016646624634342227, 32'sd0.08997726554890546, 32'sd0.13831532807237473, 32'sd0.042140566987840855, 32'sd0.05996483763772308, 32'sd-0.015153558581773252, 32'sd0.0097992516763059, 32'sd-0.16329531046384763, 32'sd-0.06436306988048504, 32'sd0.004636735289247643, 32'sd0.00020826040368658689, 32'sd-0.0104475918034155, 32'sd0.08434453380745842, 32'sd0.10882526088765239, 32'sd0.06506604248011497, 32'sd-3.9965092541218175e-125, 32'sd6.360986284187427e-126, 32'sd-2.125421546714965e-127, 32'sd7.306630497341004e-121, 32'sd-0.006234925957890461, 32'sd-0.005433771783271981, 32'sd0.03780131067487238, 32'sd-0.07340929342709232, 32'sd-0.02625200936218675, 32'sd0.03475332819090962, 32'sd-0.014274691715753228, 32'sd0.06020273274001538, 32'sd0.04864381791041066, 32'sd0.04131425796337437, 32'sd0.046547486116591735, 32'sd0.024382839359837843, 32'sd0.03415001066099973, 32'sd-0.04490841507980248, 32'sd-0.07090810604780655, 32'sd-0.17030231801042173, 32'sd-0.22181221813628102, 32'sd-0.03086859060532661, 32'sd0.06251185154906813, 32'sd-0.06468183804860385, 32'sd-0.03688665696915873, 32'sd0.09205494461764441, 32'sd-0.035476394575987565, 32'sd0.0884612720637504, 32'sd0.11131175207174543, 32'sd3.508158389028903e-126, 32'sd-8.584547951734565e-117, 32'sd0.043420339269294034, 32'sd-0.0068182750438220115, 32'sd0.0455346156746568, 32'sd-0.012185552077966995, 32'sd-0.036478452577838195, 32'sd-0.09588695982335878, 32'sd0.008070146807580754, 32'sd0.04316380586696859, 32'sd0.10108612873279105, 32'sd0.06009366264390375, 32'sd-0.05042770356491991, 32'sd0.07806866748802506, 32'sd0.09495114639714552, 32'sd-0.012867277726128666, 32'sd-0.04460599447084422, 32'sd-0.04274502018378812, 32'sd-0.011985960285788615, 32'sd-0.005388977583706392, 32'sd0.02887091741180733, 32'sd0.01079051817732676, 32'sd0.06013622684001019, 32'sd0.005940543865394309, 32'sd0.06020660028494873, 32'sd-0.007369545131267882, 32'sd0.02914745101590161, 32'sd-0.06064020938490954, 32'sd-0.04701905915303424, 32'sd-3.5488731458418265e-119, 32'sd0.005396093989985731, 32'sd-0.026352308752737887, 32'sd0.0010015459860730066, 32'sd0.006769182905656233, 32'sd-0.0428718350997916, 32'sd-0.02310299623054755, 32'sd0.07073903157216645, 32'sd0.07631939490337075, 32'sd0.10526025715193364, 32'sd0.09117818642577735, 32'sd-0.05372124834137748, 32'sd-0.044671525715006176, 32'sd-0.14263373967581924, 32'sd0.029208572739351863, 32'sd0.0015994384270099887, 32'sd0.054414112425185186, 32'sd-0.04012183008676294, 32'sd-0.1344204141669844, 32'sd-0.00731215701763739, 32'sd-0.02687143853939089, 32'sd-0.025188176231985774, 32'sd0.06240968669876307, 32'sd0.08282986217473007, 32'sd0.04563864818763962, 32'sd0.08296050389398371, 32'sd-0.028814341680537446, 32'sd0.06236149235031388, 32'sd-1.3642234121490212e-124, 32'sd0.001126736455528817, 32'sd-0.03155267336866635, 32'sd-0.05670762771628989, 32'sd-0.07598780257023685, 32'sd0.08172418566625593, 32'sd0.035550558801641576, 32'sd-0.014899296014458515, 32'sd0.07969811107755412, 32'sd-0.03863256078591552, 32'sd0.012179231433677377, 32'sd-0.08774519441089042, 32'sd-0.16998356001837694, 32'sd-0.1338323565127796, 32'sd-0.07140200605615443, 32'sd0.010552616267404514, 32'sd-0.1818747616170439, 32'sd-0.07315731119072177, 32'sd-0.12135252176725776, 32'sd-0.18016251977055248, 32'sd0.04650294557491419, 32'sd-0.08699174538797755, 32'sd0.108855932503713, 32'sd0.18240812193542402, 32'sd0.1769687443421979, 32'sd0.0784955228710059, 32'sd0.1016748040444111, 32'sd0.036699405901370476, 32'sd0.07563616178591176, 32'sd-0.01744234891644756, 32'sd-0.029199679647523378, 32'sd-0.008419381699986243, 32'sd-0.10991268512170481, 32'sd0.07509707531580138, 32'sd0.03231351706536314, 32'sd0.0799242601128159, 32'sd0.02474435107475657, 32'sd0.06638075754294971, 32'sd0.03180375299003162, 32'sd0.01937124032527781, 32'sd-0.12234256408212695, 32'sd-0.07015663470981033, 32'sd0.02523053413075123, 32'sd-0.025037892092850633, 32'sd-0.15517966935091224, 32'sd0.04968682065541657, 32'sd-0.11489612825824244, 32'sd-0.018939517413761136, 32'sd0.02005747397240631, 32'sd0.08787091082232061, 32'sd-0.03225790328290229, 32'sd-0.03776281873615222, 32'sd0.07709067579914614, 32'sd0.058430625636465255, 32'sd0.023702383657675553, 32'sd-0.006452537872141219, 32'sd0.034749682689941316, 32'sd-0.09353118672998988, 32'sd-0.07939670732366733, 32'sd0.008100082035887832, 32'sd-0.07578416151772448, 32'sd-0.02205968445314373, 32'sd0.018026197825059175, 32'sd0.17195124795839167, 32'sd0.08965474405273248, 32'sd0.1776109675394862, 32'sd-0.040073091726205254, 32'sd-0.07798130557798694, 32'sd0.012991268727102923, 32'sd-0.026104959125125504, 32'sd-0.011152994239403302, 32'sd0.03127061318508834, 32'sd-0.13843280791645665, 32'sd-0.11521429080939688, 32'sd-0.07011072840706452, 32'sd-0.0367320220510887, 32'sd0.11209286046196468, 32'sd0.15563310165574537, 32'sd0.0834870881057765, 32'sd-0.03440781293808268, 32'sd-0.022831541697978124, 32'sd0.01498010287193255, 32'sd0.01151398724954687, 32'sd0.0442121644780211, 32'sd0.001417984248296889, 32'sd-0.005610452671888452, 32'sd-0.02249449419797462, 32'sd-0.10233461741303711, 32'sd-0.023719545644245745, 32'sd-0.04954932700148617, 32'sd-0.08725820448485055, 32'sd0.16926339435487328, 32'sd0.04481168304475361, 32'sd-0.04632599160448844, 32'sd0.007555392721373275, 32'sd-0.05906867306769656, 32'sd-0.1246932312913436, 32'sd-0.09038112394631989, 32'sd-0.10987871712302498, 32'sd0.036292184170224735, 32'sd-0.06810643092434515, 32'sd-0.12475160173182631, 32'sd-0.07246264813462068, 32'sd0.07048288122464452, 32'sd0.15706364501052303, 32'sd0.16492142777603647, 32'sd0.060590432987018626, 32'sd0.042473790267658, 32'sd0.032489559825517295, 32'sd0.02246743801183653, 32'sd0.05859668516696454, 32'sd-0.00874345999571967, 32'sd0.02623782467051993, 32'sd-0.05096723646738895, 32'sd-0.06808952886116973, 32'sd0.04541834907808767, 32'sd-0.04340150820835492, 32'sd-0.2582267513307941, 32'sd0.023794038487143926, 32'sd0.052037331898711146, 32'sd0.12334264337325078, 32'sd0.16671193507193385, 32'sd0.14861112346646702, 32'sd-0.0604916426804375, 32'sd-0.015472740932561364, 32'sd-0.0014378608416661398, 32'sd-0.11913424400387888, 32'sd-0.016302075726867885, 32'sd-0.12027963089288703, 32'sd-0.12337072846715895, 32'sd-0.0115666719661459, 32'sd0.14288465685688753, 32'sd0.07571525913550309, 32'sd-0.004107400130903031, 32'sd0.08254006937994166, 32'sd0.18697304020186142, 32'sd0.06177643164779937, 32'sd-0.06723269215215816, 32'sd-0.05441858356411279, 32'sd-0.06688898563713287, 32'sd0.003217298830387905, 32'sd-0.027839492997741324, 32'sd0.06601585144826838, 32'sd-0.016589485425280496, 32'sd-0.09179596425827288, 32'sd-0.13452715491352268, 32'sd-0.05371081772687943, 32'sd-0.12172086543831542, 32'sd-0.020485491489144424, 32'sd0.11535966347855722, 32'sd0.09115156659816762, 32'sd-0.06858975803537792, 32'sd-0.005843030995217591, 32'sd0.07182159321526435, 32'sd-0.018059091435747167, 32'sd0.025363893404120798, 32'sd0.0010825604050952275, 32'sd-0.12656372399466728, 32'sd-0.12368359459625171, 32'sd0.10279645486126113, 32'sd0.04451197351106709, 32'sd0.15022293322347538, 32'sd0.044992625393408786, 32'sd-0.036167424125030295, 32'sd-0.03217263546387209, 32'sd-0.0848166036557743, 32'sd-0.050186232242672275, 32'sd-0.026759272938226313, 32'sd0.06575115692978101, 32'sd0.043503843071167635, 32'sd0.025894594331987333, 32'sd-0.00746644277043925, 32'sd-0.05222198382230063, 32'sd-0.15241528069008514, 32'sd0.016494036699788082, 32'sd0.10479298854719236, 32'sd0.10288758510615381, 32'sd0.08320914999807087, 32'sd0.0036946018783557875, 32'sd-0.07086062008377692, 32'sd-0.03969002122368726, 32'sd0.1640020454868408, 32'sd0.07515526801556408, 32'sd0.12090637923953904, 32'sd0.026689150262380456, 32'sd-0.07283081466731964, 32'sd0.007228473456277254, 32'sd-0.03925949579759248, 32'sd0.12774604739581244, 32'sd0.002555770171349697, 32'sd0.04165439184661915, 32'sd-0.0008465727762130637, 32'sd0.0465828264436003, 32'sd0.012000829353695714, 32'sd-0.10036766723553281, 32'sd0.07149176870994843, 32'sd0.014939085189622793, 32'sd-0.022283450734128952, 32'sd-0.0006284912621034259, 32'sd-0.12246729161172819, 32'sd-0.11787569529325832, 32'sd-0.11505124578186136, 32'sd0.04932472141033664, 32'sd0.01981634798091799, 32'sd-0.03487394346913426, 32'sd0.07393873409586652, 32'sd0.02575793735936772, 32'sd-0.033635952235520954, 32'sd-0.047929308855648556, 32'sd0.013459608370768079, 32'sd0.07690421138769507, 32'sd0.17456084161408056, 32'sd-0.11024400240419073, 32'sd-0.10278221767065607, 32'sd0.0061907270780120335, 32'sd-0.012298265733253112, 32'sd0.018743474257231215, 32'sd-0.006872638349980586, 32'sd0.046255215250981155, 32'sd0.10631645199934583, 32'sd-0.04266018206080319, 32'sd-0.023426547475061243, 32'sd-0.04508649890386917, 32'sd-0.005156346099030981, 32'sd0.003100587810760375, 32'sd0.01982344906762925, 32'sd0.05325580853902437, 32'sd-0.09061057886178153, 32'sd-0.06023008733990267, 32'sd-0.06220738351319141, 32'sd-0.0961350506899226, 32'sd0.05696234220681583, 32'sd0.005382078338739757, 32'sd-0.04278307793963789, 32'sd-0.1765378148802055, 32'sd-0.15228646939396945, 32'sd-0.0386323536260262, 32'sd0.017795714152444263, 32'sd0.10174067914014649, 32'sd0.15293630575653933, 32'sd0.04378140602708057, 32'sd-0.027607406487473653, 32'sd0.013794388547922082, 32'sd0.06751009008249047, 32'sd-0.1904281527986006, 32'sd-0.12446608529271878, 32'sd0.02888671236685895, 32'sd0.03327928806820995, 32'sd-0.02954723669181942, 32'sd-0.13862969831678898, 32'sd-0.017958735026336436, 32'sd0.007294973155185509, 32'sd-0.07418435969170457, 32'sd0.0322563360544526, 32'sd-0.03418227314972225, 32'sd-0.04271346404386341, 32'sd-0.02972420434650195, 32'sd-0.024158620113930593, 32'sd-0.056907493280956026, 32'sd0.010349903306915565, 32'sd-0.03130695923516379, 32'sd-0.06905945117249375, 32'sd-0.04764335083885911, 32'sd-0.12993701706145405, 32'sd-0.06833371552299766, 32'sd-0.010852666713438786, 32'sd0.07227701530334386, 32'sd0.09986874105379237, 32'sd-0.022414690491224017, 32'sd0.07173051792455698, 32'sd-0.009160180200292212, 32'sd-0.169717259580167, 32'sd-0.0772634610073829, 32'sd-0.16202816756211416, 32'sd0.0409790178848215, 32'sd-0.030522396811845348, 32'sd-0.11962840174006868, 32'sd0.04117253569356812, 32'sd-0.0799475829196195, 32'sd0.018215730875456488, 32'sd0.055906603566389296, 32'sd-0.022458345561402894, 32'sd-0.07054510437974933, 32'sd-0.03466617874284986, 32'sd-0.022305027327193902, 32'sd0.029550912682405485, 32'sd-0.10773846224766906, 32'sd-0.09652292560327434, 32'sd0.005449910884034443, 32'sd-0.046878898791046585, 32'sd-0.1545607745059143, 32'sd0.01473273433193185, 32'sd-0.03328773372074394, 32'sd0.093661022320882, 32'sd-0.03173129781851893, 32'sd-0.03758258250567767, 32'sd0.06805327677783193, 32'sd-0.06632063533858232, 32'sd0.011601633812382101, 32'sd-0.052783852716173404, 32'sd-0.19209375776849383, 32'sd-0.104989600395536, 32'sd-0.03800912111911795, 32'sd0.00041398919509469227, 32'sd0.020432978845238443, 32'sd0.10405724043035518, 32'sd0.02505674162798985, 32'sd0.045087185875931836, 32'sd1.341655886900175e-122, 32'sd-0.0762378744934119, 32'sd0.023534112876419818, 32'sd-0.015551310940748431, 32'sd-0.0012172051712131301, 32'sd-0.00850332462566963, 32'sd0.007426456506393311, 32'sd-0.042662360669088815, 32'sd-0.09814169947892927, 32'sd-0.07732468930273258, 32'sd-0.047096463297142954, 32'sd0.10033465315778044, 32'sd0.16642823192476414, 32'sd0.10157079875242057, 32'sd0.06436284932069262, 32'sd0.048716641625808875, 32'sd0.08961474287566681, 32'sd0.038997357311277736, 32'sd0.04799044199283995, 32'sd0.04268145242607179, 32'sd-0.03316810297897842, 32'sd-0.00884595615491064, 32'sd-0.04580943412458918, 32'sd-0.017386127932703208, 32'sd-0.016168548280791492, 32'sd0.012508871417885627, 32'sd-0.06747830830297684, 32'sd-0.05010363476278994, 32'sd-0.014256571085567526, 32'sd0.07816787661481069, 32'sd-0.03129670209218909, 32'sd-0.002436805153553713, 32'sd-0.04086248657259109, 32'sd-0.03984826352906631, 32'sd-0.0003949867762289301, 32'sd-0.08179701719509591, 32'sd-0.11010691317233043, 32'sd-0.17554357385381295, 32'sd-0.05259035149517808, 32'sd0.05471436009516824, 32'sd0.23164068754972023, 32'sd0.24330932359397517, 32'sd0.08299032160315298, 32'sd0.08988587015684163, 32'sd0.07504547347565119, 32'sd0.027584080129258545, 32'sd0.1207298242221687, 32'sd-0.07898605911611307, 32'sd-0.022102595189918976, 32'sd-0.07447318966116365, 32'sd-0.08774828854202313, 32'sd-0.027976284632633228, 32'sd0.0034962015321337065, 32'sd0.028866318606492174, 32'sd-0.07351755356110547, 32'sd-0.043019621124600047, 32'sd0.08495150722721605, 32'sd-0.06032427372107397, 32'sd-0.028220549059987245, 32'sd0.02527627221493188, 32'sd-0.003997758667441261, 32'sd-0.05302971334147704, 32'sd-0.143025899191992, 32'sd-0.09337921503160647, 32'sd-0.08268629447899621, 32'sd-0.040685534571189876, 32'sd-0.035530770286882264, 32'sd0.14847576414745012, 32'sd0.099597860863798, 32'sd0.10803552674441681, 32'sd0.05553224977656479, 32'sd-0.0031614179885900706, 32'sd0.005719199616394155, 32'sd-0.020130701954305052, 32'sd0.06677596570946562, 32'sd0.00032190047198881914, 32'sd-0.06836513027729159, 32'sd-0.07066046285344112, 32'sd-0.010978993924423133, 32'sd-0.0650886770551591, 32'sd-0.005501269452079921, 32'sd-0.03305708306990783, 32'sd-0.0945819181020831, 32'sd0.059587498016476836, 32'sd-3.0308222623026965e-122, 32'sd-0.08523140604654468, 32'sd0.04729012086538934, 32'sd-0.004232358381225038, 32'sd-0.13792362013546985, 32'sd-0.1386441434989491, 32'sd-0.034147524180047316, 32'sd-0.14617036723799168, 32'sd-0.15348008886983544, 32'sd-0.08330741100998884, 32'sd-0.022848345637135316, 32'sd0.16223259242108234, 32'sd0.18662824711727133, 32'sd0.011793838184246659, 32'sd0.008780971881288195, 32'sd0.08097407606538076, 32'sd0.11203729158821762, 32'sd0.07393188763089721, 32'sd-0.000860562249124359, 32'sd0.027798568486270908, 32'sd0.08510491217522867, 32'sd0.022997930881261338, 32'sd-0.14054566491118436, 32'sd-0.07353610889886636, 32'sd0.05370037171999871, 32'sd0.06035729966979121, 32'sd0.040557004543973894, 32'sd0.028762140452185628, 32'sd0.001226983837528582, 32'sd0.04676226504059297, 32'sd0.00740288483942348, 32'sd0.03209674859669555, 32'sd-0.07800496739175446, 32'sd-0.09442689785045799, 32'sd0.019110913415553484, 32'sd-0.12518692884288293, 32'sd-0.07644219818387199, 32'sd0.01944906576296541, 32'sd0.03686036773620557, 32'sd-0.026390922365948054, 32'sd0.01047134125674201, 32'sd-0.0028653889795000075, 32'sd-0.01501269558308825, 32'sd-0.02209615156515374, 32'sd0.06160835588414335, 32'sd0.03184827772124641, 32'sd-0.025376703597905025, 32'sd-0.009491793544066606, 32'sd-0.061074720384605326, 32'sd0.01938739398185239, 32'sd-0.01341194195435712, 32'sd0.09019952683370971, 32'sd0.013164554511805619, 32'sd-0.0033480294807086038, 32'sd-0.04153520036930218, 32'sd-0.025694017386843425, 32'sd0.07846246995793746, 32'sd0.08853943149374113, 32'sd0.011722520482073166, 32'sd-0.025149980868080336, 32'sd-0.011275943204600148, 32'sd-0.018261641623242595, 32'sd-0.16510494097516423, 32'sd-0.09640754666047545, 32'sd-0.11001097390252423, 32'sd0.09143989207052629, 32'sd0.0043641571671971455, 32'sd0.032258668374762704, 32'sd0.0790089757544039, 32'sd0.0621989576059945, 32'sd0.033602434456121065, 32'sd-0.016428124719941106, 32'sd0.013723249752005838, 32'sd-0.04951077432212547, 32'sd-0.010176798751340864, 32'sd0.050356026214586784, 32'sd-0.006160743152619482, 32'sd-0.027153797435943688, 32'sd-0.019412814404157954, 32'sd0.0033711387327725897, 32'sd-0.030151555893356954, 32'sd0.12140878578490555, 32'sd-0.037710736527939166, 32'sd0.05259890733065791, 32'sd6.565527360722975e-127, 32'sd0.027924112313886147, 32'sd-0.07430072084567921, 32'sd-0.007848267360346706, 32'sd0.0711755169357717, 32'sd-0.003130305056102563, 32'sd-0.1176650440127207, 32'sd-0.15044162691563404, 32'sd0.06870179239565243, 32'sd0.09934936955219369, 32'sd0.059858754759167875, 32'sd-0.017712591874242102, 32'sd0.09077887750435243, 32'sd0.0005184730294839627, 32'sd0.1743349497159667, 32'sd0.027598252361009542, 32'sd0.0627063829466556, 32'sd0.016129207870181093, 32'sd0.012010441846905773, 32'sd0.010833758409752802, 32'sd-0.00951970352441618, 32'sd0.037800993752462146, 32'sd-0.04771028367318856, 32'sd-0.053438718757321174, 32'sd0.03434103549867464, 32'sd0.08180531367699086, 32'sd0.06499292609404381, 32'sd-6.115664412464842e-115, 32'sd-2.1306710854618977e-118, 32'sd1.0591272619168101e-115, 32'sd-0.07508966035124223, 32'sd0.04146427156589811, 32'sd-0.01601953620588124, 32'sd-0.08634615205804737, 32'sd-0.058530790303575136, 32'sd-0.1628495875366739, 32'sd-0.18690482522584875, 32'sd-0.0546799754986786, 32'sd-0.05363674839554477, 32'sd0.12347370147692888, 32'sd0.014927607523840343, 32'sd-0.012611220655099488, 32'sd0.09448480361280497, 32'sd-0.0172873692446767, 32'sd-0.06556173442233224, 32'sd-0.05475818071748885, 32'sd-0.036484415808232994, 32'sd-0.06398707319582261, 32'sd-0.09647162836518107, 32'sd0.05551748229688336, 32'sd0.1560926635195623, 32'sd0.037377908180882484, 32'sd0.025229535042096116, 32'sd0.05089127433747253, 32'sd0.021587269210698284, 32'sd1.528312714084053e-121, 32'sd1.3948499996896505e-126, 32'sd-2.2074071645599558e-117, 32'sd0.05035562688788727, 32'sd0.0625476011992142, 32'sd-0.06764048114007733, 32'sd0.03623736995861305, 32'sd0.007167097815199807, 32'sd-0.04289835272816422, 32'sd-0.12179246905387693, 32'sd-0.07381542580239794, 32'sd-0.09169692707394483, 32'sd-0.06325344751667572, 32'sd-0.15293352008515482, 32'sd-0.027380881461998227, 32'sd-0.03782223853777937, 32'sd-0.010512354990803496, 32'sd-0.03136662164811003, 32'sd-0.08874076352649264, 32'sd0.03126089295361986, 32'sd0.03273453299529466, 32'sd0.08258892152275153, 32'sd0.04067377607452682, 32'sd0.0191625088776075, 32'sd0.012733508937361129, 32'sd-0.10357126742125494, 32'sd0.017409376364913947, 32'sd0.05074369767222036, 32'sd-1.2657372140911153e-115, 32'sd8.039321717667905e-121, 32'sd-6.362690819769381e-127, 32'sd1.3132922695100515e-118, 32'sd0.07032285983237126, 32'sd-0.016232499679734686, 32'sd0.12553415206721427, 32'sd0.10436840018204104, 32'sd0.04576741430878755, 32'sd-0.03646377360953577, 32'sd-0.05039270249942779, 32'sd-0.029764659666366357, 32'sd-0.06313454274108604, 32'sd0.02253655945720238, 32'sd-0.012311760805764339, 32'sd-0.09383811733034425, 32'sd-0.07261449084598344, 32'sd0.07504485079540581, 32'sd-0.00397330666295448, 32'sd-0.02210071037253804, 32'sd-0.0185495777049545, 32'sd-0.003063738003892839, 32'sd-0.020157518451380675, 32'sd0.0180146587403752, 32'sd0.0071250604871331375, 32'sd0.025376756394126898, 32'sd0.010203996886191863, 32'sd-4.460769987078691e-126, 32'sd1.759577517081319e-124, 32'sd4.301353086377586e-127, 32'sd-1.5199137101221743e-123, 32'sd-3.1990586082541884e-118, 32'sd8.111260472211538e-121, 32'sd0.08623772075628773, 32'sd0.027309231485760917, 32'sd0.020978112716522782, 32'sd0.06118607096856462, 32'sd-0.024282014025874633, 32'sd0.016220040451359354, 32'sd-0.03649001824861609, 32'sd0.025302756300631345, 32'sd-0.03880401930157288, 32'sd0.015992583059684568, 32'sd-0.028526160069614115, 32'sd-0.09348006250587118, 32'sd0.005394003781376437, 32'sd0.059146530170209856, 32'sd-0.04334943062166646, 32'sd-0.03883161900231845, 32'sd0.10735488211967222, 32'sd0.009405434424726003, 32'sd0.005956224687431784, 32'sd-0.05886628592770054, 32'sd3.312041738869503e-119, 32'sd4.2930451521641124e-125, 32'sd-3.983989886995441e-129, 32'sd-7.0765575048646605e-115},
        '{32'sd-3.7314123740096515e-123, 32'sd-9.188744563662249e-125, 32'sd-6.901372734312381e-128, 32'sd4.204532235784697e-120, 32'sd-2.869598630745413e-121, 32'sd-1.3833059358374906e-122, 32'sd-1.3991492514615377e-125, 32'sd-1.1208596957162607e-116, 32'sd-8.553868055242315e-122, 32'sd-3.494918614614154e-118, 32'sd-9.90638103297406e-121, 32'sd1.3050767567280127e-117, 32'sd0.03698150352280679, 32'sd-0.041599883118019244, 32'sd-0.00611301277348007, 32'sd-0.03758213547769738, 32'sd-3.979473361989027e-120, 32'sd-1.2287932826811293e-122, 32'sd-3.935005990895465e-123, 32'sd6.277029936685281e-117, 32'sd3.0167461963868357e-119, 32'sd-1.8090661952743953e-114, 32'sd-1.0689963445293562e-126, 32'sd-1.2738326664729396e-122, 32'sd-1.988044287565447e-121, 32'sd-7.661590103327629e-126, 32'sd2.8286137947678087e-121, 32'sd3.4045539287223987e-129, 32'sd3.4747384845215916e-119, 32'sd-1.0298904078788807e-120, 32'sd-3.938957477137292e-121, 32'sd6.478408614608202e-126, 32'sd0.026269472213179042, 32'sd-0.05095789688428745, 32'sd-0.016764652765921352, 32'sd-0.051370089517880455, 32'sd0.0012946664101747497, 32'sd0.009353801640978142, 32'sd0.05909066954488938, 32'sd-0.015697638211861358, 32'sd0.03310681742217545, 32'sd-0.040981277521368854, 32'sd-0.07077513883833883, 32'sd-0.08004763491219455, 32'sd0.04425722510078975, 32'sd0.08891999722837189, 32'sd0.05856459848945926, 32'sd-0.04153817638567568, 32'sd0.022414619065659905, 32'sd-0.07560155551510518, 32'sd0.0055392710404099845, 32'sd-0.01601276863447999, 32'sd2.1242032747245974e-126, 32'sd-3.9688848219932645e-119, 32'sd2.7568110481641068e-120, 32'sd1.1622721156145645e-115, 32'sd-8.921668698845059e-123, 32'sd3.782183729771997e-127, 32'sd-0.01137835402184866, 32'sd-0.040549694130516345, 32'sd0.010128758558999851, 32'sd0.07204255987516225, 32'sd-0.060282785177863334, 32'sd0.05337526980990945, 32'sd0.036780631958415286, 32'sd0.03384807746882166, 32'sd-0.03575937279789293, 32'sd-0.036916257764954837, 32'sd-0.05302633897402498, 32'sd0.012001162979056661, 32'sd-0.06435043463816131, 32'sd0.03012142573871813, 32'sd-0.15142987396297072, 32'sd0.0182060079096746, 32'sd0.08980785791651971, 32'sd-0.03647841416659099, 32'sd-0.002916590579695781, 32'sd-0.048666382160787766, 32'sd0.014326679642113664, 32'sd-0.08632307276205611, 32'sd-0.05045704765159653, 32'sd-0.04544850121748596, 32'sd-5.379327166126752e-124, 32'sd-5.294964589309349e-126, 32'sd-2.57060499257193e-123, 32'sd-1.0282709687056038e-120, 32'sd-0.007406327424506629, 32'sd-0.0632793775396716, 32'sd0.03679004414784448, 32'sd0.019636810540647, 32'sd0.03325627030064576, 32'sd0.050793948435601664, 32'sd0.05435739235817778, 32'sd-0.0026397945558159506, 32'sd-0.11340488692263775, 32'sd-0.024268508089780372, 32'sd0.05927946233789172, 32'sd-0.03886632454374826, 32'sd-0.023212876957073213, 32'sd-0.022956446306003388, 32'sd0.0808462738864542, 32'sd0.019162103038068777, 32'sd0.06734267265092622, 32'sd-0.11491684426382365, 32'sd-0.04043050451430033, 32'sd0.04046350181111813, 32'sd-0.018120328975876742, 32'sd0.04003652637072256, 32'sd0.02880249073933215, 32'sd-0.00861738179580492, 32'sd0.043802306535221415, 32'sd2.3505547844639063e-129, 32'sd-6.9265593790721116e-124, 32'sd0.04708910036730388, 32'sd-0.04469154458697255, 32'sd0.0247762892266328, 32'sd0.09458974733060399, 32'sd-0.02495875976362696, 32'sd-0.016482671897540165, 32'sd-0.08923094190593081, 32'sd-0.08122705216025784, 32'sd-0.18087972175028363, 32'sd-0.2296997581890913, 32'sd-0.015009079266594769, 32'sd0.08782595636208297, 32'sd0.04633327552541073, 32'sd0.05487070264118497, 32'sd0.04156793574950336, 32'sd-0.017576499312603622, 32'sd-0.0005458692426505569, 32'sd0.02281030497430041, 32'sd-0.008977744748259278, 32'sd0.025314844585586364, 32'sd0.14775467957990676, 32'sd0.0014557511350214171, 32'sd0.11100350202099829, 32'sd0.08158480745680811, 32'sd0.10904247364560153, 32'sd-0.056996208073483844, 32'sd0.012336532380284137, 32'sd-2.4218882439393344e-124, 32'sd-0.054914155948490924, 32'sd-0.002291504597776693, 32'sd0.04867271470048383, 32'sd0.012637006746763234, 32'sd-0.09989434260621159, 32'sd-0.055642071555207735, 32'sd-0.00836654584838422, 32'sd-0.12256949323448639, 32'sd-0.07235403452483573, 32'sd0.039472579173669836, 32'sd0.10443428746770037, 32'sd0.12999373823513935, 32'sd0.09829718992854941, 32'sd0.10697364791579449, 32'sd0.06422214232135823, 32'sd0.06596137684990308, 32'sd0.03415499969097053, 32'sd0.007268814568969851, 32'sd0.03558874614143251, 32'sd0.013079155052007607, 32'sd-0.0211732306700193, 32'sd0.01607418781748044, 32'sd0.0176312371603579, 32'sd0.018326698858135634, 32'sd0.011107274611154445, 32'sd-0.008002671033365001, 32'sd-0.052976969366121236, 32'sd9.189868272275318e-120, 32'sd-0.03930823505955734, 32'sd-0.08075084947314334, 32'sd-0.04960632228204131, 32'sd-0.022350208351957383, 32'sd-0.06096595297199075, 32'sd-0.11793044574760178, 32'sd-0.06687220564018306, 32'sd0.029302122370191398, 32'sd-0.11486135024527798, 32'sd0.05419556939826027, 32'sd0.06650266101842489, 32'sd-0.004161526716032232, 32'sd0.06996719835414462, 32'sd0.021782859643146624, 32'sd-0.057458258030661, 32'sd-0.02129586752542347, 32'sd-0.010797305514170137, 32'sd-0.0821675852831761, 32'sd-0.06638118644809088, 32'sd-0.06013505505643067, 32'sd-0.0537726375541305, 32'sd0.15813358562842267, 32'sd0.18897316426435176, 32'sd0.05864080476041745, 32'sd-0.16919793427637525, 32'sd-0.08696922609852063, 32'sd0.009832399288299638, 32'sd0.0007683033245202658, 32'sd0.026841161571232855, 32'sd-0.09949557920595216, 32'sd-0.02500471056159853, 32'sd-0.048622962802928146, 32'sd0.06156235501466602, 32'sd0.0027675068623676815, 32'sd-0.13363323821007808, 32'sd0.029002075707463455, 32'sd0.037097598650638504, 32'sd-0.030172622676317793, 32'sd0.060872487825971544, 32'sd0.0012988864091804193, 32'sd-0.024770210775792893, 32'sd-0.03611364214192085, 32'sd0.020151982739523004, 32'sd0.07524960365670975, 32'sd-0.013402151063776147, 32'sd0.026490594532115472, 32'sd-0.03573743188271689, 32'sd-0.0368818538628965, 32'sd-0.06460145004579433, 32'sd-0.07540924734719072, 32'sd-0.011135811717000631, 32'sd-0.003372984255677864, 32'sd-0.11234259344784221, 32'sd-0.0739712684562183, 32'sd-0.02418915306231386, 32'sd0.05295475154840487, 32'sd-0.012785627368724458, 32'sd0.06997755713070668, 32'sd-0.043307195906001086, 32'sd-0.03879928198734982, 32'sd0.020633133328952027, 32'sd-0.07080981598999776, 32'sd-0.015282330847890624, 32'sd-0.03306221068289843, 32'sd-0.05007158966836866, 32'sd-0.062000123636664156, 32'sd-0.008522267965300796, 32'sd0.011273317698861661, 32'sd0.0849847304246035, 32'sd-0.07397871741412865, 32'sd-0.0777963628873314, 32'sd0.005255177367886573, 32'sd-0.06089044196866599, 32'sd0.03317360204472336, 32'sd-0.07942146648261286, 32'sd0.06196808288727275, 32'sd0.023442711646165734, 32'sd0.007881265145553174, 32'sd-0.0446690251902064, 32'sd0.01532377138241737, 32'sd-0.04941442039049588, 32'sd-0.04420258337826459, 32'sd0.056289962252818695, 32'sd0.02227294203300099, 32'sd0.043916136063539085, 32'sd-0.053255322790156656, 32'sd-0.043106699870766416, 32'sd-0.12243625389653913, 32'sd-0.04528143773428746, 32'sd-0.16936407455750682, 32'sd-0.033367709482558634, 32'sd-0.04075893053030629, 32'sd-0.05614948219920111, 32'sd-0.005583354624310888, 32'sd0.0047449941581469935, 32'sd0.011901348215520125, 32'sd0.09378305681735614, 32'sd-0.08327291396051266, 32'sd-0.12683918982757686, 32'sd-0.15436514131935383, 32'sd0.012899698693692644, 32'sd0.10170584523616323, 32'sd0.07604803631009491, 32'sd-0.015158916895595254, 32'sd0.09387477263104721, 32'sd0.033078875424698215, 32'sd0.041158049652353694, 32'sd0.12314534834571389, 32'sd0.14331973649449853, 32'sd0.10034624504923315, 32'sd0.03006892409812426, 32'sd-0.05815857661404843, 32'sd0.011477927449140526, 32'sd-0.029632371237142158, 32'sd-0.021176357033053716, 32'sd-0.15910629974997284, 32'sd-0.10641746461459893, 32'sd-0.04238743312969185, 32'sd-0.12484239496074324, 32'sd-0.1523914097093321, 32'sd-0.04330057062711451, 32'sd0.021956220967732785, 32'sd0.10405478604293433, 32'sd0.16801694642747256, 32'sd0.09539993062038622, 32'sd0.0029715547820489776, 32'sd-0.13543788678467975, 32'sd-0.05842982347641956, 32'sd0.006122449425570022, 32'sd0.13035162594064992, 32'sd0.022573648406649282, 32'sd-0.07472533236864312, 32'sd0.06487187177115102, 32'sd0.10246421514409909, 32'sd-0.019720033457074182, 32'sd0.013032516136656114, 32'sd-0.017656505486511098, 32'sd0.0630459432471093, 32'sd0.03431948063572676, 32'sd0.03623249467899511, 32'sd-0.03542757730570834, 32'sd-0.06452289283586683, 32'sd0.04997822092646257, 32'sd-0.09726313360088579, 32'sd-0.03557335204812431, 32'sd-0.08781178106284074, 32'sd-0.08430243230457267, 32'sd-0.08744550005745892, 32'sd-0.011349191893210214, 32'sd0.06840797377578234, 32'sd0.061333905608201185, 32'sd-0.009782126860557037, 32'sd0.02661998868779684, 32'sd0.09973899629394516, 32'sd-0.02915490785832814, 32'sd0.10162263519119569, 32'sd0.19168455314345223, 32'sd0.17254195197010128, 32'sd0.038945835368994215, 32'sd-0.04618421528759972, 32'sd0.014204274573778625, 32'sd0.006725670277447634, 32'sd0.13141007771412921, 32'sd0.13782699017811834, 32'sd-0.029838889347139873, 32'sd-0.08048486344587057, 32'sd-0.014536023272213271, 32'sd-0.013925871637672066, 32'sd-0.01618030571450766, 32'sd-0.06536441189734274, 32'sd0.017924114085621806, 32'sd-0.02401976644564756, 32'sd0.09509728258535084, 32'sd0.003289787098640378, 32'sd-0.021688607935099517, 32'sd0.0020549630727540536, 32'sd0.043480182172575266, 32'sd-0.087517001391746, 32'sd-0.04321999594627309, 32'sd0.020724398137538028, 32'sd0.10776741410282188, 32'sd0.13893158083032742, 32'sd0.06315400728079072, 32'sd0.05448214077297819, 32'sd0.012910967834816886, 32'sd0.0350870460598102, 32'sd0.08967922315930768, 32'sd0.07717486036743652, 32'sd0.04382406135617138, 32'sd0.038112177349602046, 32'sd-0.002238664119716543, 32'sd0.03910080186375968, 32'sd-0.15894094198903602, 32'sd-0.06892246315763606, 32'sd-0.08522010523323008, 32'sd-0.025382663069033626, 32'sd-0.03154267160627053, 32'sd0.06521602436669505, 32'sd-0.04875208699800856, 32'sd0.09554516126768212, 32'sd0.037278459708941815, 32'sd-0.04126808607358683, 32'sd-0.06131473727559422, 32'sd-0.11289458355892973, 32'sd-0.06577531422629253, 32'sd-0.08130516519303625, 32'sd-0.015819869907934977, 32'sd0.08826816852088643, 32'sd0.14424447829405138, 32'sd0.1771028328267676, 32'sd0.027485153833057663, 32'sd-0.05529406319725737, 32'sd-0.022594873397783016, 32'sd0.028372842625283504, 32'sd0.08213921011488462, 32'sd-0.030486645860074782, 32'sd0.003986618251527829, 32'sd0.001735494977647525, 32'sd0.0459911869604292, 32'sd0.09752387463246974, 32'sd-0.03297684517174448, 32'sd0.048305111841223235, 32'sd0.00368561430012084, 32'sd-0.0029890410489131765, 32'sd-0.05203626883215955, 32'sd-0.016155485507518892, 32'sd0.10198371200411567, 32'sd-0.013842036458928867, 32'sd-0.039010802728484464, 32'sd-0.13329642629264732, 32'sd-0.14365891615501525, 32'sd-0.09886912842198911, 32'sd-0.15075483112089724, 32'sd0.00011202331271551225, 32'sd0.0022766236094042365, 32'sd0.06200850004345582, 32'sd0.14234950924500053, 32'sd-0.034316599666572446, 32'sd0.008538827610942951, 32'sd0.04070894276425516, 32'sd0.016154866837408476, 32'sd0.0681603262979347, 32'sd0.029048381306882576, 32'sd0.015130076245389444, 32'sd-0.01341413002998378, 32'sd-0.06764692451708362, 32'sd-0.10736680402689056, 32'sd-0.030781844625814795, 32'sd-0.06205411146708145, 32'sd0.03856888323222143, 32'sd0.008662620129230839, 32'sd-0.03445617244524263, 32'sd-0.04169645326180168, 32'sd0.05583486053024611, 32'sd-0.0052259933719302895, 32'sd0.005415278184579429, 32'sd-0.03486158235095136, 32'sd-0.0028863058058482853, 32'sd-0.06418338802648314, 32'sd-0.05577793635085172, 32'sd-0.06255335113387438, 32'sd0.02150146648224839, 32'sd-0.028279444431116556, 32'sd0.06154590918210219, 32'sd-0.04350857942818201, 32'sd-0.020750628468648547, 32'sd0.11015843699628837, 32'sd0.02864266924307406, 32'sd0.08078665773060222, 32'sd0.08821352727191639, 32'sd-0.012090774757526014, 32'sd0.013129392244770237, 32'sd-0.1325095553968763, 32'sd-0.11091230405954206, 32'sd-0.12237345068793533, 32'sd-0.1006123459818311, 32'sd-0.0440963135747701, 32'sd-0.064805372425943, 32'sd0.0174881695583065, 32'sd-0.029136625044125578, 32'sd-0.02643163244680949, 32'sd0.017477840502649857, 32'sd0.03765110628592766, 32'sd0.09663852434509689, 32'sd0.09031630421615641, 32'sd-0.0831063776360822, 32'sd-0.06355559464342794, 32'sd-0.04005679592738134, 32'sd-0.18696556254830082, 32'sd-0.14308829944976675, 32'sd-0.1395248082239043, 32'sd0.058795167941514535, 32'sd-0.09281315384300848, 32'sd0.02973910583727506, 32'sd-0.04312839844155437, 32'sd-0.011175626191666746, 32'sd0.1211948842292665, 32'sd0.0601190762649387, 32'sd0.012135849827632862, 32'sd-0.0662925813610042, 32'sd-0.1834126989259581, 32'sd-0.013446784238090221, 32'sd-0.07544130387728577, 32'sd-0.08002579865851313, 32'sd0.03132543548381938, 32'sd-0.015337040127177818, 32'sd-0.005898079368684539, 32'sd1.1667534350671642e-121, 32'sd-0.04919887219116013, 32'sd-0.028645564697324655, 32'sd0.01628399675085312, 32'sd0.008477415356890236, 32'sd-0.01234435659802736, 32'sd-0.014874139606188025, 32'sd-0.1675781442425755, 32'sd-0.18191778294214067, 32'sd-0.1791935308645611, 32'sd-0.2615834124856426, 32'sd-0.11421172193952249, 32'sd0.11361265459364167, 32'sd0.023719417293659745, 32'sd-0.11449524566666788, 32'sd0.013697570147065534, 32'sd0.051395123070758, 32'sd0.16365624459964384, 32'sd0.10156466693975134, 32'sd0.05874636590158745, 32'sd0.020551831257311436, 32'sd0.03523751866142835, 32'sd-0.1464665788804643, 32'sd-0.04621150922435755, 32'sd-0.12935479516228932, 32'sd0.05617794058688836, 32'sd-0.07719746015489057, 32'sd-0.06660917848013889, 32'sd0.024323171604325088, 32'sd-0.058089216145487996, 32'sd0.04491776310174501, 32'sd-0.07405588041274751, 32'sd0.13422939254920221, 32'sd0.06563519260480923, 32'sd0.062942362730818, 32'sd-0.016251177212757345, 32'sd-0.00849640386392118, 32'sd-0.03018787554118946, 32'sd0.010982698233448603, 32'sd0.08518098625526797, 32'sd0.0944634020622673, 32'sd-0.02180237501733948, 32'sd-0.1285352544475443, 32'sd-0.05003294048402363, 32'sd0.023724515361964262, 32'sd0.14747863248601617, 32'sd0.11088535618700593, 32'sd-0.039472519188885384, 32'sd0.0021948879332387137, 32'sd-0.12334837567229585, 32'sd-0.043694867083692294, 32'sd-0.09163355192750697, 32'sd0.007527982912008539, 32'sd-0.04811456009102431, 32'sd0.08037170606776992, 32'sd-0.08443395622085068, 32'sd0.004603671435681623, 32'sd-0.039911712986083724, 32'sd-0.03952710101931767, 32'sd0.04268815563782531, 32'sd0.04060445547518533, 32'sd0.024689263065537537, 32'sd0.09486733337792193, 32'sd-0.016189010271537477, 32'sd0.005424506757652609, 32'sd0.01994710691678245, 32'sd0.0021475658695756846, 32'sd-0.017758782207561587, 32'sd-0.08399083983048869, 32'sd-0.068848570391386, 32'sd-0.059981532628061524, 32'sd-0.05706283685503894, 32'sd0.005631068306207087, 32'sd0.09294140676908637, 32'sd0.13497394330978435, 32'sd-0.06321590684232962, 32'sd-0.0355015078894839, 32'sd-0.06695623799130752, 32'sd-0.1782033116332877, 32'sd-0.07504540634772697, 32'sd0.009597053733691865, 32'sd-0.0005079250973415991, 32'sd0.05991108671331239, 32'sd-0.019071015388498945, 32'sd-3.147878441149586e-119, 32'sd-0.05063498695024514, 32'sd-0.08036381162548088, 32'sd-0.05940899672561483, 32'sd-0.01862150788280709, 32'sd0.13824050110673006, 32'sd0.038305654286201966, 32'sd-0.007378041432217201, 32'sd-0.02156131202453502, 32'sd0.008341090127477751, 32'sd0.04479158263047844, 32'sd0.02111274550037564, 32'sd-0.023599216149228806, 32'sd0.023941725440384518, 32'sd-0.04410285638607148, 32'sd0.023628211196034758, 32'sd-0.005809283962473013, 32'sd0.13515075744535893, 32'sd-0.0038705969183100335, 32'sd-0.05599938979469977, 32'sd-0.22036702040940476, 32'sd-0.08495727824032505, 32'sd-0.13221648275623452, 32'sd-0.02921129008144382, 32'sd0.03505117105277342, 32'sd-0.026628793029344736, 32'sd-0.08069325607849644, 32'sd-0.004975829654576601, 32'sd-0.0006979601803021908, 32'sd-0.05548838338921164, 32'sd0.08272867616813707, 32'sd0.06628924026024145, 32'sd0.0420047248394877, 32'sd-0.06177653718259574, 32'sd-0.009675018946943812, 32'sd-0.05909500681257263, 32'sd-0.08968843628801677, 32'sd-0.04022969392219249, 32'sd0.0938258545152435, 32'sd0.10198868560397982, 32'sd-0.09331237969468915, 32'sd0.013066267879997743, 32'sd0.0839288491289848, 32'sd0.06939358327655333, 32'sd0.05599057912950219, 32'sd0.06692974352893875, 32'sd-0.031303526002591744, 32'sd-0.1597923292068891, 32'sd-0.1651078104549543, 32'sd-0.1167493537155704, 32'sd-0.2086272624184024, 32'sd-0.0793996649845482, 32'sd-0.10911196986209278, 32'sd0.004640085432271319, 32'sd0.004684455623117289, 32'sd-0.009554684755939638, 32'sd-0.010966372838878762, 32'sd-0.025072575111701054, 32'sd0.05573549634124358, 32'sd-0.03034934635742016, 32'sd0.01661133527949169, 32'sd-0.08707679578343985, 32'sd-0.04730400285085508, 32'sd0.08370894734531244, 32'sd0.006393520911963659, 32'sd0.02872292939124917, 32'sd-0.02255440938358913, 32'sd0.010401321791782275, 32'sd0.12580275572720737, 32'sd0.006836055244287957, 32'sd0.07367374184058718, 32'sd0.10273520598895669, 32'sd-0.031308366792240076, 32'sd-0.028856544818668027, 32'sd-0.08567597927128318, 32'sd-0.15684577796872012, 32'sd-0.11339655701408427, 32'sd-0.23708499502942784, 32'sd-0.09589850263986252, 32'sd-0.003368028980017624, 32'sd-0.03478880882074178, 32'sd-0.004048559017404966, 32'sd0.05999959170804036, 32'sd0.01522404183904276, 32'sd2.839656122797966e-116, 32'sd-0.020842240592025656, 32'sd-0.032145814030438924, 32'sd-0.014749586061832673, 32'sd0.043173465110023235, 32'sd0.02357791110196257, 32'sd-0.08320821700824582, 32'sd0.07050964920209575, 32'sd-0.03186775014350777, 32'sd0.017504301715768725, 32'sd0.02925114487295713, 32'sd0.0835289835724211, 32'sd0.06886108065710263, 32'sd0.025785582796110783, 32'sd0.08024951006028284, 32'sd-0.010249273075948924, 32'sd-0.05996041606567983, 32'sd-0.07285471405187774, 32'sd-0.05495756475062344, 32'sd-0.12920845856073926, 32'sd-0.03141932487514055, 32'sd-0.13707108273088925, 32'sd-0.048798921707636195, 32'sd-0.05546312454988511, 32'sd-0.033547123847923126, 32'sd0.0354803226337507, 32'sd-0.11191485352445278, 32'sd2.338189175929349e-122, 32'sd-1.274796001357001e-125, 32'sd3.372121774776245e-115, 32'sd0.004566152714825932, 32'sd0.10289567540384226, 32'sd-0.047486299890403434, 32'sd-0.13196094972034986, 32'sd-0.11014249914837025, 32'sd0.07438871137815982, 32'sd-0.0811935222727719, 32'sd-0.0867269892360328, 32'sd0.05256712107213727, 32'sd0.06336098653407048, 32'sd0.037284863511086015, 32'sd0.15010996223790113, 32'sd0.10966344342637442, 32'sd0.10062732192293578, 32'sd-0.05818848899510239, 32'sd-0.12233560035981367, 32'sd-0.20136526469337102, 32'sd-0.1870057869558165, 32'sd0.05674442604877064, 32'sd-0.0847662645309651, 32'sd-0.059036964744654606, 32'sd0.02114789436136185, 32'sd-0.0022474577717312904, 32'sd0.03820690786014069, 32'sd-0.052254321074132415, 32'sd-5.262542381441759e-116, 32'sd7.1778810570497e-121, 32'sd1.0003775833522613e-120, 32'sd-0.054530532387696104, 32'sd0.04664852752454642, 32'sd-0.06807867235775836, 32'sd-0.0833327848182814, 32'sd0.00342149808441367, 32'sd0.03375226359863163, 32'sd-0.07204968419764785, 32'sd0.06152890929150518, 32'sd-0.002157404351732162, 32'sd0.024065709803548118, 32'sd-0.055538613532653006, 32'sd0.06278962105570915, 32'sd0.02728370258536067, 32'sd0.11182231634477742, 32'sd-0.06013741455922834, 32'sd-0.16721474297000882, 32'sd-0.11482462377150904, 32'sd0.005015179549399037, 32'sd-0.03397059474658844, 32'sd-0.03277916675716374, 32'sd-0.023896000801140474, 32'sd-0.042180577295259224, 32'sd-0.04514841039886466, 32'sd0.01939486244891993, 32'sd0.08040367993799674, 32'sd-1.2487741088403254e-115, 32'sd3.339983869528033e-126, 32'sd2.1637600944426232e-127, 32'sd2.0853868106532735e-127, 32'sd-0.04213233963291629, 32'sd0.08384387459830663, 32'sd-0.010115790316460893, 32'sd-0.06337591088912711, 32'sd0.03786229678595267, 32'sd0.05249983572581087, 32'sd0.01417810374463085, 32'sd-0.09138821276343856, 32'sd0.004432776898953815, 32'sd-0.00659415436310836, 32'sd-0.07686878342799587, 32'sd-0.20660357967823437, 32'sd-0.059890959240123276, 32'sd0.000269725172342997, 32'sd-0.04473837529211354, 32'sd-0.017070534035499883, 32'sd-0.06189478877098625, 32'sd-0.05080705687098439, 32'sd-0.010700549725936542, 32'sd0.013933312683962655, 32'sd-0.0638776966514992, 32'sd-0.03987578956029812, 32'sd-0.0371357878888308, 32'sd9.542974117378244e-118, 32'sd-7.422776964800723e-122, 32'sd4.2812093556753564e-123, 32'sd-1.0286654435213316e-124, 32'sd4.1894729904963544e-125, 32'sd-3.0893589082489846e-127, 32'sd-0.0042712576945085415, 32'sd0.008398405310750106, 32'sd0.026962975238035546, 32'sd0.08214230072010408, 32'sd0.027188572279376187, 32'sd0.048489841014236715, 32'sd-0.02795445013085787, 32'sd-0.08102706801131798, 32'sd0.02577419958573807, 32'sd-0.1112806259412827, 32'sd0.04344655611498909, 32'sd-0.042066709307541916, 32'sd-0.08831975031957325, 32'sd0.004774486694366515, 32'sd0.04414269513680048, 32'sd-0.0030834554900001647, 32'sd-0.041826316468522126, 32'sd-0.04158773297688703, 32'sd0.039865717128322924, 32'sd0.024493090988456326, 32'sd8.284223457150542e-121, 32'sd5.003393454686576e-118, 32'sd2.861757082368279e-125, 32'sd-5.812868209271986e-116},
        '{32'sd3.8665452930064655e-123, 32'sd-1.3411893181403304e-119, 32'sd2.183267230219434e-121, 32'sd6.865555725711905e-125, 32'sd1.3525158280729988e-123, 32'sd-1.0623539669123623e-115, 32'sd2.0360759953223678e-117, 32'sd1.7371613797608063e-125, 32'sd4.2679789515047804e-125, 32'sd-3.6075176294311636e-117, 32'sd4.035052313719559e-117, 32'sd-3.8285627367262076e-117, 32'sd-0.015542791906511321, 32'sd0.09973378798513897, 32'sd0.07986244097251184, 32'sd0.03764249595346556, 32'sd-8.888962163976494e-127, 32'sd1.3273100829531234e-122, 32'sd-1.6121076386490225e-115, 32'sd-8.202887450840994e-119, 32'sd-4.6512084747889314e-129, 32'sd-7.769715642553756e-124, 32'sd-3.480410721713243e-119, 32'sd3.483244771327966e-127, 32'sd1.2082477776518081e-122, 32'sd3.3571958989640012e-121, 32'sd1.4723931480947387e-123, 32'sd-1.1684601433923545e-125, 32'sd-1.039220000898846e-120, 32'sd2.5013224068268752e-120, 32'sd-2.7330914368406857e-121, 32'sd-9.79722498432096e-117, 32'sd-0.041639730640038446, 32'sd0.08932977478046518, 32'sd0.005207965791741842, 32'sd0.02820879678485272, 32'sd0.12192086191699573, 32'sd-0.0034509039574701413, 32'sd0.03426203286379026, 32'sd-0.016673166596607954, 32'sd0.049823520069477316, 32'sd0.016637898418555813, 32'sd0.041308593022580435, 32'sd0.08735673460814225, 32'sd0.1048271854183185, 32'sd-0.07046957309635554, 32'sd-0.10364436500192736, 32'sd0.06872199429523844, 32'sd0.05386561429200641, 32'sd-0.033218855720049, 32'sd0.045335911939389135, 32'sd0.052019944298259096, 32'sd-2.4907620792826936e-126, 32'sd4.789616095896862e-115, 32'sd4.508376407071581e-123, 32'sd-3.8270466479596804e-118, 32'sd1.1547715136808042e-118, 32'sd-2.5191497815903816e-126, 32'sd0.01978782326181951, 32'sd0.03771961061631386, 32'sd0.04721754921871241, 32'sd-0.052743643285260294, 32'sd0.09302512243588326, 32'sd0.0998118723181109, 32'sd0.04878594113815737, 32'sd0.024612432199604403, 32'sd0.018502984117847034, 32'sd-0.10012816646007042, 32'sd-0.10374694083741734, 32'sd-0.0050216559219164025, 32'sd0.011090388236963174, 32'sd-0.06036098856193729, 32'sd0.09596495327247354, 32'sd0.020841810519165282, 32'sd0.042060024460063676, 32'sd0.0025986700777522066, 32'sd0.11726120295315522, 32'sd0.0433477414228978, 32'sd-0.04803884159868431, 32'sd-0.008213678998985055, 32'sd0.04932618785313785, 32'sd0.06331029111396932, 32'sd2.098072397915581e-117, 32'sd-7.857432936497212e-124, 32'sd-2.4003332416273904e-124, 32'sd1.4677429118104862e-125, 32'sd0.08535018901275343, 32'sd0.05745866940754711, 32'sd0.006015486218652374, 32'sd-0.03542759452736239, 32'sd-0.012087105020090397, 32'sd-0.061643010395651, 32'sd-0.044106674921774586, 32'sd-0.07284675484649736, 32'sd-0.056560346625640925, 32'sd-0.14266481048768015, 32'sd-0.16841313091266036, 32'sd0.03821208346202248, 32'sd-0.10106188504410311, 32'sd-0.11251265775683816, 32'sd-0.030591406446310945, 32'sd-0.036794600527225295, 32'sd-0.11507110732450108, 32'sd-0.07742643107628908, 32'sd0.05574488104377449, 32'sd0.12224209343058395, 32'sd-0.07044846996338348, 32'sd-0.03399616113426548, 32'sd0.029030806125165773, 32'sd0.05265069502197511, 32'sd-0.024313227452849098, 32'sd-8.918634129005407e-116, 32'sd9.95370589804402e-121, 32'sd0.028362962197632766, 32'sd-0.008806041577203109, 32'sd0.0676964942545493, 32'sd-0.08857246147944925, 32'sd-0.10936043646133421, 32'sd-0.04209775544627562, 32'sd0.009255363404615346, 32'sd-0.03973369767097779, 32'sd-0.0808393937151682, 32'sd-0.0723952143383291, 32'sd-0.05271467836883442, 32'sd-0.002881170426606948, 32'sd0.02934380407755696, 32'sd0.06832353651006218, 32'sd0.08007714045317688, 32'sd-0.01919446065755436, 32'sd0.08947044893835378, 32'sd0.03386157045098266, 32'sd-0.15593257405650351, 32'sd-0.015467593947263741, 32'sd-0.01677464940953956, 32'sd-0.04533281086132529, 32'sd-0.03840382429865339, 32'sd-0.058223301817864975, 32'sd0.005260341865618534, 32'sd-0.047238157489045106, 32'sd0.017066546361401824, 32'sd2.9988306091239024e-121, 32'sd0.039976456025518504, 32'sd0.05265515059544334, 32'sd0.011675065578525755, 32'sd-0.07057799042332684, 32'sd-0.06415922186494345, 32'sd-0.04723303902241597, 32'sd-0.013453738785768244, 32'sd-0.003613487134782273, 32'sd-0.028790525033060062, 32'sd0.08471198526448435, 32'sd-0.07542569013148512, 32'sd-0.04989578956800672, 32'sd0.09520935256060288, 32'sd0.00779163649920679, 32'sd-0.09503810039177668, 32'sd0.06394741798900229, 32'sd0.007545743701223513, 32'sd-0.09933321059195384, 32'sd-0.04578934547276171, 32'sd-0.04838018226637003, 32'sd-0.049727440382950135, 32'sd-0.10710106017424462, 32'sd-0.08293393173434445, 32'sd-0.06612640250100685, 32'sd-0.015605994494111122, 32'sd0.09394923511420257, 32'sd-0.021959974316891902, 32'sd-2.2354884410032403e-120, 32'sd-0.025926234399252592, 32'sd0.024060831626054307, 32'sd-0.011409369424503915, 32'sd0.055087069707379595, 32'sd0.07834797773422968, 32'sd-0.056978734823860004, 32'sd-0.024259995947398468, 32'sd0.00016935096964452862, 32'sd0.11649269727823877, 32'sd-0.07184950233239755, 32'sd-0.047182558709826496, 32'sd0.051500796489923666, 32'sd0.1595895705908408, 32'sd0.0445448236674525, 32'sd0.06648562328827338, 32'sd0.015626154654827404, 32'sd0.07994113016706964, 32'sd0.10928247692208776, 32'sd-0.037268947375528994, 32'sd-0.03448942318728408, 32'sd0.03959040977096572, 32'sd-0.14055102910321532, 32'sd-0.11610451375899587, 32'sd-0.17683939369764895, 32'sd-0.10530622311140424, 32'sd-0.08322191577886286, 32'sd-0.002102801904117373, 32'sd-0.0023918204931104837, 32'sd0.02106853619236696, 32'sd-0.03441079230278235, 32'sd0.011672987780841916, 32'sd0.009967875238238102, 32'sd0.00847981261211249, 32'sd0.04986645039007227, 32'sd0.017777557956504222, 32'sd0.05992946082521828, 32'sd0.034712233862372065, 32'sd-0.04577223389560276, 32'sd0.008132869039501249, 32'sd-0.03392335659816493, 32'sd0.0469622577382673, 32'sd0.0803760307263558, 32'sd0.1600538049824023, 32'sd0.044869912547441465, 32'sd0.037710161449181774, 32'sd0.09949772769019462, 32'sd0.014052685773124742, 32'sd-0.09152139218003352, 32'sd-0.017378859443018594, 32'sd-0.0783497604437949, 32'sd-0.10729397325933795, 32'sd-0.044560708494560494, 32'sd0.05120144895138769, 32'sd-0.04229749794511294, 32'sd-0.017744356650118462, 32'sd0.007016524590277876, 32'sd-0.018108462171412428, 32'sd0.03488684091682226, 32'sd0.0038924332006603918, 32'sd0.03183157523196472, 32'sd-0.021939777632603633, 32'sd0.0373838979082132, 32'sd0.03448712025757594, 32'sd0.0727308154708586, 32'sd0.11368095427499388, 32'sd0.13471304503083784, 32'sd-0.008639704660645018, 32'sd0.06673910042984767, 32'sd0.02223152869486537, 32'sd0.07725319217535762, 32'sd0.12723121334628099, 32'sd-0.011923951681745586, 32'sd-0.08789705073735021, 32'sd0.1241726856014276, 32'sd0.16742721135350702, 32'sd0.08938994350576954, 32'sd0.02069891613906729, 32'sd-0.06108450628301641, 32'sd-0.13721205290395103, 32'sd-0.025590942412951647, 32'sd-0.061906377242199155, 32'sd-0.0025500231662038244, 32'sd-0.02851238247162281, 32'sd0.07544688366844592, 32'sd-0.0014356789470212827, 32'sd0.028424248247837132, 32'sd0.0064471971705251365, 32'sd-0.02190486086137032, 32'sd0.05631974246396157, 32'sd-0.009037163648358802, 32'sd0.11298956239299526, 32'sd0.0398378356817066, 32'sd-0.06619177185968808, 32'sd0.11395344643579444, 32'sd0.10773110611030715, 32'sd-0.009926950420331666, 32'sd-0.07935844704700784, 32'sd-0.024336897920579775, 32'sd-0.08468542339149543, 32'sd-0.04807206996111526, 32'sd0.0707219833050669, 32'sd-0.026940946336664835, 32'sd0.15040963970007637, 32'sd0.07785689739231516, 32'sd-0.08859983758943464, 32'sd-0.05615243929071112, 32'sd-0.09147347207865736, 32'sd0.05085742673172811, 32'sd-0.08902985189248236, 32'sd-0.12474096919315067, 32'sd-0.021179337894569224, 32'sd-0.03727733740858712, 32'sd0.045290712526473646, 32'sd0.02137302271378418, 32'sd-0.1595744650318592, 32'sd-0.06752198024930596, 32'sd0.035385627382344575, 32'sd0.11100331000157525, 32'sd0.08149806299990896, 32'sd0.022673686983469374, 32'sd-0.03213915393735027, 32'sd0.008345152504735357, 32'sd0.09547902809656279, 32'sd-0.13073950552938418, 32'sd0.05108952727565591, 32'sd-0.19363788589292494, 32'sd-0.14908268220007745, 32'sd0.07575884171304045, 32'sd-0.050319885921103855, 32'sd0.12042125252271506, 32'sd0.13771017324091495, 32'sd0.14319351337533784, 32'sd-0.08202952305351463, 32'sd-0.07117148213294092, 32'sd-0.11330168663155749, 32'sd-0.11775045026948348, 32'sd-0.04215080945902118, 32'sd-0.023279349313568738, 32'sd0.027757434152558696, 32'sd0.0393323113551106, 32'sd0.024766743330635672, 32'sd-0.06916008885939344, 32'sd0.060413658798103925, 32'sd0.053391877946374545, 32'sd0.045690262957983035, 32'sd0.06350897868034687, 32'sd0.02176117864412325, 32'sd0.029555948697400265, 32'sd-0.04650807330223057, 32'sd-0.057861605921508456, 32'sd0.07775967464406533, 32'sd0.026021953384292907, 32'sd-0.1376604960018968, 32'sd-0.200451321493273, 32'sd0.036015374857087064, 32'sd-0.01281197402184239, 32'sd0.046188354846344266, 32'sd0.13415494055464414, 32'sd0.07071831836284219, 32'sd0.138263154436285, 32'sd0.023209863046787953, 32'sd0.05642062591670353, 32'sd-0.08383125880622265, 32'sd0.017968102091053248, 32'sd0.09598132708941595, 32'sd0.051414001663168986, 32'sd0.04067577328712673, 32'sd-0.03492982604133661, 32'sd0.06423603451841661, 32'sd0.07453942069278766, 32'sd-0.008597068603496212, 32'sd-0.0015150020079436736, 32'sd-0.10724471766708339, 32'sd-0.010455549073531268, 32'sd-0.04677294582928072, 32'sd0.03740344491039019, 32'sd-0.0028784089839403683, 32'sd0.00030034538982010066, 32'sd-0.04459040980940287, 32'sd0.08636850145217993, 32'sd-0.19619001223854352, 32'sd-0.19453879304563418, 32'sd-0.1259432200218224, 32'sd0.0038477403856009996, 32'sd0.08730249337649773, 32'sd0.15441695673553632, 32'sd0.17695074451771978, 32'sd0.10841987183691044, 32'sd-0.013073015720050029, 32'sd-0.026582441499541722, 32'sd-0.009735881040276721, 32'sd-0.09751081244984161, 32'sd0.007152610938118622, 32'sd0.025428675407879377, 32'sd-0.05846468611845592, 32'sd0.01672510920023662, 32'sd0.0001540419825028713, 32'sd0.08539229786940931, 32'sd0.011481568249599032, 32'sd0.0006878291887869722, 32'sd-0.0026158363823199815, 32'sd0.03327951657051103, 32'sd-0.038879920049291715, 32'sd0.055421483349721135, 32'sd-0.030974780275998086, 32'sd0.047995661306560446, 32'sd-0.04443216148006862, 32'sd-0.029740717507122483, 32'sd-0.12275789204877646, 32'sd-0.2240609523271551, 32'sd-0.026596672073395305, 32'sd-0.06879789547950005, 32'sd0.04075965675842386, 32'sd0.14236725342741294, 32'sd0.11043595173736602, 32'sd0.05824781442958735, 32'sd0.012096890389148124, 32'sd-0.00799148448576253, 32'sd-0.022878598665901004, 32'sd-0.08110876120224103, 32'sd0.058655779826679584, 32'sd0.0007464755488207466, 32'sd0.06002736857372944, 32'sd-0.007415015922526762, 32'sd0.037474355458353883, 32'sd0.07636364188653343, 32'sd-0.07383209063653762, 32'sd-0.03871182936181057, 32'sd-0.035963727660119175, 32'sd0.018788408969383795, 32'sd-0.08022039992932488, 32'sd-0.07304265436260661, 32'sd-0.10559572692724287, 32'sd0.05715738231188085, 32'sd0.0275509121496764, 32'sd-0.018083819016144913, 32'sd-0.09512435875164317, 32'sd-0.17429682882317762, 32'sd-0.08792483880171992, 32'sd0.026474747017949163, 32'sd0.08757175517538389, 32'sd0.10510601614722571, 32'sd0.1880369452732042, 32'sd-0.013718782924911906, 32'sd-0.04814125243223269, 32'sd0.026754866749204513, 32'sd0.13297741681233088, 32'sd-0.09271446288013406, 32'sd0.034499080774834406, 32'sd-0.03140757060996053, 32'sd0.03606495628890194, 32'sd0.012611606681699378, 32'sd-0.1227064457675583, 32'sd-0.05030923631943627, 32'sd-0.11984107651238655, 32'sd-0.05757501344908143, 32'sd-0.16516998669551688, 32'sd-0.008517718663626661, 32'sd0.022850595895270387, 32'sd-0.00885013820479336, 32'sd0.012973419995206847, 32'sd0.04221112978057467, 32'sd-0.1104558792447656, 32'sd-0.26641501205939816, 32'sd-0.2290560009428543, 32'sd-0.07782248121013578, 32'sd-0.040541126280773915, 32'sd0.061982446558895, 32'sd-0.027805181376346615, 32'sd0.1083975112207649, 32'sd0.12099970029848801, 32'sd-0.06643347407922243, 32'sd-0.05262013126030697, 32'sd0.02593412420812764, 32'sd-0.016341310176469684, 32'sd-0.07418064726957659, 32'sd-0.0054765107176913035, 32'sd-0.019208651309666848, 32'sd0.0604364122804189, 32'sd0.037542327559589264, 32'sd0.03983339846910872, 32'sd0.015508175057355106, 32'sd-0.05885943620107223, 32'sd-0.005559614785982375, 32'sd-0.1065192988921232, 32'sd0.024581448615262007, 32'sd0.05919364735106015, 32'sd-0.0768809710789125, 32'sd-0.0934587030978163, 32'sd-0.04907360276495064, 32'sd-0.08124975690457242, 32'sd-0.2837880136012388, 32'sd-0.08665970337212245, 32'sd0.05114397396613948, 32'sd0.11398730426674426, 32'sd0.011817377295181548, 32'sd0.057718098954399256, 32'sd-0.055519697957617985, 32'sd0.034030341582517804, 32'sd0.03904762750583442, 32'sd0.0210143340940132, 32'sd-0.032035315850336935, 32'sd0.1406725514040904, 32'sd0.014261269808800154, 32'sd-0.0028892560560435953, 32'sd-0.09989738817676096, 32'sd-0.0748669779492865, 32'sd-3.551390515523722e-116, 32'sd0.0017219639135385722, 32'sd-0.05444668633074861, 32'sd-0.06942757025312965, 32'sd-0.03297714112353913, 32'sd-0.07134573712273051, 32'sd-0.06119120475687368, 32'sd-0.005899724558750088, 32'sd-0.0548791124286216, 32'sd-0.00870426082716355, 32'sd-0.19430777134003474, 32'sd-0.23039004893831094, 32'sd-0.17668661434075922, 32'sd0.040994188909117525, 32'sd0.08252306728017379, 32'sd0.07216171357773735, 32'sd0.12642684143787813, 32'sd0.04256784623421604, 32'sd0.12111631495990954, 32'sd-0.09535214310950585, 32'sd-0.0247759208835724, 32'sd-0.15371953835371316, 32'sd-0.07255936977796143, 32'sd-0.040143603169324873, 32'sd-0.09695205481481753, 32'sd-0.098127636536533, 32'sd-0.0509945602303694, 32'sd0.043938365340323124, 32'sd0.013614024208587703, 32'sd0.09199427418608977, 32'sd0.050331121939367805, 32'sd-0.040868915023775536, 32'sd-0.13556059952041055, 32'sd-0.10118434711924247, 32'sd-0.05765914551663688, 32'sd-0.03591086515003899, 32'sd-0.06776896318933591, 32'sd-0.135752024673015, 32'sd-0.19859951637704004, 32'sd-0.2048787258381763, 32'sd-0.037470239185544194, 32'sd0.1033202480909476, 32'sd0.03165752764666917, 32'sd0.004536152131726594, 32'sd0.08086647193454104, 32'sd-0.03890225401841975, 32'sd-0.003645626300201125, 32'sd-0.023735263182296934, 32'sd-0.08053960124614944, 32'sd-0.21643276813101087, 32'sd-0.03213668504776425, 32'sd0.04674745654545141, 32'sd0.08593260184295472, 32'sd0.04958499898533693, 32'sd0.07678041878415186, 32'sd0.053742735870375334, 32'sd0.0016670217426060412, 32'sd-0.036587979987515076, 32'sd-0.058195392937553166, 32'sd0.021378717431252598, 32'sd-0.08269853466888301, 32'sd-0.025685473963150542, 32'sd-0.04668829952802366, 32'sd0.10528377621799133, 32'sd-0.052724438239528756, 32'sd-0.11008887208373744, 32'sd-0.04716244301977125, 32'sd-0.09559998796431553, 32'sd0.17585050449171455, 32'sd0.1514755258913901, 32'sd0.15254771355220087, 32'sd0.02830727581016348, 32'sd0.06864758652775785, 32'sd0.0819268243023684, 32'sd-0.028922164392735993, 32'sd-0.02238516600415389, 32'sd-0.11099812746801553, 32'sd-0.13129463690272972, 32'sd-0.13998587249499278, 32'sd-0.042848467950901546, 32'sd0.07416836475229267, 32'sd-0.018910987671831754, 32'sd0.0781499820632307, 32'sd0.020126632970219303, 32'sd-1.4693062329198571e-124, 32'sd0.025171048220807266, 32'sd0.0024952109801194733, 32'sd0.05098571274594225, 32'sd-0.026610714979909262, 32'sd-0.07353052474752157, 32'sd0.0025267422529117833, 32'sd0.05203406443970177, 32'sd0.08300786044040087, 32'sd-0.06256324266558863, 32'sd-0.0763023099678695, 32'sd0.0014315522188207887, 32'sd0.17826045519591313, 32'sd0.11070628131540008, 32'sd0.07896861299056245, 32'sd0.05209414703058042, 32'sd0.06286344156645167, 32'sd-0.09575600322058819, 32'sd0.01818197067485877, 32'sd0.015443872259974399, 32'sd-0.08484988054584085, 32'sd0.03716431908722603, 32'sd-0.13399782013185224, 32'sd0.04580037227592119, 32'sd0.13371530053311695, 32'sd-0.011128261710215921, 32'sd0.008492727067398077, 32'sd-0.0024950749563946023, 32'sd-0.012089869154296851, 32'sd0.06963030486234166, 32'sd0.05266073934586863, 32'sd-0.027214013617125735, 32'sd-0.07674982932703449, 32'sd-0.05965154934525515, 32'sd-0.09045622955567176, 32'sd-0.09437558123396889, 32'sd0.004038487644721484, 32'sd0.008914144213798894, 32'sd-0.05151414012161788, 32'sd-0.10579398797427086, 32'sd0.10492551890984238, 32'sd0.08489408913692406, 32'sd-0.008603387859196001, 32'sd0.06175095184459222, 32'sd-0.05575167810818352, 32'sd-0.01651091511410463, 32'sd0.0779490225324285, 32'sd0.03306576043724371, 32'sd-0.043497220327757276, 32'sd0.051612651335042364, 32'sd0.07442372236542492, 32'sd0.06368694871040137, 32'sd0.11424712859611348, 32'sd-0.06459079224054022, 32'sd-0.046932216041554835, 32'sd-0.03663354252437142, 32'sd-0.03302002832110125, 32'sd-0.03344878679963444, 32'sd0.02831575427440462, 32'sd-0.0707201502659765, 32'sd-0.11061981811548181, 32'sd-0.1281969425237293, 32'sd-0.0005488753263665175, 32'sd-0.0682445163917489, 32'sd0.13628194279687847, 32'sd-0.02377127691945131, 32'sd-0.13779020039620057, 32'sd-0.10553380193879286, 32'sd-0.03320798394485101, 32'sd0.021357269445465718, 32'sd0.09552718305796483, 32'sd0.0672107793457655, 32'sd0.07786826836068887, 32'sd0.10879309935027598, 32'sd0.027261137812617468, 32'sd-0.14422032181768846, 32'sd-0.02106371122332912, 32'sd-0.11841021968908903, 32'sd0.00310096991632984, 32'sd-0.037249714429150566, 32'sd0.030166746107855077, 32'sd-0.0016719523206021665, 32'sd-0.05566182644249689, 32'sd0.024872495856178387, 32'sd2.984011469442441e-123, 32'sd-0.04281884834325188, 32'sd0.02000893147896624, 32'sd0.0023408989923391706, 32'sd-0.08942906389959235, 32'sd-0.050992458030018346, 32'sd-0.02272011514696404, 32'sd-0.029365251990133366, 32'sd-0.04807832303041411, 32'sd0.01652948755509271, 32'sd-0.11869434556456566, 32'sd0.02679347493672572, 32'sd-0.010281271938066234, 32'sd0.02020875087296379, 32'sd0.0433840515291852, 32'sd-0.028181101446995527, 32'sd-0.032832543880643335, 32'sd-0.0428671800308385, 32'sd-0.0853652859634928, 32'sd0.0918347865419159, 32'sd0.008583619422772025, 32'sd-0.010905036111252993, 32'sd-0.03205937984915893, 32'sd-0.03355775213461087, 32'sd-0.08581586146469303, 32'sd0.01213481916512429, 32'sd-0.0014277799689394021, 32'sd3.553713245152009e-122, 32'sd2.142286613692255e-116, 32'sd-3.972925445496038e-117, 32'sd-0.006975578949610026, 32'sd-0.073091533578401, 32'sd-0.12113764519531776, 32'sd-0.19272654167643544, 32'sd-0.027396225360482036, 32'sd-0.04801469152652971, 32'sd-0.06893710948820644, 32'sd-0.025733326889479075, 32'sd-0.05499095642109174, 32'sd-0.04611087178073587, 32'sd-0.1576301159336207, 32'sd0.07741560179932108, 32'sd0.02592758132856896, 32'sd-0.01787830747775879, 32'sd0.034553582800283554, 32'sd0.006435679931802812, 32'sd0.037565265163781364, 32'sd0.05771885555962895, 32'sd0.021712434990400698, 32'sd-0.06678172669558852, 32'sd0.0172273515658659, 32'sd-0.015051017388715839, 32'sd0.01576422373962277, 32'sd0.01774154296630109, 32'sd0.0003912127531433309, 32'sd4.864663249257479e-121, 32'sd7.568592217713429e-115, 32'sd-4.868277858135341e-123, 32'sd0.036894182816523645, 32'sd-0.006141406785739145, 32'sd-0.07730781626264804, 32'sd-0.11981444477357901, 32'sd-0.002240935251631085, 32'sd-0.06181259729816423, 32'sd-0.11936841488705466, 32'sd-0.09907065667606892, 32'sd-0.019467387267101288, 32'sd0.0002627362364295857, 32'sd0.011433075660210264, 32'sd-0.009683770330576444, 32'sd0.11505879169747668, 32'sd0.008698814406516321, 32'sd0.010823831065454185, 32'sd0.05874930468706749, 32'sd0.053257165274538, 32'sd0.04579838651134764, 32'sd0.07093114433690627, 32'sd0.020307903268598205, 32'sd-0.03805475583106028, 32'sd0.04865813620613905, 32'sd-0.006042858134450543, 32'sd0.04813198583242716, 32'sd0.0008906012775716615, 32'sd-5.637560927262124e-124, 32'sd7.059819962478974e-122, 32'sd1.077222281044353e-124, 32'sd-8.824412525128658e-120, 32'sd0.03393895520642883, 32'sd0.03673919644309346, 32'sd-0.05196178747815047, 32'sd-0.11998492569462538, 32'sd-0.07884996834025428, 32'sd0.0999088947416422, 32'sd0.12907753496191493, 32'sd0.07950149407403674, 32'sd0.0013338232369564525, 32'sd-0.058933564244764904, 32'sd0.07273568549528568, 32'sd0.1283798227624553, 32'sd-0.050810700500419505, 32'sd0.026692922313087137, 32'sd0.04113432007898991, 32'sd0.12188682548815839, 32'sd0.10669052777152437, 32'sd0.10717099714889117, 32'sd-0.01475228217893097, 32'sd0.002019203335242476, 32'sd0.01618590697808983, 32'sd0.024353440589577825, 32'sd-0.0035294188166756064, 32'sd6.853831486517139e-124, 32'sd1.6435415290358032e-127, 32'sd2.9064946071032736e-124, 32'sd7.160946484585685e-116, 32'sd-8.796330172855624e-125, 32'sd5.360320354674621e-116, 32'sd0.07639684796430046, 32'sd0.0025115573654057493, 32'sd-0.02261536502111449, 32'sd0.08798994872369717, 32'sd0.05901762634633665, 32'sd-0.051541909193142624, 32'sd0.05958586860455273, 32'sd0.08584263303412733, 32'sd-0.0035592150518832058, 32'sd0.013724309840809672, 32'sd-0.00045645334681834444, 32'sd0.038582976233803926, 32'sd0.029127497382215872, 32'sd0.011597561415025921, 32'sd0.024846610373999246, 32'sd-0.019564805586634947, 32'sd-0.03531908672002156, 32'sd0.04685916768847087, 32'sd0.0957333765019705, 32'sd0.10624638420482144, 32'sd-9.883228592657915e-121, 32'sd5.0151109122621836e-124, 32'sd1.293937020308293e-125, 32'sd-1.294573682985486e-126},
        '{32'sd-4.623930999104525e-123, 32'sd1.549413430546416e-119, 32'sd4.6568855300702144e-126, 32'sd-1.4337087978070613e-118, 32'sd4.356473927166638e-115, 32'sd3.3954779955136504e-122, 32'sd4.6195610000324806e-127, 32'sd-5.570637863032211e-115, 32'sd9.532155925571006e-120, 32'sd-1.8177765690062756e-123, 32'sd-4.7254051197110444e-123, 32'sd9.512481375479111e-120, 32'sd-0.09391372575453244, 32'sd-0.08631013676219108, 32'sd-0.0756199607683161, 32'sd-0.05952468845089372, 32'sd-1.4126061885853526e-124, 32'sd-4.2705592838754054e-126, 32'sd1.0342404397524594e-122, 32'sd3.1476915037747745e-119, 32'sd7.2328056620324574e-127, 32'sd4.514855284263552e-116, 32'sd1.0188004667818416e-124, 32'sd-5.094693253177587e-125, 32'sd-6.064475165047776e-126, 32'sd3.170182760547296e-126, 32'sd-5.168037318889037e-118, 32'sd1.0970047271351268e-119, 32'sd3.244421226574775e-121, 32'sd5.553313527269376e-126, 32'sd2.0676059072469508e-117, 32'sd-6.534392174306378e-117, 32'sd-0.045185032077266304, 32'sd-0.07975845344622448, 32'sd-0.008607825328093698, 32'sd-0.1284031238494566, 32'sd-0.031025037645750198, 32'sd0.06903617640766035, 32'sd0.04350333458136847, 32'sd-0.08447941820855631, 32'sd-0.08076600866652116, 32'sd-0.049190784681491635, 32'sd0.019328959389259794, 32'sd0.0725858523280165, 32'sd-0.003045965337628817, 32'sd0.00777541663157423, 32'sd0.01701698045421649, 32'sd-0.011495747404076107, 32'sd-0.1460887173497326, 32'sd-0.1174505960116593, 32'sd0.011226109884462392, 32'sd0.041640209500685706, 32'sd6.853197072765812e-125, 32'sd-1.780043971681699e-121, 32'sd8.615165282938275e-127, 32'sd-6.94791362439833e-124, 32'sd-1.349191567291176e-123, 32'sd-1.0127716196351918e-124, 32'sd-0.03424803878186208, 32'sd-0.0578350747138232, 32'sd0.0019203585630448027, 32'sd0.05483308173509278, 32'sd-0.1370802845749815, 32'sd0.057236992324791854, 32'sd0.058937398817411175, 32'sd0.12378152896881384, 32'sd0.10558326530577485, 32'sd-0.058520362546026314, 32'sd-0.028720171985489526, 32'sd-0.04433671889910119, 32'sd0.028547237816590333, 32'sd0.039972305958691515, 32'sd-0.1133614491699537, 32'sd-0.0798013463487427, 32'sd0.03222821789819077, 32'sd-0.041833290916482566, 32'sd-0.06982089995198218, 32'sd0.019234089900351463, 32'sd-0.055579516643722814, 32'sd-0.08901144471011045, 32'sd-0.0665319369353923, 32'sd-0.087306615941121, 32'sd6.848156014230048e-126, 32'sd5.395042624382355e-127, 32'sd3.0058611522590715e-120, 32'sd9.812934294163562e-121, 32'sd-0.03905792135703172, 32'sd-0.0501634989173912, 32'sd0.0007586387927903484, 32'sd-0.14707058424207373, 32'sd-0.24509165984344258, 32'sd-0.15006111427901203, 32'sd-0.04957486391584145, 32'sd-0.011348010570707693, 32'sd0.04756179670545912, 32'sd-0.040314163964386605, 32'sd-0.01758972399793736, 32'sd0.03320397226844511, 32'sd0.028539828151724123, 32'sd-0.03303021050414839, 32'sd-0.004708853663626064, 32'sd-0.04760029158000871, 32'sd-0.021327899377477044, 32'sd0.03036022704943649, 32'sd0.046093262628693635, 32'sd-0.0009373246539480752, 32'sd-0.07456519356506146, 32'sd0.05861468511141961, 32'sd-0.09187780322924147, 32'sd-0.08804030284524193, 32'sd-0.0543682713352912, 32'sd8.621977441987611e-117, 32'sd5.396391914092754e-125, 32'sd0.042562678854740174, 32'sd0.05924266233278199, 32'sd-0.11064972073497671, 32'sd-0.013180376885348849, 32'sd-0.06336490799283934, 32'sd-0.0032655495014941144, 32'sd-0.07218676752802486, 32'sd0.062101710131849584, 32'sd0.13431262188677215, 32'sd0.1610739882892237, 32'sd0.08268113382025533, 32'sd0.004657685287987665, 32'sd0.03245781279417616, 32'sd0.14734988790615097, 32'sd0.09912191975743205, 32'sd-0.11063678060749259, 32'sd-0.06987670247978345, 32'sd-0.05912136908014426, 32'sd-0.02044811504241141, 32'sd0.12702766415943498, 32'sd0.04800210972744815, 32'sd0.06738989721953442, 32'sd-0.017693360416004007, 32'sd0.009057531885151468, 32'sd-0.023413780262147417, 32'sd-0.04982219063474162, 32'sd0.05787713737849982, 32'sd2.774822766906043e-120, 32'sd-0.024529758606435758, 32'sd0.03366006778817135, 32'sd0.03200060640432191, 32'sd0.0976424539107853, 32'sd0.04500117400467474, 32'sd-0.06684007953459359, 32'sd0.03663459522023018, 32'sd0.12043018306988326, 32'sd0.10832905171859938, 32'sd0.15180881864756923, 32'sd0.0996818878090917, 32'sd0.08918713038982991, 32'sd-0.028739243529352115, 32'sd-0.039547318573760155, 32'sd0.012169279985587927, 32'sd-0.009296018887186572, 32'sd-0.13003315543909108, 32'sd-0.05050923146219685, 32'sd-0.14364626426475852, 32'sd-0.024003925518563105, 32'sd-0.0469840730459605, 32'sd0.00857167102434765, 32'sd0.09128209719324308, 32'sd0.042955247288625466, 32'sd-0.008510745789219166, 32'sd-0.04881256508908346, 32'sd-0.03425732983022939, 32'sd-4.277955086667472e-121, 32'sd-0.07021957025136365, 32'sd0.009144752029787588, 32'sd0.021499724248196055, 32'sd-0.01196813759186309, 32'sd-0.02537313620205344, 32'sd0.10363736225570809, 32'sd0.10598581535198047, 32'sd0.06616087399373786, 32'sd0.09160090177601041, 32'sd0.053303531752528395, 32'sd0.17541708600941264, 32'sd0.07495887965623207, 32'sd0.03465760252853549, 32'sd-0.04344210340817885, 32'sd-0.03307364583489054, 32'sd-0.07935209833244335, 32'sd-0.012249528990944482, 32'sd-0.12659620884026368, 32'sd0.02804361457543395, 32'sd-0.12111122007738627, 32'sd-0.08202777113473173, 32'sd-0.0840045154708998, 32'sd0.03716411066348896, 32'sd0.08879105446327272, 32'sd-0.05351089641953869, 32'sd-0.052444120149312975, 32'sd0.04326506236609246, 32'sd-0.05281940428933796, 32'sd0.039536038349441076, 32'sd0.02665847751398297, 32'sd-0.07492748603179432, 32'sd-0.0005996108963745551, 32'sd0.10793831446389714, 32'sd-0.021379926426365076, 32'sd0.01395862802272827, 32'sd-0.011655960609510824, 32'sd0.03757897692451613, 32'sd0.08387152398869939, 32'sd-0.005219334161128827, 32'sd0.0409631860123245, 32'sd0.12894224650200342, 32'sd0.027222416440026147, 32'sd-0.05129897793431953, 32'sd-0.03711953800107243, 32'sd0.07459923384396137, 32'sd-0.010112164492436508, 32'sd0.010447129068932404, 32'sd-0.009051822574646583, 32'sd0.12308021625515807, 32'sd0.14032939587413493, 32'sd0.02997914384488085, 32'sd-0.07355818394401775, 32'sd0.04627823795762278, 32'sd0.08968953553863089, 32'sd-0.02873693911930468, 32'sd-0.03753625372947863, 32'sd0.0062082492946372615, 32'sd-0.08191309779286704, 32'sd-0.010390545708491043, 32'sd-0.07217288749555408, 32'sd0.02349519061038616, 32'sd-0.007424356742337499, 32'sd-0.022881535467725662, 32'sd0.08801544053217275, 32'sd0.1713161903901985, 32'sd0.11685740071704638, 32'sd0.01192434741689817, 32'sd-0.051605776259235146, 32'sd-0.010801581531299427, 32'sd0.10321748327695367, 32'sd0.052689318941209026, 32'sd0.009690405048489474, 32'sd-0.042415550952278495, 32'sd-0.0560809547252212, 32'sd-0.001762225467896605, 32'sd-0.05699633508223839, 32'sd-0.009729215827745984, 32'sd0.014839535535599498, 32'sd-0.04232075674664601, 32'sd-0.08359114712458934, 32'sd0.05297972159312726, 32'sd0.06932083660832743, 32'sd0.1107472624240101, 32'sd-0.11605796627814789, 32'sd-0.024102134534151668, 32'sd-0.05122196077741608, 32'sd0.032161249537574065, 32'sd-0.05112286686998579, 32'sd-0.005936886178250401, 32'sd0.04241692606460404, 32'sd-0.03536228062709009, 32'sd0.15650524779914143, 32'sd0.1541979429487752, 32'sd0.07081853510579539, 32'sd-0.1411963434889722, 32'sd-0.35304884928880775, 32'sd-0.17645393882091825, 32'sd-0.018422700449270493, 32'sd0.0022869335155855206, 32'sd0.044344198742051984, 32'sd-0.037445979527110616, 32'sd-0.01621292238782528, 32'sd0.14914505095859515, 32'sd-0.05886544119689598, 32'sd-0.09329078886113339, 32'sd-0.0670059843891697, 32'sd0.04455078334956921, 32'sd0.10024038118352341, 32'sd0.031811227425462475, 32'sd0.06475081671238246, 32'sd0.036878495956020975, 32'sd-0.054703625643105026, 32'sd-0.12536836307376603, 32'sd-0.15504794813117423, 32'sd0.08767423580570928, 32'sd0.006301557755495724, 32'sd0.10162125546876517, 32'sd0.11606110052807316, 32'sd0.0800254682502393, 32'sd0.21236060960909514, 32'sd0.1946666503254671, 32'sd0.018196072383770946, 32'sd-0.16438461476501912, 32'sd-0.22135996261036905, 32'sd-0.16830633183788304, 32'sd0.10072818339882292, 32'sd-0.04854057938933814, 32'sd-0.025052743465423005, 32'sd0.008932567726356803, 32'sd0.11086290063242807, 32'sd-0.015212599254997006, 32'sd-0.008174018198917346, 32'sd-0.049637445260986915, 32'sd-0.06237148560286162, 32'sd0.0914964529984983, 32'sd0.14236282081251606, 32'sd-0.024347174424182296, 32'sd-0.03176009426062136, 32'sd0.06069025684997109, 32'sd-0.07324694595093066, 32'sd-0.08791953609549205, 32'sd-0.01481763500109581, 32'sd-0.04580718841968223, 32'sd0.04579421549309302, 32'sd-0.013568743749900693, 32'sd-0.033444777458202235, 32'sd0.10285294826744273, 32'sd0.13759108606154138, 32'sd0.17080826336131713, 32'sd0.07969715521854104, 32'sd-0.013139520153476773, 32'sd-0.07794871849058455, 32'sd-0.009679529652821418, 32'sd-0.0057920967283413, 32'sd-0.023198254711583422, 32'sd-0.05789392783478247, 32'sd-0.028182443294404964, 32'sd-0.047588105841784654, 32'sd0.039386496827932015, 32'sd-0.05558499264242389, 32'sd-0.02023331517181963, 32'sd-0.11584466487116897, 32'sd0.010226476473764368, 32'sd0.0693362076458463, 32'sd-0.033307275754318987, 32'sd0.0977550477088042, 32'sd-0.09103198608685413, 32'sd-0.07316878085115713, 32'sd-0.049238214904045875, 32'sd-0.13444157052361924, 32'sd0.047329688092426256, 32'sd-0.07055315445967662, 32'sd0.03658158984815595, 32'sd0.1823723386103775, 32'sd0.18295186915101228, 32'sd0.08918763261271354, 32'sd0.2033337545424886, 32'sd0.006076942271734678, 32'sd0.09493198118028673, 32'sd0.12060566438661746, 32'sd0.06996121115209226, 32'sd-0.09149531352574708, 32'sd-0.08607860527727176, 32'sd-0.07633658320100516, 32'sd-0.06109189536035465, 32'sd-0.08951009640223273, 32'sd0.003962666362927504, 32'sd-0.04911178082218784, 32'sd-0.0056032589985536615, 32'sd-0.17400367095906877, 32'sd-0.04882551856388908, 32'sd0.05850893272015398, 32'sd-0.016449603435592878, 32'sd-0.018214239981320213, 32'sd-0.08013712113792144, 32'sd-0.05460915807178699, 32'sd0.012618186738316405, 32'sd-0.11270991030157594, 32'sd0.025369290294088027, 32'sd-0.07171755567248751, 32'sd0.04895436221602678, 32'sd0.11454345846144137, 32'sd0.05816520208564436, 32'sd0.05069098477374763, 32'sd0.10538019152276644, 32'sd0.1484594309921115, 32'sd0.21844034994807865, 32'sd0.01719266743056445, 32'sd0.0710348548952712, 32'sd0.008600046044787556, 32'sd0.02226958090662137, 32'sd-0.10667379294861687, 32'sd-0.048418806602512965, 32'sd-0.003716901856849939, 32'sd0.13099829067750748, 32'sd-0.0663072475165354, 32'sd-0.04902252089693935, 32'sd0.05848050983900438, 32'sd-0.11543751588953911, 32'sd-0.10632313095162531, 32'sd0.018896655052508888, 32'sd0.05812107825978606, 32'sd-0.11437900181245754, 32'sd0.06276086941881594, 32'sd-0.052496449483294426, 32'sd0.00876338560745874, 32'sd-0.10200646424617715, 32'sd-0.06463137847789749, 32'sd0.13138506056078889, 32'sd0.09431114789251083, 32'sd0.03389848953014858, 32'sd0.014497859718890574, 32'sd0.06548868363778311, 32'sd0.0392429388015682, 32'sd0.06484271671640551, 32'sd0.001776207330267139, 32'sd-0.06671619057754766, 32'sd-0.002861366896030529, 32'sd-0.06447705559282708, 32'sd-0.09479955042310426, 32'sd0.10645318993819457, 32'sd0.09065065677352954, 32'sd-0.05240794502988784, 32'sd-0.04954462217250642, 32'sd0.015444574169478321, 32'sd-0.01993555414844273, 32'sd-0.063974299797899, 32'sd-0.03921401440177973, 32'sd0.08800359851173713, 32'sd0.005582096089547033, 32'sd-0.0072519471391310425, 32'sd0.07645561306081, 32'sd0.011134414655420864, 32'sd-0.07535350817011757, 32'sd-0.046111346387973026, 32'sd-0.05002505889338046, 32'sd0.05938317686153527, 32'sd0.03762169772852311, 32'sd-0.06053991983479075, 32'sd-0.06640801242046608, 32'sd0.1161375556402319, 32'sd0.11981759909422417, 32'sd0.16015046359495652, 32'sd0.055853149097485864, 32'sd0.08707453793206635, 32'sd0.00590883890941332, 32'sd-0.02630500150704106, 32'sd0.04617691091399669, 32'sd-0.054687020122306064, 32'sd0.0018350226566478814, 32'sd0.05559048497058243, 32'sd0.035179582244830046, 32'sd-0.03832789591197569, 32'sd0.014255175712810686, 32'sd-0.052495827865184565, 32'sd0.04261676474542926, 32'sd0.040455700001783355, 32'sd-0.03180618280131027, 32'sd0.04161670191351337, 32'sd0.04205481259122395, 32'sd0.03341238920057051, 32'sd-0.02474935776170409, 32'sd-0.16009206781413102, 32'sd-0.0015783969373155174, 32'sd0.024413298346015053, 32'sd-0.1343140725675718, 32'sd-0.08327555211250513, 32'sd-0.09882369479732893, 32'sd-0.10275312549611904, 32'sd0.11462266227817573, 32'sd0.15758802597499777, 32'sd0.0840530182175427, 32'sd0.0730041482927201, 32'sd-0.11094773758980062, 32'sd-0.03390756126907035, 32'sd0.04811149497192697, 32'sd-0.12886622810478568, 32'sd0.06923337425531985, 32'sd0.03655306659617483, 32'sd0.025998603943809623, 32'sd-0.06747366984620469, 32'sd-0.09118928914471498, 32'sd0.09983602830221963, 32'sd0.03009108321179587, 32'sd0.009749272736900681, 32'sd0.07452578173700672, 32'sd0.030420559175268716, 32'sd2.6820924255619847e-115, 32'sd-0.003296315129500217, 32'sd0.0016231876329127972, 32'sd0.04982006102397521, 32'sd-0.04297992773066165, 32'sd-0.03321439493888892, 32'sd0.0004928003214618085, 32'sd-0.19231496805173648, 32'sd-0.08671047962164692, 32'sd-0.03183054675116069, 32'sd0.1214338963270753, 32'sd0.07943234784559049, 32'sd0.008590488221499746, 32'sd0.05866182035993936, 32'sd0.06056133143330911, 32'sd-0.06176617382637231, 32'sd0.046707567732321195, 32'sd-0.2161707238261382, 32'sd-0.09125325515705841, 32'sd-0.009150348668578287, 32'sd0.07135972956711098, 32'sd-0.009256876576041575, 32'sd0.04595766649373873, 32'sd-0.013591750242691684, 32'sd0.1215549227577316, 32'sd-0.010402508983882413, 32'sd-0.07878423283641814, 32'sd-0.07908450868841872, 32'sd-0.10270097508815487, 32'sd0.08446278905841069, 32'sd-0.004015877390524237, 32'sd0.05395764635357323, 32'sd-0.07445446625250518, 32'sd-0.033640518832653815, 32'sd0.05463378992492346, 32'sd-0.08721816027433311, 32'sd-0.08169201165333939, 32'sd0.07486827347918446, 32'sd-0.017091237534429513, 32'sd-0.017603376720813364, 32'sd0.00639748594477856, 32'sd0.03204244742172148, 32'sd0.07178487160049568, 32'sd-0.08540030352961632, 32'sd-0.1693517753041934, 32'sd-0.21005479705079846, 32'sd-0.15046523902768377, 32'sd-0.019888270178874463, 32'sd0.08268455596086874, 32'sd0.023163100010281237, 32'sd-0.09985109941099345, 32'sd-0.0561271207084113, 32'sd0.1180501505048832, 32'sd0.036540370046289516, 32'sd0.01963643161633199, 32'sd-0.08442473295471212, 32'sd-0.08763810503869839, 32'sd0.04512308956192816, 32'sd-0.020014165178200122, 32'sd0.12023832755448208, 32'sd-0.08303411329763818, 32'sd0.014209620994427274, 32'sd0.06660451740092357, 32'sd-0.021157962855948127, 32'sd0.10538431407208336, 32'sd0.1199625982715188, 32'sd-0.04494446572053335, 32'sd-0.09636283446028589, 32'sd-0.01903709669145347, 32'sd0.131130365595847, 32'sd0.0327309937517749, 32'sd0.13740182938179465, 32'sd-0.12338034778059793, 32'sd-0.24504237839471835, 32'sd-0.13064087565543248, 32'sd-0.09105526664879113, 32'sd0.07608347874279289, 32'sd0.08899248167700743, 32'sd0.09142499899354874, 32'sd-0.04663032480921686, 32'sd0.01451816277481194, 32'sd-0.0683318256253534, 32'sd0.020682695140268475, 32'sd-0.10199185059717378, 32'sd8.689459024853579e-127, 32'sd0.0760285206421125, 32'sd-0.0011833008571071988, 32'sd0.005180689749190124, 32'sd0.05157673747791978, 32'sd-0.07922766140569241, 32'sd-0.03549372243120131, 32'sd0.0027375158719669976, 32'sd0.11255756388845257, 32'sd0.07946074852352933, 32'sd0.0429080042208083, 32'sd0.053947109783174345, 32'sd-0.04042644157469542, 32'sd-0.01496029211570518, 32'sd0.06909246888511493, 32'sd0.07480031050626357, 32'sd-0.04931503479218743, 32'sd-0.08625686276252433, 32'sd-0.04778812692525403, 32'sd-0.03864622367711202, 32'sd0.15767596978698256, 32'sd0.012862437300447293, 32'sd0.04099973357616554, 32'sd0.07054938869585085, 32'sd-0.039030186110696696, 32'sd-0.04454593115988734, 32'sd7.170553945941778e-05, 32'sd-0.08010346584940459, 32'sd-0.06313211666717151, 32'sd-0.09290605949985764, 32'sd-0.046708380633292856, 32'sd0.06520004776195201, 32'sd-0.0011406314711534832, 32'sd-0.029968562887297344, 32'sd0.028326899771576573, 32'sd0.10571545310240334, 32'sd0.0860075491877154, 32'sd0.09386087438598746, 32'sd-0.05011154915977902, 32'sd-0.07611640820812474, 32'sd-0.1532660669331857, 32'sd-0.05910014413934812, 32'sd0.015346082739730205, 32'sd0.2549299795635999, 32'sd0.02853285154500029, 32'sd0.012442891049466278, 32'sd-0.02688907013030464, 32'sd0.025643249372630253, 32'sd0.09897967057661887, 32'sd0.13589075350656749, 32'sd0.06198036570630989, 32'sd0.027765410866165973, 32'sd-0.05582265356045176, 32'sd-0.03185171851255871, 32'sd0.03436636220094451, 32'sd-0.02798436928238954, 32'sd-0.08025514456350538, 32'sd0.06086495757306238, 32'sd0.02705201218930871, 32'sd0.019567737706896075, 32'sd-0.03529019713582814, 32'sd-0.16146532019280097, 32'sd-0.11455771175063473, 32'sd0.059611632537624956, 32'sd0.07416969271270829, 32'sd0.0457999530288883, 32'sd0.1240565156751605, 32'sd0.047880638633971205, 32'sd-0.055060002081581655, 32'sd-0.12309747607834304, 32'sd0.01950859446604505, 32'sd0.03761098374308249, 32'sd0.045591106829034354, 32'sd0.016368641078534498, 32'sd0.10103353920776256, 32'sd0.035654869319780326, 32'sd0.08905647019227571, 32'sd0.051685684240349354, 32'sd0.039118165693969385, 32'sd0.11873371149084538, 32'sd-0.048053698853325034, 32'sd0.021647790260385314, 32'sd-0.014407498774948931, 32'sd-0.06477029820876022, 32'sd7.204287061710062e-122, 32'sd-0.08233522768796678, 32'sd0.07922136745942522, 32'sd-0.0008941445108500758, 32'sd0.10449151069973199, 32'sd-0.02189995923963861, 32'sd-0.03850816343756476, 32'sd-0.0008719995253884155, 32'sd-0.004003661539307073, 32'sd0.023462446726658034, 32'sd-0.024551496901361186, 32'sd0.007808403600016389, 32'sd0.005158410427645053, 32'sd0.06738420966018603, 32'sd-0.039469327214177945, 32'sd-0.07545942961498556, 32'sd0.09343698303047111, 32'sd0.08314745277831417, 32'sd0.06194785482398006, 32'sd0.16581435295646735, 32'sd0.012485658880287544, 32'sd0.04049190863168544, 32'sd0.05854488522791949, 32'sd-0.027616822410499967, 32'sd-0.10063784464871432, 32'sd-0.08191511011056232, 32'sd-0.0824823388649068, 32'sd-1.2038786280253566e-120, 32'sd3.6203516034168517e-122, 32'sd-2.150222966820401e-114, 32'sd-0.012647105939925447, 32'sd-0.11514947115336645, 32'sd-0.10144122881275162, 32'sd-0.10562585300016339, 32'sd-0.05477237009558161, 32'sd0.03678883501555147, 32'sd-0.010052179050816158, 32'sd0.03914745969476788, 32'sd-0.006534758133416301, 32'sd0.07869910005918437, 32'sd0.0372279364585457, 32'sd0.08316585941189661, 32'sd-0.10770600369610918, 32'sd0.011925615018822104, 32'sd-0.005734891325421604, 32'sd0.017622542826667812, 32'sd0.08755464324514925, 32'sd0.09876021955072396, 32'sd0.05538066101442363, 32'sd-0.012521462805261297, 32'sd0.0647035860803245, 32'sd0.059037581215224844, 32'sd-0.019493729607479957, 32'sd-0.048497757061565845, 32'sd-0.06894175884510792, 32'sd3.546892165420612e-122, 32'sd3.206972253809323e-119, 32'sd-3.7114347725819405e-120, 32'sd0.04667219336805518, 32'sd-0.10828261961000182, 32'sd0.05764366665076213, 32'sd-0.012960926636113534, 32'sd-0.1460780985502841, 32'sd-0.13339680436339682, 32'sd-0.049813328635328925, 32'sd0.07728354874160306, 32'sd0.06920236965552481, 32'sd0.07539427665499907, 32'sd0.056051548699771025, 32'sd0.025523885749870353, 32'sd-0.06023301744969952, 32'sd0.08927588553960965, 32'sd-0.08255956033715241, 32'sd0.0374584464924939, 32'sd0.029888273778826774, 32'sd0.03387298669835896, 32'sd0.007037967458292037, 32'sd-0.07377048972372453, 32'sd-0.03754737141172916, 32'sd0.017070831813447696, 32'sd-0.006790270935300843, 32'sd-0.11243313088564433, 32'sd-0.04101096547506352, 32'sd1.723238036017202e-125, 32'sd-7.01037350062688e-116, 32'sd-2.0973162731293997e-124, 32'sd-1.6503097864817195e-119, 32'sd-0.03758721589006595, 32'sd-0.09144740444080605, 32'sd-0.1269821920815692, 32'sd-0.02651100969089915, 32'sd0.0002184723241099606, 32'sd0.10150860132437743, 32'sd-0.0804507675291323, 32'sd-0.03396295804785196, 32'sd0.031833676613578936, 32'sd0.12896391426133164, 32'sd-0.025181293728227035, 32'sd0.02111302133490943, 32'sd0.046796969919260065, 32'sd-0.003845914226243194, 32'sd0.10208721979893942, 32'sd-0.027099800325832837, 32'sd-0.02706004056911829, 32'sd0.033290933507538915, 32'sd0.014212851325444573, 32'sd0.0016328618985172049, 32'sd0.02918779696663182, 32'sd0.06914470436346919, 32'sd-0.05867814442929009, 32'sd-2.3661215450336176e-118, 32'sd-1.078736338124847e-124, 32'sd-3.165768108578592e-120, 32'sd3.3122535143281506e-122, 32'sd1.194783656648207e-121, 32'sd-1.0347854681408892e-120, 32'sd-0.00783241341967864, 32'sd-0.08642046475984896, 32'sd-0.0868535958231665, 32'sd-0.1015540039366501, 32'sd-0.02858307501379818, 32'sd0.06508646375118678, 32'sd0.08135869014915997, 32'sd-0.05228949328908758, 32'sd0.0452038809374335, 32'sd0.01647923329863423, 32'sd-0.04316430755616572, 32'sd-0.0844783439221961, 32'sd-0.11150648013755447, 32'sd-0.04269577496039759, 32'sd-0.034718349849923495, 32'sd0.01351327858485556, 32'sd0.030077435326187195, 32'sd-0.13324387988383582, 32'sd-0.08227513337263241, 32'sd-0.031667574716951245, 32'sd-4.314710845067995e-125, 32'sd1.0752649196070771e-121, 32'sd1.144926066783627e-120, 32'sd-5.2640832127582545e-120},
        '{32'sd-3.5502677824488845e-119, 32'sd-7.072355669930852e-115, 32'sd-6.211286067885274e-127, 32'sd5.309286526635024e-117, 32'sd-1.046041687084867e-120, 32'sd2.872743517212762e-114, 32'sd-4.914972029442641e-117, 32'sd-1.198508656806461e-122, 32'sd1.181610139121439e-116, 32'sd-3.1366896436502027e-123, 32'sd4.2845391139733274e-125, 32'sd-4.556027630312202e-118, 32'sd0.041603584893698496, 32'sd0.09427929118724468, 32'sd0.07392584298471153, 32'sd0.013780016136292131, 32'sd1.2670486314023798e-122, 32'sd-1.4179499365042462e-121, 32'sd2.026646542962708e-125, 32'sd1.2422725584529878e-122, 32'sd-5.691091010104585e-123, 32'sd1.128284167048965e-119, 32'sd3.7941641271518735e-117, 32'sd-1.1599654496642495e-121, 32'sd-2.264023016540429e-120, 32'sd-1.802038451684928e-125, 32'sd-2.0828418043611438e-119, 32'sd-1.718962622894927e-125, 32'sd8.06587633620706e-118, 32'sd7.050809438673415e-124, 32'sd7.536723899160601e-118, 32'sd9.143505255117798e-125, 32'sd-0.005838964895366798, 32'sd0.025618514601179948, 32'sd0.14158290779074686, 32'sd0.09920657092841564, 32'sd0.05472009632532598, 32'sd0.08004326163854136, 32'sd-0.01653576721380181, 32'sd0.047059483730557274, 32'sd0.027115551329365092, 32'sd0.0397383681949938, 32'sd-0.055445745417760074, 32'sd0.05110488871568899, 32'sd-0.03522205138052197, 32'sd0.02582276289120577, 32'sd0.02747931783669602, 32'sd0.05615987421375007, 32'sd0.0013042917107391886, 32'sd0.11288481005493056, 32'sd0.026033864531162923, 32'sd0.04527822880395795, 32'sd-2.0526452375577489e-128, 32'sd6.812549768653982e-121, 32'sd1.580485779584317e-127, 32'sd-8.423517183879579e-117, 32'sd3.461485470459258e-119, 32'sd-2.941894528822352e-116, 32'sd0.07432563249410318, 32'sd0.040243305550814144, 32'sd0.03917288416093552, 32'sd-0.0011978417288437673, 32'sd0.011727969820502757, 32'sd0.060167795186576174, 32'sd0.10629820728769786, 32'sd-0.03824153225878257, 32'sd-0.07397152905968805, 32'sd-0.0312753035492138, 32'sd0.07217551719688911, 32'sd-0.0503588217900023, 32'sd0.020283871857209593, 32'sd0.037406602354087236, 32'sd-0.019519552019554194, 32'sd-0.05061970081562519, 32'sd0.07160748761463993, 32'sd0.059260487454629494, 32'sd0.010631828074220133, 32'sd0.07549871846197133, 32'sd0.0919656091304041, 32'sd0.12541438024570414, 32'sd0.031162302224416523, 32'sd0.0760513395077252, 32'sd-2.4849366852163586e-118, 32'sd-2.672800970972401e-124, 32'sd-4.5186398520002147e-125, 32'sd4.873138025334387e-123, 32'sd-0.0797721194325064, 32'sd0.03540129761784789, 32'sd0.01910653119941039, 32'sd-0.12300925985863174, 32'sd-0.003635301585292764, 32'sd-0.021401254601962082, 32'sd0.059380616368490444, 32'sd0.05248680061303563, 32'sd-0.008830717841952324, 32'sd0.04237137861413835, 32'sd-0.06478596707515055, 32'sd-0.04782905844963342, 32'sd-0.09103979822252277, 32'sd-0.046717299957100916, 32'sd-0.04894884580967372, 32'sd-0.09272069843129596, 32'sd0.1223023002991136, 32'sd-0.020078006651248155, 32'sd0.016589272903724073, 32'sd0.10600091189974252, 32'sd-0.013660829221540995, 32'sd-0.16395690096863758, 32'sd0.007055663138125004, 32'sd-0.04482408735666993, 32'sd0.0227925740884268, 32'sd-9.667018295052996e-124, 32'sd3.4799028171587475e-116, 32'sd0.028216775431644785, 32'sd0.007139673082188997, 32'sd0.0003714619074414387, 32'sd-0.08406396150701223, 32'sd-0.028197855410946125, 32'sd0.04658397440687743, 32'sd0.11539837477561006, 32'sd0.05442390041980925, 32'sd0.0887791959609218, 32'sd0.011692960262729127, 32'sd0.0911730826603991, 32'sd0.15663990298939892, 32'sd0.17709465475252076, 32'sd-0.004037701953530479, 32'sd-0.023641062177688226, 32'sd-0.13649603464863191, 32'sd-0.09047302783772533, 32'sd0.021883508255295375, 32'sd-0.0025637727503376078, 32'sd-0.04050913891288619, 32'sd0.12438208300552853, 32'sd0.021887001403367443, 32'sd-0.04279668441568743, 32'sd-0.06590966960100911, 32'sd0.015733714175907722, 32'sd0.004895061309980519, 32'sd0.022712814008306343, 32'sd-2.430366760814319e-115, 32'sd0.08178355094034216, 32'sd-0.0246918545459369, 32'sd-0.027411640989774375, 32'sd0.0449690270360683, 32'sd0.07514790643014675, 32'sd0.06680648557482433, 32'sd0.19175868439903468, 32'sd0.08334121741645253, 32'sd-0.02705167516196924, 32'sd0.12679490998239507, 32'sd0.04378359465595527, 32'sd0.11271989346941617, 32'sd0.10026749741787133, 32'sd-0.045387283039392705, 32'sd0.03697600851894559, 32'sd0.11585256260674652, 32'sd-0.08551451465879502, 32'sd0.001664993979677544, 32'sd0.0660811467687929, 32'sd0.03487721432419814, 32'sd-0.05180642593922548, 32'sd0.01729113562387331, 32'sd-0.07997790829182351, 32'sd-0.09241366098234588, 32'sd-0.025062643949276354, 32'sd-0.011566572585298442, 32'sd0.017920972154565878, 32'sd-1.3059305006138494e-123, 32'sd0.020719739067123395, 32'sd0.04444396179092641, 32'sd0.01856454533847385, 32'sd0.10040085419199718, 32'sd0.006663942467139324, 32'sd-0.02344375317987135, 32'sd0.04471775659355957, 32'sd0.007563673619520993, 32'sd0.050521353538528574, 32'sd-0.05464866866561278, 32'sd-0.03353102200285044, 32'sd0.00244690650644801, 32'sd-0.048044761407423524, 32'sd0.05600964811228129, 32'sd0.1181251127124799, 32'sd0.06366739137284702, 32'sd0.15995013900326144, 32'sd0.09093922431752578, 32'sd0.02720241843427529, 32'sd0.003562261747528563, 32'sd0.04145585945973074, 32'sd-0.013735543762266206, 32'sd-0.0873668153414062, 32'sd-0.07574809618383797, 32'sd0.05823920625893238, 32'sd0.04995901815357751, 32'sd-0.005558890640385713, 32'sd0.05175321088955504, 32'sd0.03449895677395268, 32'sd0.08134399063574481, 32'sd0.017921937780978007, 32'sd0.035399390370487546, 32'sd-0.06220795129648507, 32'sd-0.029577512172511304, 32'sd-0.023826262103193184, 32'sd-0.04432082603903991, 32'sd-0.1185671520882836, 32'sd-0.026886258076753235, 32'sd-0.18238202812061152, 32'sd-0.1431959518750872, 32'sd-0.022644090460858704, 32'sd0.02069809235863896, 32'sd0.07061132873766966, 32'sd0.05031457537343487, 32'sd0.11152778995439322, 32'sd0.11949988541837954, 32'sd0.07676421109558158, 32'sd0.008810798562358078, 32'sd0.07516737047462149, 32'sd0.0073559462629482425, 32'sd-0.08450543757238316, 32'sd-0.07395018623686826, 32'sd-0.02049139019260137, 32'sd0.010042674417409931, 32'sd0.103142739272712, 32'sd0.06085034942834092, 32'sd-0.04710102342129773, 32'sd0.006603334151930225, 32'sd-0.05873129657873025, 32'sd0.006621658639421438, 32'sd-0.09979015659472153, 32'sd-0.022203935316618482, 32'sd-0.029333762061509103, 32'sd0.14311773439376274, 32'sd-0.1249078306166178, 32'sd-0.06836337478530302, 32'sd-0.010475223112901555, 32'sd-0.12052787951703842, 32'sd-0.009976663633624745, 32'sd-0.03333159637677286, 32'sd-0.0034571783816014982, 32'sd-0.0974173018261565, 32'sd0.032948917785478066, 32'sd-0.07083294447485199, 32'sd0.04174209379528556, 32'sd0.025264366121085895, 32'sd0.058143464246429126, 32'sd0.08879660790390966, 32'sd0.037500595959001286, 32'sd-0.1260516636133636, 32'sd-0.07838796225809903, 32'sd0.01582153875089079, 32'sd-0.05142196348309954, 32'sd0.05124338059555944, 32'sd0.009832741961107302, 32'sd0.038262993981405716, 32'sd0.10575005935189916, 32'sd0.06678489468401493, 32'sd-0.1322911677508437, 32'sd-0.07044154497292937, 32'sd-0.0897816933983356, 32'sd-0.05996448473405117, 32'sd-0.1265748692945251, 32'sd-0.03347533737635694, 32'sd0.012886558603209187, 32'sd-0.12944773065115556, 32'sd0.02544672056292102, 32'sd0.03189616636990819, 32'sd0.12021853202331755, 32'sd-0.06130550570352322, 32'sd-0.14275415002044642, 32'sd-0.1601634620017828, 32'sd0.005092610464783461, 32'sd-0.024399954005055086, 32'sd-0.0031637045914405656, 32'sd0.06959629686988919, 32'sd0.08068974143632918, 32'sd-0.009715929200944454, 32'sd0.06220511891185563, 32'sd-0.085697372663246, 32'sd0.012868859573947374, 32'sd-0.013136735865831292, 32'sd-0.010931603225520942, 32'sd0.055605273201693256, 32'sd0.10544568643730491, 32'sd0.07021756178385781, 32'sd-0.07017792772420632, 32'sd0.05527757750702358, 32'sd0.00396624399362676, 32'sd0.012633305086003141, 32'sd-0.08938288737146943, 32'sd0.028474724948892364, 32'sd0.03704325422065581, 32'sd0.020129685566823652, 32'sd0.00027511941642470553, 32'sd0.12112738598061591, 32'sd-0.01880725392275845, 32'sd-0.08615516931303371, 32'sd-0.07806382141915004, 32'sd-0.09247511806784454, 32'sd-0.02268369427906742, 32'sd0.027063137625697252, 32'sd-0.05339051192462883, 32'sd0.0038871468846007925, 32'sd0.08998590212119187, 32'sd0.09334577983580211, 32'sd-0.06415900446653297, 32'sd0.0400912386154252, 32'sd0.0642809087767291, 32'sd0.0035206762321685786, 32'sd0.09081044772725196, 32'sd-0.06384187524091522, 32'sd0.05918734665326347, 32'sd0.026485665217331034, 32'sd-0.024440590708596235, 32'sd-0.0969064377490957, 32'sd-0.0699966770062687, 32'sd-0.06037244621378468, 32'sd-0.06681769946628924, 32'sd0.08749109248585624, 32'sd-0.0351377578879075, 32'sd-0.024588782393707997, 32'sd-0.06526468821085758, 32'sd0.04152534514107821, 32'sd-0.07785927420605668, 32'sd-0.03168278537797879, 32'sd0.12003994305296106, 32'sd0.01906165850103962, 32'sd0.010716425246721003, 32'sd0.11154848704850882, 32'sd0.05296731368749152, 32'sd0.05354010038783832, 32'sd0.11477684321115214, 32'sd-0.0719386999281314, 32'sd-0.02663558883738547, 32'sd0.09896622925799309, 32'sd0.10153242021167266, 32'sd0.038678409651519356, 32'sd0.0211254231676079, 32'sd0.05931951433895621, 32'sd-0.016941397635569864, 32'sd0.009777401565505283, 32'sd0.014756206559785537, 32'sd-0.10987886592805926, 32'sd-0.05253673682604727, 32'sd-0.09847280896329878, 32'sd0.008758470413216233, 32'sd0.04366477636037609, 32'sd-0.0075343274255441055, 32'sd-0.04083211288906754, 32'sd0.014355001100712146, 32'sd0.009363947682588676, 32'sd0.07643795613644122, 32'sd0.23087501980614417, 32'sd0.024829620854648685, 32'sd0.0916507380007836, 32'sd-0.0057634734013620355, 32'sd0.058521135988872854, 32'sd0.01923785427992546, 32'sd0.016734346239373227, 32'sd0.05856472368834852, 32'sd0.06459288158569504, 32'sd0.02887991235418394, 32'sd-0.12390929143386145, 32'sd-0.07776415265662599, 32'sd-0.005674537644872946, 32'sd0.09215497964787538, 32'sd-0.04012102830462114, 32'sd-0.03001059123618009, 32'sd0.016531356433755487, 32'sd0.043921966042403025, 32'sd0.024078589635330286, 32'sd-0.012979116494296977, 32'sd0.020192693664635167, 32'sd-0.1275849910281675, 32'sd-0.04030931325796083, 32'sd0.024352159383635955, 32'sd0.048952451855553275, 32'sd-0.02656137175248659, 32'sd0.16672268229181073, 32'sd0.16636362344276973, 32'sd0.1256841108594014, 32'sd0.13911682228031955, 32'sd-0.010414636046707731, 32'sd-0.0255914481386219, 32'sd-0.04545451584478587, 32'sd-0.014969647395557761, 32'sd0.09748814596562742, 32'sd-0.02691366774951058, 32'sd0.06330511796280161, 32'sd-0.06315187579503878, 32'sd-0.03721793166892084, 32'sd0.028796505356114412, 32'sd-0.037530678357628126, 32'sd0.09194295618951141, 32'sd0.09396095569464796, 32'sd-0.04437297895416538, 32'sd-0.010299800272706928, 32'sd0.1273554682016868, 32'sd0.026468511814248828, 32'sd0.06267834599793354, 32'sd-0.0809569772733799, 32'sd0.021418535165484854, 32'sd0.038287942508845915, 32'sd0.07091128512390446, 32'sd0.14635356216918569, 32'sd0.14662128553176504, 32'sd0.11264135788148717, 32'sd0.09576301401189498, 32'sd0.13638526921284846, 32'sd-0.017635770996206845, 32'sd-0.08160435067858239, 32'sd-0.01703165734493616, 32'sd0.010359970515318966, 32'sd-0.012037737305095303, 32'sd0.034658184776758805, 32'sd0.01835921107031988, 32'sd0.018814941585470174, 32'sd0.06371198995260142, 32'sd0.06335729197769666, 32'sd-0.014951737797056663, 32'sd0.017963650477281948, 32'sd-0.02033616413067889, 32'sd0.0028009589550432733, 32'sd0.01777274755796888, 32'sd0.06778007923538906, 32'sd-0.03362060066821327, 32'sd0.05235661189079831, 32'sd-0.006293612979173293, 32'sd-0.03536303663970448, 32'sd-0.00853303292794106, 32'sd0.06774682853065814, 32'sd0.07036250899958887, 32'sd0.1766421525777784, 32'sd0.0956380126759839, 32'sd-0.004441879421005704, 32'sd-0.08184735603381256, 32'sd0.05716947595931025, 32'sd0.03509200281696349, 32'sd0.05496266458151502, 32'sd-0.02800493869907827, 32'sd-0.0024821166657081786, 32'sd0.009773627788963991, 32'sd0.040067864215863364, 32'sd0.052904050873509106, 32'sd-0.07859539195438008, 32'sd0.04388408915425091, 32'sd0.06444862259752562, 32'sd0.015343876041908719, 32'sd0.024892127494021244, 32'sd0.02873201649788522, 32'sd0.06745206503864566, 32'sd-0.041727353431016516, 32'sd-0.03725569288364928, 32'sd-0.026083210011999303, 32'sd0.010124967939641983, 32'sd0.048899066101090724, 32'sd-0.0823776981378142, 32'sd-0.009327807120136212, 32'sd0.013681187625282299, 32'sd-0.06011474636704405, 32'sd-0.022981742717471516, 32'sd-0.09814040330713523, 32'sd-0.135242733096199, 32'sd-0.18302308174194806, 32'sd0.012758081639544155, 32'sd0.0025366107511502504, 32'sd-0.029414250231982318, 32'sd-0.08798684184429176, 32'sd0.03639926045104329, 32'sd0.007472655248047935, 32'sd0.004447447197803317, 32'sd0.0009333309373681409, 32'sd-0.028569131891343785, 32'sd-0.013954173170684528, 32'sd-0.03681313637227658, 32'sd-0.07725927808356284, 32'sd2.6966910733918535e-119, 32'sd-0.01920176942295423, 32'sd0.02039827319207355, 32'sd-0.017637437785652705, 32'sd-0.051334249138509265, 32'sd-0.09926680880683558, 32'sd-0.13955449090030353, 32'sd0.019865729126524186, 32'sd-0.17834668609614113, 32'sd-0.07983170762974792, 32'sd-0.12820354022129973, 32'sd-0.13561331788076902, 32'sd-0.19272015743891727, 32'sd-0.012578097486645344, 32'sd-0.010728861337912133, 32'sd-0.11958525583018874, 32'sd-0.12558308402817372, 32'sd0.004455312267369483, 32'sd0.07041887447441822, 32'sd0.049508442549787, 32'sd0.06926231043633495, 32'sd0.11008648955773294, 32'sd-0.05756361061450237, 32'sd0.031316994275772315, 32'sd0.024534818477016926, 32'sd0.05260577426947494, 32'sd-0.061606413596681155, 32'sd0.01003100177267718, 32'sd0.0020177749535067765, 32'sd0.03259923741624409, 32'sd-0.006044486957478466, 32'sd-0.09365683577532279, 32'sd-0.0436678871938688, 32'sd-0.10227869723293889, 32'sd-0.06909090769061353, 32'sd-0.030908170713862097, 32'sd-0.030894110216094554, 32'sd-0.08301683358764184, 32'sd-0.2245696061086488, 32'sd-0.20197133000213066, 32'sd-0.21657939193982736, 32'sd-0.12822966282730952, 32'sd0.07185592246680464, 32'sd-0.05845403043654569, 32'sd-0.012144696316566724, 32'sd0.0330911944340048, 32'sd-0.05294917883219984, 32'sd-0.004783256411228716, 32'sd-0.010861089900919154, 32'sd-0.018247881567862344, 32'sd-0.06923853127999714, 32'sd-0.1383404188789655, 32'sd-0.0771837621669836, 32'sd0.041961013429027, 32'sd0.1233883546273772, 32'sd0.0033158962116731304, 32'sd0.02896959723142891, 32'sd0.04107395445978675, 32'sd0.020682138254780106, 32'sd-0.07672027749210364, 32'sd-0.12163987566234136, 32'sd-0.05686507532328867, 32'sd-0.04878361833793668, 32'sd-0.10994753438312828, 32'sd-0.02922279097922159, 32'sd-0.07760170951870113, 32'sd-0.06018630013150097, 32'sd-0.18605328504829513, 32'sd-0.09773389679739217, 32'sd-0.039600563427111164, 32'sd-0.004424083645655625, 32'sd-0.035922130986558345, 32'sd-0.11089023883926709, 32'sd-0.09278652503513027, 32'sd0.1110314407998378, 32'sd0.0426050896734652, 32'sd-0.02127755181174438, 32'sd-0.011499130366040885, 32'sd-0.05172566242528335, 32'sd-0.08556838935813961, 32'sd0.0027779039468102495, 32'sd0.05945798017761562, 32'sd-0.01304786076375951, 32'sd0.07763178352103436, 32'sd-8.63022270839524e-117, 32'sd0.016021296937048003, 32'sd0.027630040799242524, 32'sd-0.03236687202407663, 32'sd-0.04057063558764523, 32'sd0.016374166423561504, 32'sd-0.019136117201890585, 32'sd-0.05757824125865207, 32'sd-0.02085475432668004, 32'sd0.029697209920105588, 32'sd0.02018781379446456, 32'sd0.034780826789720394, 32'sd0.03819233920599021, 32'sd0.07489262249221779, 32'sd0.03714913364610568, 32'sd-0.16624336568942807, 32'sd-0.1527924695592863, 32'sd0.031856854265906454, 32'sd-0.03248611713362379, 32'sd-0.027160833370531923, 32'sd-0.025160981075720186, 32'sd0.03258244843885117, 32'sd-0.028938181636690444, 32'sd-0.03340078552891361, 32'sd0.046982461218715035, 32'sd-0.05194356368991839, 32'sd0.10314489431336675, 32'sd0.04532563534684803, 32'sd0.049964760249711644, 32'sd0.01652612268402011, 32'sd0.0600021497094355, 32'sd0.1358517520458424, 32'sd0.1334251656719831, 32'sd0.0542844917322168, 32'sd0.022364620670693686, 32'sd0.00883564397021991, 32'sd-0.05234137220623037, 32'sd0.019112349403043075, 32'sd0.13064267884801584, 32'sd0.0751434989146184, 32'sd0.08912643996131002, 32'sd0.020600697821665095, 32'sd-0.05581461842698109, 32'sd0.018049367571831836, 32'sd-0.0656200304421023, 32'sd-0.0711550429311502, 32'sd-0.022660371662751103, 32'sd-0.09154005777147436, 32'sd0.05890564821300669, 32'sd-0.06095989182673816, 32'sd-0.042502747840112126, 32'sd-0.07551889280288514, 32'sd-0.10360244506290699, 32'sd-0.011707139916980575, 32'sd0.07988423950470694, 32'sd0.020461625549320236, 32'sd0.07309833779911791, 32'sd0.0053909640766795315, 32'sd-0.0032403450076109526, 32'sd0.10537031345750898, 32'sd0.05468849468654896, 32'sd-0.04055100241650348, 32'sd0.10761170271383687, 32'sd-0.015088646329052437, 32'sd0.08434021548109441, 32'sd0.06769335276796509, 32'sd0.07382383989004968, 32'sd0.08798783784523355, 32'sd0.0813232895517562, 32'sd0.12750909143217454, 32'sd0.13793118281620967, 32'sd-0.026124792648714975, 32'sd-0.07287930842775316, 32'sd0.05263252054875788, 32'sd0.0688351143217866, 32'sd-0.05835963229079778, 32'sd-0.019970373580580656, 32'sd-0.09845774777902024, 32'sd-0.1869411959591064, 32'sd-0.01781010303050337, 32'sd-0.09430357159238136, 32'sd0.06778073718140615, 32'sd0.023763132092452195, 32'sd0.06629743525529828, 32'sd-1.3016006856864665e-124, 32'sd0.01802354304538098, 32'sd0.005602068772800611, 32'sd0.027989816429764874, 32'sd0.02870411140845815, 32'sd0.05420963564565671, 32'sd0.10348777456111179, 32'sd0.10308249250038806, 32'sd0.049685216016332745, 32'sd0.16395635019546537, 32'sd0.12945427293025405, 32'sd0.0026474487925091652, 32'sd-0.01898880524985663, 32'sd0.08972071480792196, 32'sd0.008283443109700995, 32'sd-0.061881893289687497, 32'sd0.02968751382359669, 32'sd0.03895167850950791, 32'sd0.09791589848283397, 32'sd-0.023982729537003353, 32'sd-0.00020541702270885707, 32'sd0.008987977189790757, 32'sd-0.03654458913945581, 32'sd0.010195580334105087, 32'sd-0.003415797909369518, 32'sd-0.06617833522807849, 32'sd-0.013024003638176112, 32'sd3.609351722299843e-116, 32'sd-1.9598589838752186e-117, 32'sd2.076389909603565e-117, 32'sd-0.031969609741152726, 32'sd0.08259774083511733, 32'sd0.05780049672937926, 32'sd0.025521263385842815, 32'sd-0.0142981393244737, 32'sd0.13929917615196266, 32'sd0.13126645018644922, 32'sd-0.022933790630920003, 32'sd0.04365041767352106, 32'sd-0.10206151407921857, 32'sd-0.02761263267446664, 32'sd0.04775140444754464, 32'sd-0.061220955011171016, 32'sd-0.06888166395624765, 32'sd-0.07900916549012647, 32'sd0.009397025210683436, 32'sd-0.009496354559110482, 32'sd-0.07662485619453605, 32'sd-0.04954142786240692, 32'sd-0.021417502593830316, 32'sd-0.02160286585793625, 32'sd-0.010457320657450088, 32'sd-0.025205953285584556, 32'sd-0.010283936458594892, 32'sd0.02441013535848292, 32'sd2.0905776161454046e-117, 32'sd5.822430467643609e-126, 32'sd-2.7920285692533394e-116, 32'sd0.06604997528375947, 32'sd-0.07466096835032761, 32'sd-0.03497953274826979, 32'sd0.1021140547996501, 32'sd-0.010282872222554675, 32'sd0.02673047980642802, 32'sd0.03248619914079396, 32'sd-0.08220146877864325, 32'sd-0.003419645504722621, 32'sd-0.01646462530917025, 32'sd-0.04678989271191215, 32'sd0.05819542988406973, 32'sd0.005476040579214769, 32'sd-0.015120917063468709, 32'sd-0.061227619252293454, 32'sd-0.0038489830030710107, 32'sd0.047310977953482755, 32'sd-0.0646406614470694, 32'sd-0.07891211122829563, 32'sd-0.0686856481482174, 32'sd-0.03631337783359555, 32'sd0.06215563010374875, 32'sd-0.014939982379022634, 32'sd0.06015802583989731, 32'sd0.025568468821506412, 32'sd-1.9411246766550117e-123, 32'sd-1.4312867682850058e-118, 32'sd-2.3484093729153248e-125, 32'sd-6.386320932792821e-117, 32'sd0.04117621892342671, 32'sd-0.03542912357248172, 32'sd-0.019322652904807076, 32'sd-0.00729422637034283, 32'sd0.0015036465295633927, 32'sd0.020301633977068093, 32'sd0.05712628678651124, 32'sd0.0492897978092563, 32'sd-0.0632214664938346, 32'sd-0.04445749359981658, 32'sd-0.009511984926159652, 32'sd-0.13013768486066915, 32'sd-0.027400453577965486, 32'sd0.05616561400565517, 32'sd0.07862051762384097, 32'sd0.00963098207744717, 32'sd0.05004449444553628, 32'sd-0.07594192327008663, 32'sd-0.011940592918125544, 32'sd-0.030379949885485206, 32'sd0.055446170883919774, 32'sd-0.0076141332876254585, 32'sd0.025509465307502165, 32'sd2.073230163171752e-126, 32'sd-3.354728843315941e-120, 32'sd6.893256403843519e-120, 32'sd3.307235580286653e-120, 32'sd-3.0602579529650993e-121, 32'sd4.3634384034647455e-128, 32'sd0.07215677176886195, 32'sd0.09325246332219515, 32'sd-0.0017309918181828295, 32'sd0.09011037531667643, 32'sd-0.0013720463960287378, 32'sd-0.04639097228479943, 32'sd0.0261139894464124, 32'sd0.0909351361992627, 32'sd0.031604652447136686, 32'sd0.021578967720356855, 32'sd-0.027688516205223047, 32'sd-0.06399961184112067, 32'sd-0.019406516467088582, 32'sd-0.012699208199282778, 32'sd0.0763153168509916, 32'sd0.03520831471054831, 32'sd0.02774770598000089, 32'sd-0.020719573051321185, 32'sd-0.021603180469688316, 32'sd0.02420302165450233, 32'sd7.152159638681702e-125, 32'sd1.0405806432273694e-120, 32'sd-1.4799565554185108e-124, 32'sd-1.0581635716070972e-119},
        '{32'sd-6.918966035447998e-115, 32'sd-1.8378315090572044e-116, 32'sd3.907366371320888e-124, 32'sd-6.944053304847761e-115, 32'sd-3.15353166705128e-124, 32'sd3.1521798416661185e-116, 32'sd3.1110900130993015e-122, 32'sd-5.884324253228559e-129, 32'sd2.679961835421944e-118, 32'sd1.8874345363398816e-117, 32'sd8.407271707924129e-122, 32'sd2.3948621641605215e-124, 32'sd0.0147727399594456, 32'sd0.0666591427259206, 32'sd0.0912022529894863, 32'sd0.07498793722816743, 32'sd-5.758971593471708e-121, 32'sd-7.305983888277439e-117, 32'sd2.114008786690929e-116, 32'sd2.150005308498399e-127, 32'sd-1.9455073809734786e-127, 32'sd-4.02407721377909e-129, 32'sd-1.733128463075431e-125, 32'sd-3.544275196994516e-124, 32'sd-1.498277444044281e-127, 32'sd-5.755126738380817e-128, 32'sd-1.5791537653670654e-117, 32'sd-2.444312600588478e-125, 32'sd-2.7117400281192538e-124, 32'sd7.452360028561115e-127, 32'sd2.406521380663943e-114, 32'sd8.348119646420476e-125, 32'sd-0.024566578968505025, 32'sd-0.011325307655389211, 32'sd-0.023208157070392, 32'sd0.0635297180641687, 32'sd0.007226586155027382, 32'sd-0.06554018972346298, 32'sd0.021514963118864572, 32'sd0.07859577279969453, 32'sd0.06035601565406585, 32'sd0.004102551106880829, 32'sd-0.011121790069391655, 32'sd0.01140780573156378, 32'sd0.05448323114269064, 32'sd-0.06436079056502286, 32'sd0.01759464620200035, 32'sd0.12329176237148157, 32'sd0.0010502542169791682, 32'sd0.09618487187756197, 32'sd0.08894133306429872, 32'sd0.047446364559151286, 32'sd-7.375360900603556e-127, 32'sd-2.997447845039547e-115, 32'sd1.8244423868551381e-124, 32'sd-3.96343232563445e-118, 32'sd-1.5124367356878907e-115, 32'sd-2.710031943365495e-114, 32'sd0.07826559836145439, 32'sd0.02037463517461603, 32'sd0.05686043397236619, 32'sd0.08457144592372336, 32'sd0.09397579907610626, 32'sd0.04109978982282005, 32'sd0.011262484627706407, 32'sd0.04218363143842316, 32'sd0.046006670923603325, 32'sd0.09698875580498417, 32'sd0.0324290678371029, 32'sd0.052959959840332985, 32'sd0.09451405088722994, 32'sd-0.04085173299213526, 32'sd-0.06788132553844939, 32'sd0.2632519978889562, 32'sd0.14315974991828756, 32'sd0.05016717072693093, 32'sd-0.06530617063264049, 32'sd0.07885702223054025, 32'sd0.13573817644491468, 32'sd0.15691084866535043, 32'sd-0.027668656591106094, 32'sd0.09899489961578618, 32'sd-5.581894731741659e-121, 32'sd3.696044281777464e-125, 32'sd-2.1735691476588106e-116, 32'sd-1.9060441793906803e-128, 32'sd0.04673865577509815, 32'sd0.007223679798554418, 32'sd-0.02616099571124953, 32'sd0.09843229052071022, 32'sd-0.018217320444150475, 32'sd-0.07717854500641895, 32'sd0.11270786705781308, 32'sd0.06522511348618916, 32'sd0.048981273029134166, 32'sd-0.10466606195581064, 32'sd0.0009746788450805645, 32'sd-0.12794641504301843, 32'sd-0.0039276316719152925, 32'sd0.1799416841780363, 32'sd0.04598751952063366, 32'sd0.015016836409355768, 32'sd0.09033934422357218, 32'sd0.07055382680557701, 32'sd0.027076348651049305, 32'sd0.07765533353421826, 32'sd0.03588411940259469, 32'sd0.02748776307379601, 32'sd0.0647082015957121, 32'sd-0.046650867538146006, 32'sd0.06830976372539194, 32'sd3.2157101279024714e-119, 32'sd-3.3532418199167676e-121, 32'sd0.013689204040303694, 32'sd0.029723313905146057, 32'sd-0.08026424792063411, 32'sd-0.07164031677316451, 32'sd-0.08140329030109486, 32'sd-0.04215162852088256, 32'sd-0.1972579201498312, 32'sd-0.07308550799555037, 32'sd-0.021338349855352, 32'sd-0.004294116947673651, 32'sd0.0334754492123434, 32'sd-0.04517556768395173, 32'sd-0.05568547556596783, 32'sd-0.06714010851858379, 32'sd-0.037800225609161534, 32'sd0.056567052766888136, 32'sd0.09922560551695316, 32'sd-0.03335961700893997, 32'sd0.0610482050680288, 32'sd0.01737892621784217, 32'sd0.04362926658372602, 32'sd-0.08321497503989454, 32'sd0.06995764881730293, 32'sd0.006739080597744233, 32'sd-0.007939361566755817, 32'sd-0.01314739492432812, 32'sd-0.010404153201530186, 32'sd6.318505432102952e-126, 32'sd0.004702429969979997, 32'sd-0.03253811316513569, 32'sd0.099800821487899, 32'sd-0.03488614408665371, 32'sd-0.08219207982793011, 32'sd-0.04018804340535368, 32'sd-0.08619876394483476, 32'sd-0.03571085440039482, 32'sd-0.08244628205672153, 32'sd-0.024013181854522933, 32'sd-0.12124536795617115, 32'sd0.023232722665857596, 32'sd-0.041836854737080084, 32'sd-0.02192931749701411, 32'sd-0.0658555678806316, 32'sd0.08806232704603065, 32'sd0.14678759019229679, 32'sd0.06813720882025551, 32'sd0.03981129961945354, 32'sd0.12033613328478843, 32'sd0.03040668269038952, 32'sd0.028527862076652363, 32'sd0.09441932006841629, 32'sd0.1246437487331419, 32'sd0.010049716820861055, 32'sd-0.011450745419537821, 32'sd0.02150206178842989, 32'sd4.524830204204394e-121, 32'sd0.05187925912874503, 32'sd0.031334989868160204, 32'sd0.13475366709530387, 32'sd0.010555377779972593, 32'sd0.04884214741998038, 32'sd-0.0005672053042147651, 32'sd0.09021647393026529, 32'sd-0.02524796330147114, 32'sd-0.01874656161851507, 32'sd-0.021485526565875365, 32'sd0.024691026168667172, 32'sd0.10378866916584864, 32'sd0.03695647433599746, 32'sd0.057407790611394616, 32'sd0.051388019236594605, 32'sd0.061911769956971036, 32'sd-0.06307450314627977, 32'sd0.0030935406591609533, 32'sd0.11295096663886157, 32'sd-0.06748682048326753, 32'sd-0.11115634403841636, 32'sd-0.01416793901498248, 32'sd0.11268258928396795, 32'sd0.06371805282474478, 32'sd0.011384796405318464, 32'sd0.026252912986627852, 32'sd0.11024151115200044, 32'sd0.07755225011793339, 32'sd0.03445403606313923, 32'sd-0.03502979387952057, 32'sd-0.07405289042133563, 32'sd0.011893323184583571, 32'sd-0.03738691012586967, 32'sd0.100466422624606, 32'sd-0.002924103949681299, 32'sd0.022805631703708272, 32'sd-0.09899731235992139, 32'sd-0.016864727790656377, 32'sd-0.018371637447952897, 32'sd0.04942110975355909, 32'sd0.04902846030838115, 32'sd0.006387362059140722, 32'sd-0.0788013089753786, 32'sd-0.10955983727451817, 32'sd-0.10709390971162526, 32'sd0.015153903257061379, 32'sd-0.17472224057869926, 32'sd-0.09985956162752604, 32'sd-0.28061090471295125, 32'sd-0.22562740415027835, 32'sd-0.08784954981750298, 32'sd-0.027792577917400866, 32'sd-0.014871768981150538, 32'sd-0.11236890197131169, 32'sd-0.0646138418220925, 32'sd0.013639709178433646, 32'sd0.01196592515834811, 32'sd-0.16502018717939068, 32'sd-0.19194430374227922, 32'sd-0.10811977403876814, 32'sd-0.0873967809447918, 32'sd0.044045981749223896, 32'sd0.009232904516286486, 32'sd0.09442772984923872, 32'sd-0.05911947978950835, 32'sd0.032158094762560374, 32'sd0.12305880130844651, 32'sd-0.004002883374871775, 32'sd-0.00015554389363682446, 32'sd-0.025151490014364, 32'sd-0.19715925315884655, 32'sd-0.12240196104084915, 32'sd-0.10037438830131731, 32'sd-0.26036753816308195, 32'sd-0.2549468637891234, 32'sd-0.24035874693231102, 32'sd-0.30519465368647264, 32'sd-0.3101569610902757, 32'sd-0.1564489214589816, 32'sd-0.14534148934055863, 32'sd-0.14750106601538518, 32'sd-0.07313783633883272, 32'sd0.06448299820811257, 32'sd0.03411028754096227, 32'sd-0.07342354074702752, 32'sd0.014308162335376995, 32'sd-0.047076359981189184, 32'sd-0.09211869605783847, 32'sd-0.008095650384968357, 32'sd-0.08286612743172873, 32'sd0.06396278431302933, 32'sd0.027342534766656056, 32'sd0.06346247589568178, 32'sd-0.013561323410726862, 32'sd-0.04708981672746817, 32'sd0.0890864643114677, 32'sd-0.11175279610714052, 32'sd-0.10880468748426934, 32'sd-0.09497804076735344, 32'sd-0.25057386826036077, 32'sd-0.14868891875270795, 32'sd-0.22320026516481178, 32'sd-0.20840411093752634, 32'sd-0.15626853341851762, 32'sd-0.1332019367945063, 32'sd-0.10019411540053101, 32'sd-0.08741210325121213, 32'sd0.03735441923330027, 32'sd-0.07846652750049571, 32'sd0.07384204522600846, 32'sd-0.04781348738274109, 32'sd-0.023675460667686027, 32'sd0.047555313801556316, 32'sd-0.05820530411273295, 32'sd0.02573688498949188, 32'sd0.04530872727229653, 32'sd0.08933830685526692, 32'sd0.11457833216820949, 32'sd0.06764763997382428, 32'sd-0.00483093345251556, 32'sd-0.02853067625688896, 32'sd-0.03982522192095271, 32'sd0.011199737072917498, 32'sd0.003150304810624445, 32'sd-0.11150586082046218, 32'sd-0.14098443278628794, 32'sd-0.16859504060748812, 32'sd-0.17171139872954028, 32'sd-0.012613970264769092, 32'sd-0.03577975738732305, 32'sd-0.0897305723918594, 32'sd-0.08085897390191435, 32'sd-0.09084808588349923, 32'sd-0.12665922862589413, 32'sd0.05922697297075176, 32'sd0.11868339391418621, 32'sd0.049279455326683694, 32'sd-0.05132700675924988, 32'sd-0.08998901579838035, 32'sd0.025807863677293243, 32'sd0.009924633609235511, 32'sd-0.02435953711031974, 32'sd-0.11377940371699329, 32'sd-0.06407341815529531, 32'sd-0.07267382592995489, 32'sd0.05674395069887074, 32'sd-0.016868419412221104, 32'sd0.08570869490993069, 32'sd-0.10267845691563207, 32'sd0.014114228744218913, 32'sd0.08561362593361677, 32'sd0.016918491830270378, 32'sd-0.039058039424004404, 32'sd0.04903827916156811, 32'sd-0.08801229122759228, 32'sd0.01340838496819618, 32'sd-0.0916536266712377, 32'sd-0.036571699482879534, 32'sd0.07801301419997356, 32'sd0.005252412741390663, 32'sd-0.03263174494214362, 32'sd-0.0031512579310215057, 32'sd0.18139077501821693, 32'sd0.11992699626674434, 32'sd0.06551790036318768, 32'sd-0.011982458810990007, 32'sd0.023557736119272928, 32'sd0.06324141346163326, 32'sd0.018437712712654094, 32'sd-0.024998091503296644, 32'sd-0.007046106575946222, 32'sd-0.07747913497771315, 32'sd-0.08064668509826435, 32'sd-0.06557977967224106, 32'sd0.0609594695572429, 32'sd-0.044623499859351594, 32'sd0.03921199786975338, 32'sd0.006239597242360536, 32'sd0.09643903092410153, 32'sd-0.024350787154470366, 32'sd0.12695602217656263, 32'sd0.1611716169482534, 32'sd-0.011037429144382946, 32'sd0.0021392953025171197, 32'sd-0.03615551661600219, 32'sd-0.08577162441847686, 32'sd-0.006440220356238746, 32'sd-0.05340459318545418, 32'sd-0.03976235972578375, 32'sd0.14637680928052338, 32'sd0.007642721893609484, 32'sd0.007809830298127056, 32'sd-0.029778019490820585, 32'sd-0.04246493673948882, 32'sd-0.029589445292573516, 32'sd0.029288259910042136, 32'sd0.04019278680257097, 32'sd-0.09271114333513802, 32'sd-0.037044934383682206, 32'sd-0.1985246582652107, 32'sd-0.0684790334714664, 32'sd-0.0944812694961435, 32'sd0.03660052037160486, 32'sd0.07785268458768366, 32'sd0.06144880260783731, 32'sd-0.04675490603641234, 32'sd-0.04410986904490677, 32'sd-0.013342005721070546, 32'sd0.1463942454437622, 32'sd0.18487381089363103, 32'sd0.11916217449484379, 32'sd0.09078626961425607, 32'sd0.05322802155969025, 32'sd0.05444183323364678, 32'sd0.06335808704297743, 32'sd-0.03610202794751165, 32'sd-0.07463254077275916, 32'sd-0.035399218239182934, 32'sd-0.01014078591370288, 32'sd-0.006809168659431075, 32'sd-0.07107531363155717, 32'sd-0.0007803491072869108, 32'sd-0.05139690511154692, 32'sd0.014545451714850392, 32'sd-0.025428901094704272, 32'sd0.01696493806807748, 32'sd-0.022841826693328505, 32'sd-0.03709383285038025, 32'sd-0.0849974677848479, 32'sd-0.02080585201847254, 32'sd0.04584335268245547, 32'sd-0.07567019943435677, 32'sd-0.006692735876515707, 32'sd0.11842290752668319, 32'sd0.0194442073918741, 32'sd-0.037415573415569704, 32'sd0.1115935252453972, 32'sd0.1188981475503667, 32'sd0.12608261959212042, 32'sd0.21611556692043174, 32'sd0.08170367235722337, 32'sd0.11405182353247205, 32'sd0.08581102944862018, 32'sd-0.05513067015221997, 32'sd-0.0499607246179168, 32'sd-0.01424082509165081, 32'sd-0.07922474247850318, 32'sd-0.11915523730673727, 32'sd0.050845611978335585, 32'sd-0.0028089642413353373, 32'sd-0.005050006764764639, 32'sd0.00027579927346394037, 32'sd-0.04978905518176387, 32'sd-0.04897434386560564, 32'sd-0.003732844350994, 32'sd0.022057125464577425, 32'sd-0.054877901418787206, 32'sd0.09687439898076314, 32'sd-0.07844490895277562, 32'sd-0.035518309742987204, 32'sd-0.10485994282963748, 32'sd-0.02598143521205868, 32'sd0.05011385402621348, 32'sd0.09917853991337691, 32'sd0.08604532636327004, 32'sd0.08329376287191795, 32'sd0.10218610592291302, 32'sd0.20238441568203375, 32'sd0.11459334292760598, 32'sd0.11659115541758593, 32'sd0.144027228768408, 32'sd-0.02506559308479352, 32'sd0.09755993789734851, 32'sd-0.0024897599451524093, 32'sd-0.004621555840212071, 32'sd0.09358253320168698, 32'sd-0.01076776375287303, 32'sd-0.10059635888216126, 32'sd-0.052996323418221684, 32'sd0.017745083773636317, 32'sd0.03157764028385914, 32'sd-0.060307697860592174, 32'sd-0.06628687877838255, 32'sd-0.0943643133979758, 32'sd-0.1298342386063965, 32'sd-0.018551677599601916, 32'sd-0.09954260614921415, 32'sd-0.1331887867319902, 32'sd-0.08921203901768297, 32'sd0.06748931141599437, 32'sd0.021034282910431336, 32'sd-0.002189889133749366, 32'sd-0.023210614895661216, 32'sd-0.025897339322672956, 32'sd0.04419609006967639, 32'sd0.011149803155045148, 32'sd0.23223138559890555, 32'sd0.06400914555321233, 32'sd0.08538923754325406, 32'sd0.10252942110334161, 32'sd0.15096742784012288, 32'sd0.13560628190894278, 32'sd0.17101688538465, 32'sd0.11208388045134779, 32'sd-0.000489898896504607, 32'sd0.0641818565981785, 32'sd0.05144736085088446, 32'sd-5.5441491808728455e-118, 32'sd0.03783310691883226, 32'sd-0.009613055128337222, 32'sd0.06101748252652768, 32'sd-0.022900646784986198, 32'sd-0.038756146932917096, 32'sd0.05453395419232856, 32'sd-0.04457378658050499, 32'sd0.019120243748515085, 32'sd-0.010201273460523944, 32'sd0.02069178277045704, 32'sd-0.03825100282050938, 32'sd0.007472077441238331, 32'sd-0.08686074170784715, 32'sd-0.12012702301040434, 32'sd-0.0831534978686, 32'sd0.08359180034950141, 32'sd0.15636076913093439, 32'sd0.1092164818746941, 32'sd-0.009395998380260564, 32'sd0.11369353702929365, 32'sd0.16879865534041705, 32'sd0.09469061729480187, 32'sd-0.025503864840519478, 32'sd0.00044275864797571954, 32'sd-0.051236050076623595, 32'sd0.0020092038026060803, 32'sd0.05336127950171922, 32'sd-0.0012575298423220481, 32'sd0.010443667856098444, 32'sd0.09911794845422169, 32'sd-0.022375097497362745, 32'sd-0.042535910190635726, 32'sd0.02979564217003809, 32'sd-0.029551697820716705, 32'sd0.008944845089490611, 32'sd0.05983453113267737, 32'sd0.028026302186421305, 32'sd-0.03440322457038332, 32'sd-0.023693267717704858, 32'sd-0.06224755937318001, 32'sd0.00885563311437782, 32'sd0.04633694839420502, 32'sd-0.06707736809254486, 32'sd-0.006317371050676853, 32'sd0.10884614697928617, 32'sd0.08423493176862923, 32'sd0.14389505951981701, 32'sd0.11937039327425411, 32'sd0.12797426780848042, 32'sd0.09074199684411711, 32'sd0.045893030987376675, 32'sd-0.03548228575859409, 32'sd0.0697344427230585, 32'sd0.053364258057406744, 32'sd0.0083683267390705, 32'sd0.015844669027278043, 32'sd-0.09511172664706902, 32'sd0.11817770633886228, 32'sd-0.07397951558060499, 32'sd-0.043694647478329886, 32'sd-0.043555370426653084, 32'sd-0.12520906436908, 32'sd0.0031876460118190424, 32'sd0.0688883143133051, 32'sd0.03483517242605912, 32'sd0.00815774113266575, 32'sd0.0629431297119156, 32'sd-0.06065557818203473, 32'sd-0.06031029674059078, 32'sd0.060412584028806136, 32'sd-0.09400760860306037, 32'sd0.029583989728726515, 32'sd0.08512822487112233, 32'sd0.032959690571240416, 32'sd0.019581893608230014, 32'sd0.057662268545660415, 32'sd-0.0062255937751427475, 32'sd0.026457703605660285, 32'sd0.1325455428002976, 32'sd-0.039369587587939396, 32'sd0.10078021754911902, 32'sd0.0004934740706944328, 32'sd0.07878666227487127, 32'sd4.373816741767108e-127, 32'sd-0.006546573099360819, 32'sd0.033223132631551536, 32'sd-0.04629750637322829, 32'sd0.024351755249551302, 32'sd0.009806575563439265, 32'sd-0.011263019049448993, 32'sd-0.029416401375806055, 32'sd-0.03696757833182964, 32'sd0.06512368969907086, 32'sd0.027496665566881646, 32'sd0.0306330376468471, 32'sd-0.03995935235633798, 32'sd0.04588947948908815, 32'sd-0.021633168051411727, 32'sd-0.02552525265367142, 32'sd-0.048408771741243584, 32'sd0.039830884406048976, 32'sd-0.020462109708174605, 32'sd0.11957088657887956, 32'sd0.1108014214505435, 32'sd0.1093725046479096, 32'sd0.12351002398769059, 32'sd0.0060787985110372965, 32'sd-0.038506406320692146, 32'sd0.03277362987867337, 32'sd-0.04172685781366554, 32'sd0.026900522975754848, 32'sd0.028894383556064315, 32'sd-0.06152276713885309, 32'sd-0.05185876222848538, 32'sd-0.09807921976481014, 32'sd-0.009554744922987338, 32'sd0.06467079624630394, 32'sd0.03145877421360855, 32'sd0.059740212849834246, 32'sd-0.0028428854307516772, 32'sd0.037771264918932304, 32'sd0.01706931946267158, 32'sd-0.03208573391063834, 32'sd0.08629745150758253, 32'sd-0.023537754142094636, 32'sd0.0014866005659198553, 32'sd-0.0593459178449964, 32'sd-0.06960448428297568, 32'sd-0.1058673537650215, 32'sd-0.049965263971601684, 32'sd0.11633418835650247, 32'sd0.14641468710087271, 32'sd0.0021206865233682573, 32'sd0.06547295731240307, 32'sd0.06655113138601362, 32'sd-0.09351990424697314, 32'sd-0.00015862011652645054, 32'sd0.04048291757583582, 32'sd0.03417859134632975, 32'sd0.031115181208867162, 32'sd0.05884517115488653, 32'sd0.026038887764651783, 32'sd0.00898621930561767, 32'sd-0.042188685595547164, 32'sd0.03327468113521261, 32'sd0.07643687137769972, 32'sd0.11975766757790601, 32'sd-0.00877440246934862, 32'sd0.08537171039244353, 32'sd0.053605314165001784, 32'sd0.04418439334627972, 32'sd-0.04458668050407981, 32'sd-0.059964047171560175, 32'sd-0.105408281216178, 32'sd-0.10362057706609179, 32'sd-0.182692503656182, 32'sd-0.15223736079323416, 32'sd-0.12483218078506066, 32'sd0.008874906568644108, 32'sd-0.03160837098440288, 32'sd0.00804696827308926, 32'sd0.016551686372499534, 32'sd-0.04426766516578098, 32'sd-0.05460027281342034, 32'sd-0.025588374658713078, 32'sd-0.03779178393731754, 32'sd0.010765018868556667, 32'sd1.329735624871677e-122, 32'sd0.04049967838445972, 32'sd0.017670758524882948, 32'sd-0.02519833771862671, 32'sd0.03534944761198037, 32'sd0.053117722319360336, 32'sd0.034079368125232844, 32'sd0.006965666411478971, 32'sd0.004657788593694559, 32'sd0.04504829577279735, 32'sd0.06946093663084361, 32'sd-0.01982890462305264, 32'sd-0.007238920713907144, 32'sd0.05641992579328293, 32'sd-0.14940499410881625, 32'sd-0.16867953771252675, 32'sd-0.11320582808083798, 32'sd-0.13188056985890567, 32'sd-0.2062883385913878, 32'sd-0.10805434008906722, 32'sd-0.08566959777674077, 32'sd-0.09848336105652374, 32'sd-0.0008123920521811696, 32'sd-0.17821899179308165, 32'sd0.02157174631130677, 32'sd0.03574900286226731, 32'sd-0.1176201260984867, 32'sd1.589159571471902e-117, 32'sd-2.8743266593475415e-116, 32'sd-6.693017257396632e-117, 32'sd-0.007914621662858619, 32'sd0.046154925908892384, 32'sd0.01634341402201367, 32'sd-0.014465545689015683, 32'sd-0.0054117318965723644, 32'sd0.04069009498333224, 32'sd-0.018279485383901076, 32'sd-0.09550527953966886, 32'sd-0.13286653298150364, 32'sd-0.09867073398236317, 32'sd-0.06856515425896692, 32'sd-0.018049378184205222, 32'sd-0.07379640526235792, 32'sd-0.04388147387328128, 32'sd-0.04219631166633167, 32'sd-0.11010356304380037, 32'sd-0.09675353205276042, 32'sd-0.17689585574270622, 32'sd-0.09285628533728657, 32'sd-0.014453375441838645, 32'sd0.024779071184708706, 32'sd-0.18706874177145522, 32'sd-0.02126906922828956, 32'sd0.06637327651857529, 32'sd0.048108801249528974, 32'sd1.4185498716850059e-127, 32'sd3.957572057931639e-116, 32'sd2.2115733079064242e-119, 32'sd0.013716894887006592, 32'sd0.05961539886076337, 32'sd-0.049029754211750806, 32'sd0.05316025864354813, 32'sd0.0027114716648788304, 32'sd-0.0495684793922966, 32'sd-0.07761744331017088, 32'sd0.10151342733131183, 32'sd-0.061792524502183296, 32'sd0.022213985060673645, 32'sd-0.009910493013342308, 32'sd-0.047822436500912675, 32'sd-0.015186097458265031, 32'sd0.08675047859592563, 32'sd0.11947970554380281, 32'sd-0.19011781961803403, 32'sd-0.10843871566822125, 32'sd-0.06918903887973589, 32'sd-0.0861844471232264, 32'sd-0.023932896191376313, 32'sd-0.10556983960248097, 32'sd-0.13720173297830893, 32'sd-0.05738303378158762, 32'sd0.027664683940401835, 32'sd-0.029748304122597612, 32'sd2.7329597742919267e-116, 32'sd1.6253039413062978e-115, 32'sd2.684138433233128e-119, 32'sd-1.2213191532521612e-118, 32'sd0.06484245281135749, 32'sd0.07833824677993342, 32'sd0.035669920532121036, 32'sd-0.00026244928112674113, 32'sd0.00292111377007904, 32'sd-0.052173777141705194, 32'sd0.053084807331676816, 32'sd-0.06632837079120103, 32'sd-0.07100765641312282, 32'sd0.09864915063727368, 32'sd0.05030500427177719, 32'sd0.12285576790026659, 32'sd-0.09842584223642913, 32'sd0.016946602800710146, 32'sd0.042080958199920374, 32'sd-0.050570766448799175, 32'sd-0.017413193305741675, 32'sd0.09177450920997232, 32'sd-0.012777981567752032, 32'sd0.023065146231617897, 32'sd-0.0577027918637151, 32'sd0.04110719922353432, 32'sd0.061049398996102726, 32'sd1.3393684488950626e-122, 32'sd9.445983996056385e-125, 32'sd1.7119314671100102e-122, 32'sd3.9099505735440673e-118, 32'sd-8.555450686206016e-119, 32'sd2.7355227640484566e-125, 32'sd0.07619195580090603, 32'sd0.05359359097110981, 32'sd0.046764842052725845, 32'sd-0.014772137055357005, 32'sd-0.008506606527672603, 32'sd0.049453314479649506, 32'sd0.024896372430258416, 32'sd0.08228885949758817, 32'sd0.06203749465596387, 32'sd0.07972712218594438, 32'sd0.03416809255810912, 32'sd-0.018042695110527123, 32'sd0.07958846246149541, 32'sd0.03880766019840791, 32'sd0.03434304126819887, 32'sd-0.03723401642123291, 32'sd0.023043029554306812, 32'sd-0.05090516586010707, 32'sd-0.051316394526446894, 32'sd0.041518038279159925, 32'sd-7.19574568508432e-115, 32'sd1.927021235783931e-121, 32'sd9.461751447970494e-126, 32'sd-3.092565963350739e-120},
        '{32'sd3.29232835998905e-123, 32'sd2.15479737012033e-127, 32'sd-2.4896314571761586e-116, 32'sd-2.972970949355999e-116, 32'sd3.848669205990335e-127, 32'sd1.415250495559326e-118, 32'sd-2.616454904237217e-125, 32'sd1.169888220873787e-116, 32'sd-2.1730761239497156e-119, 32'sd-3.8535243733009223e-119, 32'sd-1.4956121194119657e-126, 32'sd6.101383497897952e-121, 32'sd0.009011349027757817, 32'sd0.021117054083991862, 32'sd-0.0094264285467419, 32'sd0.0178066198541402, 32'sd2.6719659786185304e-120, 32'sd-3.488739938072159e-126, 32'sd9.108068978103719e-123, 32'sd5.4848702015267314e-123, 32'sd3.346973503890056e-114, 32'sd2.895942243683968e-116, 32'sd-6.141591702060094e-115, 32'sd-7.186333748630596e-118, 32'sd1.128411893562875e-125, 32'sd1.8799744620214712e-120, 32'sd-1.4359417203741432e-116, 32'sd3.712102649022245e-119, 32'sd6.464132475000709e-123, 32'sd-1.1389971263380594e-116, 32'sd-2.75107660627643e-119, 32'sd1.9749671294270245e-119, 32'sd0.03922656325088632, 32'sd0.01287548736953918, 32'sd0.044106126395271575, 32'sd0.05396632555766461, 32'sd0.036775947175931537, 32'sd0.04431292940194917, 32'sd0.06579912445612668, 32'sd0.047178390931581625, 32'sd0.11079325201984268, 32'sd0.09471697027313418, 32'sd0.01342399379112632, 32'sd0.085506798242656, 32'sd0.009207209652371361, 32'sd0.08791166813150131, 32'sd0.013944376110392738, 32'sd0.09347091516819354, 32'sd0.07476649860181032, 32'sd0.01635398358345191, 32'sd0.09281383400384134, 32'sd0.010326337919182247, 32'sd1.8340865492952006e-123, 32'sd-5.108900304550255e-118, 32'sd3.1026249419540116e-119, 32'sd-8.794995723315203e-127, 32'sd3.395808375409381e-120, 32'sd-1.0266451388030318e-121, 32'sd0.01796236858020632, 32'sd-0.026276241387395354, 32'sd0.014418766524876477, 32'sd0.019912994734004787, 32'sd0.017624641712050092, 32'sd-0.047675474450316904, 32'sd-0.011881315076016235, 32'sd-0.03277945306939692, 32'sd4.2596550224753506e-05, 32'sd0.18631782649959705, 32'sd-0.01525385876889325, 32'sd-0.011591274748069738, 32'sd0.09541925682983039, 32'sd0.03187441130884832, 32'sd-0.020253880377138628, 32'sd0.1717266647379927, 32'sd0.07014707952125192, 32'sd0.1859481760381541, 32'sd0.12117116203432693, 32'sd0.0761750062254329, 32'sd0.061004338210280416, 32'sd0.07060910375710754, 32'sd0.03803458550480682, 32'sd-0.0062471233405936724, 32'sd1.1402043226580418e-118, 32'sd2.591433855004067e-126, 32'sd-4.0209045079411775e-123, 32'sd2.2622281749460775e-120, 32'sd0.06101600046689864, 32'sd0.034575662036257955, 32'sd-0.006296225100555857, 32'sd-0.10325600708525973, 32'sd-0.04395128444520148, 32'sd-0.1293892008056253, 32'sd0.1169626905003403, 32'sd0.0728417927041973, 32'sd0.01472244446560199, 32'sd0.0866072358732956, 32'sd0.13963833437503856, 32'sd0.19309586241312882, 32'sd0.1013363299232891, 32'sd0.04798015397937835, 32'sd-0.029029676913156804, 32'sd0.019009385077446178, 32'sd-0.008678995901529008, 32'sd-0.010154003024539933, 32'sd0.05806479474861527, 32'sd0.002470736297355055, 32'sd-0.14085217654594095, 32'sd-0.0640385044354691, 32'sd-0.09621614155389997, 32'sd-0.04982101046921551, 32'sd0.01502760523455737, 32'sd4.9814955224732675e-121, 32'sd6.827713912019901e-115, 32'sd0.04590375812090651, 32'sd-0.06724057308283957, 32'sd0.10259630583311041, 32'sd-0.0037157138566871225, 32'sd-0.04609152875071377, 32'sd0.0243162312864718, 32'sd-0.0843026000332709, 32'sd0.057271269738145184, 32'sd-0.007357094998091634, 32'sd-0.009041437607631705, 32'sd-0.034232197944414275, 32'sd-0.03201287824261578, 32'sd0.04021883555552985, 32'sd0.011837069604710147, 32'sd0.0603461671780636, 32'sd0.05521956246734945, 32'sd0.05926199339923011, 32'sd0.04672447487088049, 32'sd-0.01909349436963365, 32'sd0.07620798068151378, 32'sd0.05110118896920459, 32'sd0.025681647817616563, 32'sd-0.03332867513476895, 32'sd-0.05548144721408836, 32'sd0.044753018355752405, 32'sd-0.1053438308234824, 32'sd0.10433437509768666, 32'sd1.3734521678740562e-123, 32'sd0.05876502899257139, 32'sd0.02417941269988027, 32'sd-0.10947211751031125, 32'sd-0.07347388924786605, 32'sd-0.07895435674119708, 32'sd-0.17520779115518048, 32'sd0.004098744565924451, 32'sd0.0031013904478011424, 32'sd0.10403339897150939, 32'sd0.0704979795059223, 32'sd-0.0658569234072838, 32'sd-0.1118251048769434, 32'sd0.07295894232675418, 32'sd0.02397740509888276, 32'sd0.04242442066543259, 32'sd0.006257562828824181, 32'sd0.10553452554589778, 32'sd0.02886208299395285, 32'sd0.053354120141109504, 32'sd0.06251311039726215, 32'sd0.07341686581116214, 32'sd0.1087962772186377, 32'sd0.10224345463238892, 32'sd0.08394145709362803, 32'sd-0.02479345397473907, 32'sd-0.017924067608497792, 32'sd-0.011720230401023757, 32'sd-1.6210893830799453e-115, 32'sd0.07842254807642902, 32'sd-0.0011956615652302246, 32'sd-0.0046137473362709, 32'sd0.07494172131883194, 32'sd0.04870051961891474, 32'sd-0.03492891307845244, 32'sd-0.11440452623892126, 32'sd0.010872854186370967, 32'sd0.019307522771146883, 32'sd0.035064560456315036, 32'sd-0.01489605895453771, 32'sd0.09551661958464829, 32'sd0.04327238214782093, 32'sd0.00806774888218298, 32'sd-0.022761642514837796, 32'sd0.025850383767318755, 32'sd0.0747989439829067, 32'sd0.16714391525332445, 32'sd0.03045971021810322, 32'sd-0.025928634002912895, 32'sd-0.07314170711129461, 32'sd0.07733452248068334, 32'sd-0.09549632534411746, 32'sd0.10856007250076263, 32'sd0.016765395574197556, 32'sd0.05912986331108688, 32'sd-0.08721070446962964, 32'sd0.06586325306295604, 32'sd0.007813572941118495, 32'sd-0.010762066934662222, 32'sd0.0009322977369508572, 32'sd0.10766283609482868, 32'sd-0.04472762531514785, 32'sd-0.14737500906236078, 32'sd-0.0681783094311409, 32'sd0.00320196893879094, 32'sd-0.04929697253498948, 32'sd0.04807843400573899, 32'sd0.14278973743484075, 32'sd0.08105865031775512, 32'sd0.024643203670930935, 32'sd0.0697148664536125, 32'sd-0.004132904628378205, 32'sd0.042063974194884425, 32'sd0.15506985335050755, 32'sd0.18063198395496816, 32'sd0.06463233059092838, 32'sd0.12355309900188434, 32'sd0.13062895077636932, 32'sd-0.010688408903392302, 32'sd-0.020552154611155202, 32'sd-0.07090173228326563, 32'sd0.04874875393037611, 32'sd0.011696225781014622, 32'sd-0.006587212950685642, 32'sd0.047927359416996385, 32'sd0.1149102468423918, 32'sd-0.005527928798454577, 32'sd0.036964784460326465, 32'sd0.022346869911308437, 32'sd-0.06044074786154735, 32'sd-0.1649865542088067, 32'sd0.03542734798648112, 32'sd0.03433982259657623, 32'sd-0.014214763936384055, 32'sd-0.03321914555959744, 32'sd0.11656233575444692, 32'sd0.20518489032614903, 32'sd0.06008727789793834, 32'sd0.05898715692487242, 32'sd0.017478106049311715, 32'sd0.0576428788611468, 32'sd-0.026180703730519162, 32'sd0.017674856817654804, 32'sd0.08356015385849769, 32'sd0.086402451398253, 32'sd0.09149644313912901, 32'sd-0.018870892298435783, 32'sd-0.08785267055098371, 32'sd-0.013568348093912504, 32'sd0.031902432584422866, 32'sd0.07764692932885094, 32'sd-0.0650407664181471, 32'sd0.047096130977260064, 32'sd0.14347273699612292, 32'sd-0.058575761732904935, 32'sd0.024116292193768957, 32'sd0.07138074434527905, 32'sd-0.035437831897839944, 32'sd0.013896413307710414, 32'sd-0.01406024031391041, 32'sd0.02163004799179125, 32'sd-0.13996656602367188, 32'sd-0.1530261991326143, 32'sd0.018324127090502677, 32'sd0.06950427261264691, 32'sd0.1492985914052522, 32'sd-0.04022652415495682, 32'sd-0.1478298909271317, 32'sd-0.29235907055691135, 32'sd-0.263105308908342, 32'sd-0.04364695835641982, 32'sd0.0197586285441524, 32'sd0.0774686289008026, 32'sd-0.03715025897824273, 32'sd0.07036631775997264, 32'sd-0.08471504675010061, 32'sd0.030644643145308344, 32'sd-0.03021104731857054, 32'sd-0.052494336134582695, 32'sd0.009344833971523244, 32'sd0.06853641428133868, 32'sd0.068102074062931, 32'sd0.10233804293772776, 32'sd-0.04718493871188932, 32'sd0.08695638138322134, 32'sd-0.03366556675391725, 32'sd-0.09238006033066228, 32'sd-0.10837054801138798, 32'sd-0.0018640667831014224, 32'sd-0.04620508593563558, 32'sd0.08973132527921981, 32'sd0.13763247851802124, 32'sd0.10976739635932276, 32'sd0.12734294472988086, 32'sd-0.2111663820684731, 32'sd-0.2534532014520114, 32'sd-0.22771553699180314, 32'sd-0.14809523548950287, 32'sd-0.020748436329962018, 32'sd0.011313501174610587, 32'sd-0.06505726646315578, 32'sd-0.06904564469938583, 32'sd-0.07110576789807554, 32'sd-0.16085846686078867, 32'sd-0.04526994167105706, 32'sd-0.03137365420192408, 32'sd0.01628641184489667, 32'sd0.05723771299131878, 32'sd0.09747736782639183, 32'sd0.09738692564106556, 32'sd-0.021800739242954614, 32'sd0.1016864397331036, 32'sd-0.06668475386240419, 32'sd0.07386066314527233, 32'sd-0.013971968782193402, 32'sd-0.015296342912717182, 32'sd0.008724041062120972, 32'sd0.12979294850098816, 32'sd0.05158297211293178, 32'sd0.17273869609189998, 32'sd0.15020038759559526, 32'sd0.004622572055761712, 32'sd-0.28546060293077663, 32'sd-0.16763302061238403, 32'sd-0.08419528805988045, 32'sd0.038378326159702277, 32'sd0.10249371612577927, 32'sd-0.044110063620749894, 32'sd-0.13235274748364595, 32'sd-0.13238786321566268, 32'sd-0.19104066505865575, 32'sd-0.1507718353861752, 32'sd-0.09302972134169496, 32'sd-0.003883960663833833, 32'sd0.04324240622121864, 32'sd0.0003127312535741326, 32'sd0.029830004909045978, 32'sd-0.018706015327259767, 32'sd0.002835623666837836, 32'sd-0.06976965465061567, 32'sd0.01741933959914203, 32'sd-0.043831549481012755, 32'sd0.02280828033583623, 32'sd0.06947207448970642, 32'sd0.09194841818082697, 32'sd0.0561674638979548, 32'sd0.11700225456564431, 32'sd0.08736485434681332, 32'sd-0.04365964673733296, 32'sd-0.14032731875432877, 32'sd-0.2688683602412705, 32'sd-0.0837083538229681, 32'sd-0.006792282288375316, 32'sd-0.04152827281202562, 32'sd0.13682890564445957, 32'sd-0.1712304113201523, 32'sd-0.08523342230105861, 32'sd-0.0322264636778186, 32'sd-0.20731140863493253, 32'sd-0.16798120995325927, 32'sd-0.03693545776837753, 32'sd-0.07578583746280819, 32'sd0.04171445072405631, 32'sd0.003663768443104629, 32'sd-0.0005305729662920192, 32'sd-0.027285654146583637, 32'sd0.0901938109555187, 32'sd-0.021045308789063615, 32'sd0.0746513214086102, 32'sd0.06599782552717014, 32'sd0.11891364338341694, 32'sd0.10615456465945847, 32'sd0.10066949146299163, 32'sd0.0889218489853354, 32'sd0.10733405151618004, 32'sd-0.050861762384971775, 32'sd-0.02825411661380632, 32'sd-0.17161602177038163, 32'sd-0.12764972499445865, 32'sd-0.18927384472136247, 32'sd-0.14426353119860166, 32'sd-0.04269843283824782, 32'sd-0.026668392300303188, 32'sd0.042006851795336496, 32'sd-0.04636631578083491, 32'sd-0.03409129448043841, 32'sd-0.15449062232122632, 32'sd-0.1494476061824381, 32'sd0.07831618743613059, 32'sd-0.05722757950875229, 32'sd-0.05936961357306102, 32'sd-0.01999073898640506, 32'sd-0.012642752287029399, 32'sd-0.0381008142151622, 32'sd0.013387668237379169, 32'sd-0.07298930838492751, 32'sd0.07647659915070124, 32'sd0.03843952723161786, 32'sd-0.042775026381928746, 32'sd-0.0037992770849993936, 32'sd0.05918303865691512, 32'sd0.03285117630017239, 32'sd-0.050454308194488914, 32'sd-0.05733641246015394, 32'sd-0.034820867060395964, 32'sd-0.1337743375237706, 32'sd-0.18550353564627928, 32'sd-0.13903652112440015, 32'sd-0.0525148471037643, 32'sd-0.11834413180727779, 32'sd-0.04774324357569708, 32'sd0.024141566997997868, 32'sd0.006319855931917247, 32'sd0.029016267245949377, 32'sd-0.056345659621280804, 32'sd-0.13255881521814009, 32'sd0.01160788479457839, 32'sd-0.1470599010043192, 32'sd0.02464993466728495, 32'sd0.08049342839906014, 32'sd-0.027072634549970012, 32'sd0.0004494768510348108, 32'sd0.10710777614335319, 32'sd0.015193019155061244, 32'sd-0.01730791066486657, 32'sd0.025562715514405577, 32'sd-0.13099261882760438, 32'sd-0.03351948234484264, 32'sd-0.17851138138066874, 32'sd-0.08388447606387206, 32'sd-0.01295922792881174, 32'sd-0.09867207033617331, 32'sd-0.0849945625318262, 32'sd-0.03068526609069271, 32'sd-0.09719072126449128, 32'sd-0.11152223795256784, 32'sd-0.06455327443852577, 32'sd0.0029222577593157073, 32'sd0.08171576186921545, 32'sd0.0037293571567983885, 32'sd-0.06435299639037104, 32'sd0.08391958421315399, 32'sd-0.037016759347492934, 32'sd-0.019942345270101993, 32'sd0.026361511608852094, 32'sd-0.10130238642116061, 32'sd-0.021086639801689094, 32'sd0.04636867091468933, 32'sd0.004388720457276989, 32'sd0.03413153889190147, 32'sd0.05886558998201901, 32'sd0.0368430289366832, 32'sd-0.1395640588128784, 32'sd-0.10217149986937904, 32'sd-0.15566124342158483, 32'sd-0.10118933294845195, 32'sd-0.12254139006507361, 32'sd-0.04524269672069336, 32'sd0.05357306377947084, 32'sd0.017491243323368294, 32'sd-0.004786128870306192, 32'sd-0.1711327067432045, 32'sd-0.098447168884029, 32'sd-0.05425888749648357, 32'sd-0.06716750364211971, 32'sd0.04887986030109002, 32'sd0.08104381885707677, 32'sd0.02840982133533433, 32'sd0.03364346623163494, 32'sd0.08940224547076536, 32'sd0.13354565818296135, 32'sd-0.02920859597451489, 32'sd-0.01967863611043591, 32'sd-0.038727970305619024, 32'sd0.018122332223881234, 32'sd-0.04278539812672915, 32'sd3.962699236461415e-123, 32'sd0.014152423209941152, 32'sd-0.04873986840256607, 32'sd0.008790556380317434, 32'sd-0.11724923898269472, 32'sd-0.0996009567760251, 32'sd-0.03518136207297982, 32'sd0.07104787491247888, 32'sd-0.15028360703199078, 32'sd-0.10160690938166125, 32'sd0.06609167992962868, 32'sd-0.11478271016217624, 32'sd-0.093905837354635, 32'sd-0.04214244068154242, 32'sd-0.14104808000512034, 32'sd-0.19236800935096954, 32'sd-0.10988450833821006, 32'sd0.008679517198661122, 32'sd0.1219973904152167, 32'sd0.11091711367940645, 32'sd0.0651800532049905, 32'sd0.07727156559153889, 32'sd0.07573989416614657, 32'sd-0.06038834138081081, 32'sd0.06628106801730396, 32'sd-0.025647045822311143, 32'sd-0.012623010315616063, 32'sd0.0707034408441079, 32'sd-0.00444046582264758, 32'sd0.08760285436497421, 32'sd0.05621743372713205, 32'sd0.02978189901273923, 32'sd-0.07706911526975867, 32'sd-0.17232812662725025, 32'sd-0.10086976497847186, 32'sd-0.04319767900313911, 32'sd-0.05826598772712946, 32'sd0.002814269738873369, 32'sd-0.012607787328846936, 32'sd-0.07119349710895632, 32'sd0.03467272678301698, 32'sd-0.15449811603965036, 32'sd-0.16109572043933607, 32'sd-0.17565244462018598, 32'sd-0.06691275851756773, 32'sd-0.007946321134811434, 32'sd0.07774851123402043, 32'sd0.023510858930890825, 32'sd0.06681096739680242, 32'sd0.05389172058598325, 32'sd-0.041380567202110516, 32'sd0.005942658690820356, 32'sd-0.06822648643163762, 32'sd-0.08017052061205268, 32'sd0.016103554237897798, 32'sd-0.04253319950505363, 32'sd0.009409246025441204, 32'sd0.022988156265422215, 32'sd0.09320097431330011, 32'sd0.04984905790160351, 32'sd-0.018444876741853435, 32'sd-0.0525159653690005, 32'sd-0.07474171740020966, 32'sd-0.056383065313121386, 32'sd-0.14501818426709778, 32'sd-0.06077374697846712, 32'sd-0.19736310853768851, 32'sd-0.031402322430803896, 32'sd-0.037089168221681706, 32'sd-0.004213140819520603, 32'sd-0.0763187787657035, 32'sd-0.12893779402505526, 32'sd-0.037777539135020514, 32'sd0.10507341176890968, 32'sd0.05855844678078963, 32'sd-0.09361528668459017, 32'sd0.0875058212658959, 32'sd-0.05338548557568469, 32'sd0.050792039435518556, 32'sd-0.034345390557936395, 32'sd-0.0031624240151308567, 32'sd-0.0003000489091336682, 32'sd-0.03925298665232678, 32'sd-0.05489596863560852, 32'sd-3.790147288667311e-119, 32'sd-0.042062222351671126, 32'sd-0.08913928811456077, 32'sd0.10007874543752836, 32'sd0.024531493732157714, 32'sd-0.10742587014221433, 32'sd-0.05509031373364264, 32'sd-0.06881357609967662, 32'sd-0.0071998455862457705, 32'sd-0.013155323843886159, 32'sd-0.06055042136155552, 32'sd0.009703255724976823, 32'sd0.028723077797002106, 32'sd0.02126806420282581, 32'sd0.04644835819336841, 32'sd-0.002788088799393394, 32'sd-0.048141218026738625, 32'sd-0.03963694896010656, 32'sd-0.09388705700365492, 32'sd-0.0411933531447801, 32'sd0.030270798219719133, 32'sd0.005888739197524865, 32'sd0.06679454497241005, 32'sd0.05321551698979974, 32'sd-0.00734328205759397, 32'sd-0.08482873619560291, 32'sd-0.04896088703731161, 32'sd0.03938994125170029, 32'sd0.04535033929616786, 32'sd0.028599860796931602, 32'sd0.01837533284614366, 32'sd0.000878159855774577, 32'sd0.0020328065765989915, 32'sd-0.13669600450083533, 32'sd-0.09051392784069992, 32'sd-0.1250412677447097, 32'sd0.008582255755961528, 32'sd0.05141740701483902, 32'sd0.05652055026584591, 32'sd0.08006822578052761, 32'sd0.13909193223699087, 32'sd0.14043038691044887, 32'sd0.0884389358645901, 32'sd0.12275143164828636, 32'sd0.013857717165634042, 32'sd-0.03385401365097722, 32'sd0.02873710856787318, 32'sd-0.10442954903411157, 32'sd-0.015876569966321887, 32'sd0.04810408829416166, 32'sd0.12928697037415074, 32'sd0.021140897130665533, 32'sd-0.09006876638411156, 32'sd-0.018127152288852002, 32'sd0.012199217803739107, 32'sd-0.016869610334605184, 32'sd0.02824860747841814, 32'sd0.04010837194954168, 32'sd-0.018857849383321534, 32'sd-0.08269334390045442, 32'sd-0.04437080261879513, 32'sd-0.08918031180340046, 32'sd-0.15150715395918266, 32'sd-0.11982470682942765, 32'sd0.0023617876083418883, 32'sd0.056580245458263345, 32'sd-0.06035384577194287, 32'sd0.14092839096894033, 32'sd0.16205349616167086, 32'sd0.15599726868261884, 32'sd-0.003487249367156006, 32'sd0.1550409374286064, 32'sd0.18451346926484796, 32'sd-0.06446095565534378, 32'sd0.009362448370534675, 32'sd0.004301597108434175, 32'sd0.026832863771531407, 32'sd-0.08627937254689738, 32'sd0.06148888287618797, 32'sd0.06698694207506281, 32'sd-0.08571424661063755, 32'sd-0.132788341601685, 32'sd0.045050463673198905, 32'sd0.06513397922570241, 32'sd-2.1708707061370033e-127, 32'sd0.05523930620682579, 32'sd-0.0282822438714662, 32'sd0.011590708999937287, 32'sd-0.06650535268983163, 32'sd0.040699010578647464, 32'sd-0.03796038335681349, 32'sd0.015515113093025635, 32'sd0.034883142970775605, 32'sd0.10903003525450816, 32'sd0.11658299868951584, 32'sd0.14129523257460325, 32'sd0.044395241742166136, 32'sd0.07772455446742481, 32'sd0.06961037628584753, 32'sd0.016719676028824047, 32'sd-0.031725658248218935, 32'sd0.11334435349247333, 32'sd0.07900964632689605, 32'sd0.06583728912026808, 32'sd-0.1261211650946622, 32'sd-0.015117889201166508, 32'sd-0.004051795390631003, 32'sd0.09241602742984166, 32'sd-0.1048462072959383, 32'sd-0.10246877810024732, 32'sd-0.01090101373569802, 32'sd4.3617634543407303e-122, 32'sd-2.623243146627509e-122, 32'sd-4.7969311755681075e-129, 32'sd0.0025615217368587, 32'sd-0.023354496624552898, 32'sd0.03786454991822104, 32'sd0.07736872374709103, 32'sd0.03691246479505837, 32'sd0.06539929188580952, 32'sd0.16219273632555184, 32'sd0.209730863982502, 32'sd0.1352651550860545, 32'sd0.011472745720273639, 32'sd0.10277589309680457, 32'sd-0.009602948184026436, 32'sd0.03606973286478353, 32'sd0.09727673943776745, 32'sd0.08450095994348462, 32'sd0.1266167182417977, 32'sd0.1019674543140877, 32'sd0.1495516579833551, 32'sd-0.06071514478696683, 32'sd-0.03296663905133585, 32'sd-0.0029951128407539056, 32'sd-0.1050702102178598, 32'sd0.001260469675039101, 32'sd0.049173187365180886, 32'sd0.02272367039023608, 32'sd1.0285481442363402e-119, 32'sd-4.863506894779109e-127, 32'sd-4.874500825880841e-123, 32'sd-0.0160572842810474, 32'sd0.0373348646338777, 32'sd-0.01280304663821434, 32'sd-0.016840236378408792, 32'sd0.031184913497772034, 32'sd0.11184985877734052, 32'sd0.0645968046881024, 32'sd0.16416692599662627, 32'sd0.006518250925789916, 32'sd0.04210036899034018, 32'sd0.08975714167911368, 32'sd0.12790152279245715, 32'sd-0.1048542500770137, 32'sd-0.006505238473652445, 32'sd-0.02339100559523084, 32'sd0.0130131227691091, 32'sd0.018023879109005762, 32'sd0.014303425247033494, 32'sd0.11271034440387952, 32'sd-0.05058184498454483, 32'sd0.008027274351762478, 32'sd-0.007108878033630089, 32'sd0.002707306688029642, 32'sd-0.00670336451894657, 32'sd0.07306046424479358, 32'sd-2.1110341548608268e-119, 32'sd2.076836201097574e-117, 32'sd-1.1821509009281003e-121, 32'sd1.0211617841978798e-120, 32'sd0.020231590794618493, 32'sd0.04277992441372465, 32'sd-0.1482060127724277, 32'sd-0.023160932824266952, 32'sd0.034449468420314565, 32'sd-0.026018213258953864, 32'sd0.11977134985126073, 32'sd0.04287209113226752, 32'sd0.05239755555000962, 32'sd0.1474045202797834, 32'sd0.056945466975692395, 32'sd-0.003916609843355927, 32'sd0.09106442991261932, 32'sd0.12335591209740729, 32'sd0.035161409006117056, 32'sd0.07060507599791864, 32'sd0.03945501977198847, 32'sd-0.0799997159308905, 32'sd-0.05706785973573222, 32'sd-0.048926782881877795, 32'sd-0.024797105726176424, 32'sd-0.012167224706807046, 32'sd0.023482899703437945, 32'sd-2.628925132047927e-121, 32'sd1.6137253275161974e-115, 32'sd-7.433039422476896e-115, 32'sd-6.431337471154935e-127, 32'sd-1.7015398108253827e-126, 32'sd2.6226419133016735e-125, 32'sd0.09443042752381407, 32'sd0.013513878814201647, 32'sd-0.01792619632120952, 32'sd0.08616146185735334, 32'sd0.06415815868336464, 32'sd0.013071032831208567, 32'sd0.015124122820938328, 32'sd0.04672750507404765, 32'sd0.0650540459094202, 32'sd0.10353399772380674, 32'sd0.01096745076728269, 32'sd0.040593361105209065, 32'sd-0.02357851309094428, 32'sd0.12953263418473238, 32'sd0.0018531217966617777, 32'sd0.0038091795684126726, 32'sd-0.0010141864911508644, 32'sd-0.015015581982542242, 32'sd-0.011665052595110446, 32'sd0.019375728439875253, 32'sd-3.7900837736976324e-122, 32'sd-2.625910146497655e-119, 32'sd-2.689673124678537e-124, 32'sd5.209870900506999e-118},
        '{32'sd-4.963021604824245e-115, 32'sd5.1902553978247746e-126, 32'sd5.730051323098458e-125, 32'sd1.313916584104527e-126, 32'sd-1.697400632837211e-121, 32'sd-2.547163601687575e-122, 32'sd-2.7836136623306796e-123, 32'sd-1.3188572745419073e-117, 32'sd-1.0505622148352857e-124, 32'sd-5.081937622007938e-118, 32'sd7.720499004881737e-123, 32'sd6.240517699308852e-124, 32'sd0.041603735823194266, 32'sd-0.044981764097226214, 32'sd0.07425714371613462, 32'sd0.0855230411184068, 32'sd6.3573336085892624e-127, 32'sd7.879898006910994e-127, 32'sd-1.5765559740072215e-117, 32'sd-1.8640399554972862e-125, 32'sd3.590619915288838e-122, 32'sd1.2521555509931131e-117, 32'sd-2.11669148916708e-124, 32'sd3.348446431751269e-123, 32'sd2.0123090973335696e-118, 32'sd1.5142686547272657e-119, 32'sd-3.358551156460452e-121, 32'sd1.0066144452798187e-122, 32'sd6.633215443048932e-118, 32'sd-2.5056145193509065e-124, 32'sd9.100397300228472e-118, 32'sd2.039880754628471e-127, 32'sd-0.035813269615102825, 32'sd0.05257075738491231, 32'sd0.08468551913415061, 32'sd0.0017010309888880108, 32'sd-0.04509027101083048, 32'sd0.07483569197052004, 32'sd-0.010386916013671798, 32'sd-0.0853076923204324, 32'sd-0.11155564267416523, 32'sd-0.016066915887257924, 32'sd0.01958887368772185, 32'sd0.006434152122977391, 32'sd0.07735753173037727, 32'sd-0.0741869053975554, 32'sd-0.06649201125933354, 32'sd-0.010071900039379007, 32'sd-0.02569122115070218, 32'sd-0.060205876365691975, 32'sd-0.012799171087438253, 32'sd-0.018952587037407435, 32'sd-4.283145558415494e-118, 32'sd-2.0105118012862036e-123, 32'sd-4.224805864788299e-125, 32'sd1.8190116893596383e-123, 32'sd4.787381912076311e-123, 32'sd-1.1108297261035896e-124, 32'sd-0.01474546023262422, 32'sd-0.056283136883080585, 32'sd-0.11886196568274085, 32'sd-0.09178280153990272, 32'sd0.002781575951497858, 32'sd0.062441019100526664, 32'sd-0.04294581759907293, 32'sd-0.0959092108316785, 32'sd-0.029663725736000797, 32'sd-0.019934524409104187, 32'sd-0.1701783817132324, 32'sd-0.03844507671075384, 32'sd-0.13410174939833627, 32'sd-0.09360764068840793, 32'sd0.032278141960220476, 32'sd-0.08555133529517234, 32'sd-0.017303511368192845, 32'sd0.08469902741832916, 32'sd-0.04501024124139598, 32'sd0.019649773668133, 32'sd-0.13170285948301969, 32'sd-0.0521119988114955, 32'sd0.025780937391968867, 32'sd-0.010529735189782756, 32'sd-2.7094034194303004e-124, 32'sd-3.5348010345180936e-122, 32'sd5.404737460235472e-125, 32'sd-1.5490405061186628e-115, 32'sd0.010477714801189697, 32'sd0.07191444409102976, 32'sd0.02103502144868551, 32'sd0.04336361713690903, 32'sd-0.051769515927344315, 32'sd-0.04264543986898663, 32'sd-0.10556571972289863, 32'sd0.06235295237779247, 32'sd-0.03182488037528903, 32'sd-0.12559950157997918, 32'sd-0.06714309382792745, 32'sd-0.14809199383587904, 32'sd-0.05453800673832778, 32'sd0.06121621809603992, 32'sd0.04819968975484705, 32'sd-0.0984976776833093, 32'sd-0.17025928162608742, 32'sd-0.062366176336587434, 32'sd-0.020897511471103233, 32'sd-0.051732809553632256, 32'sd0.039093760233170474, 32'sd-0.0606605199528422, 32'sd0.07501239438085726, 32'sd0.023820023092700312, 32'sd0.03354625000207151, 32'sd2.2424054801188887e-121, 32'sd-4.2070112870333694e-125, 32'sd-0.030236851100196038, 32'sd0.05140207017452937, 32'sd0.004877002628226055, 32'sd-0.031222370250169412, 32'sd-0.06508824147978727, 32'sd-0.014673473950311995, 32'sd-0.06437732757764512, 32'sd-0.20223244174921234, 32'sd-0.07756520414110459, 32'sd-0.10595610369034333, 32'sd-0.06521769625057514, 32'sd0.016212243242528675, 32'sd-0.08706114534992933, 32'sd-0.06833843752148283, 32'sd-0.03991300602883398, 32'sd-0.034700910066221675, 32'sd-0.01597257450226885, 32'sd0.01085775878691212, 32'sd-0.05409492744892822, 32'sd0.08406508934567192, 32'sd-0.030265663208291584, 32'sd0.05397332611329921, 32'sd-0.1102638985861296, 32'sd-0.09342454492808064, 32'sd0.04881517505470907, 32'sd0.07943833287243873, 32'sd0.011759960983660594, 32'sd6.246640189796453e-126, 32'sd-0.036057133846532655, 32'sd-0.09845346125193853, 32'sd0.028234814692583904, 32'sd0.002302259290873083, 32'sd-0.1308139440477556, 32'sd-0.11844995719554746, 32'sd-0.12505778272893045, 32'sd-0.0873672353576418, 32'sd-0.10793308531483216, 32'sd-0.00011837788153880775, 32'sd0.005163928791703905, 32'sd0.0033622634796710506, 32'sd0.2216361726684412, 32'sd0.11785567206247019, 32'sd0.06423575358154486, 32'sd-0.09377889115855227, 32'sd-0.0638831761737295, 32'sd-0.0022565566843066333, 32'sd0.06890252921583365, 32'sd-0.031096292396796437, 32'sd-0.1477217061669388, 32'sd-0.01347165987641195, 32'sd-0.18314782643509797, 32'sd-0.08568794919687588, 32'sd-0.06275241248018246, 32'sd0.03937537783487291, 32'sd-0.021278409698954694, 32'sd1.9099559498239014e-126, 32'sd-0.021836352324224567, 32'sd-0.025237586459404573, 32'sd-0.09655260031656063, 32'sd-0.01984902225001604, 32'sd-0.17431082688825314, 32'sd-0.10586357700617997, 32'sd-0.0392660600043972, 32'sd-0.0462436068206241, 32'sd-0.025472991211180074, 32'sd-0.012368633650252602, 32'sd0.0187755088609978, 32'sd0.03359822264764267, 32'sd0.03310980857008125, 32'sd0.00618473149109053, 32'sd0.022887018272571877, 32'sd0.08806093967151096, 32'sd0.08564956485617782, 32'sd0.10787691277642478, 32'sd-0.00024039726618409288, 32'sd0.057436947283954355, 32'sd0.05923281893700201, 32'sd0.04298092931066576, 32'sd-0.07026616913819063, 32'sd-0.029579682438400753, 32'sd-0.01474913795880013, 32'sd-0.12189127828539671, 32'sd0.05617446521302801, 32'sd0.03291776962523219, 32'sd-0.014758590309879756, 32'sd0.013943778562079292, 32'sd-0.018965753986590974, 32'sd0.05754646902575603, 32'sd-0.14522586892483896, 32'sd-0.14954919049307472, 32'sd-0.06274699326400703, 32'sd-0.03987263098287641, 32'sd0.003490252661274567, 32'sd0.05697631502734696, 32'sd0.026591397280921043, 32'sd0.006687649393673594, 32'sd-0.04714851296837404, 32'sd0.00416233879335064, 32'sd0.0027834531175522717, 32'sd0.09260285380330982, 32'sd0.07372489029106083, 32'sd0.14255761908616624, 32'sd0.13516666377379336, 32'sd0.03461191325378464, 32'sd-0.010169338416292986, 32'sd-0.009338285317254546, 32'sd0.029039143509671347, 32'sd0.09713779772440558, 32'sd0.026847617245739447, 32'sd-0.1457448755200146, 32'sd-0.02235936491021628, 32'sd0.018814970024011834, 32'sd0.016486643695630937, 32'sd0.068543545852803, 32'sd-0.08043415270346979, 32'sd-0.04649893003091061, 32'sd-0.0017639776501819423, 32'sd0.010216353137961712, 32'sd-0.08450057290761737, 32'sd-0.014375109197134295, 32'sd-0.038089303253873996, 32'sd0.05691204429254232, 32'sd-0.020906036381089683, 32'sd-0.013068409068733477, 32'sd-0.0639364645956002, 32'sd0.07609772685149155, 32'sd0.23549726093936188, 32'sd0.26404015803920305, 32'sd0.16445525085402754, 32'sd0.040945959003659896, 32'sd0.1240704257181296, 32'sd0.002900505200510723, 32'sd0.03845129242550998, 32'sd-0.04791680017215445, 32'sd0.06131338305935754, 32'sd0.04375817048506077, 32'sd0.09594898839568484, 32'sd-0.0714389561740386, 32'sd-0.05025056380367117, 32'sd-0.06787861642885384, 32'sd-0.07997202499447698, 32'sd-0.04796970818192791, 32'sd-0.059274479616662164, 32'sd0.049764978261543746, 32'sd-0.07900960457252713, 32'sd0.12543519305387765, 32'sd0.027624766077126245, 32'sd-0.053403146828452375, 32'sd0.017935851866587405, 32'sd0.07915100627978833, 32'sd-0.028445997463553477, 32'sd-0.009081363573029853, 32'sd0.06640527289522838, 32'sd0.02526601529409053, 32'sd0.07321342809245873, 32'sd0.11736221799442212, 32'sd0.042666468271174554, 32'sd0.06853821110452518, 32'sd0.07101229826326026, 32'sd0.22597082107980226, 32'sd0.06969673806664539, 32'sd-0.039231225092355874, 32'sd0.0005447584551175886, 32'sd0.058600475022252504, 32'sd-0.002228164183167295, 32'sd-0.059586071882134835, 32'sd-0.041923927078502086, 32'sd0.030719748922035106, 32'sd0.0029016884184387736, 32'sd-0.05611158438668365, 32'sd0.06998948208155732, 32'sd0.021193376723262727, 32'sd0.05579560020924045, 32'sd0.011827362362885325, 32'sd-0.06346771236335948, 32'sd-0.04186230523166935, 32'sd0.0059753459376413525, 32'sd0.06376781170632408, 32'sd0.10032878311092298, 32'sd0.027460253717197368, 32'sd-0.0401858694320515, 32'sd0.003317244362276784, 32'sd0.018212573366421392, 32'sd-0.05302156631370333, 32'sd-0.04656550052983124, 32'sd-0.018851720712766935, 32'sd0.01915151475173127, 32'sd0.12881288932307836, 32'sd0.12421167824279779, 32'sd0.07008998847299147, 32'sd0.02453940072941113, 32'sd0.07128292122377008, 32'sd-0.025245534450622154, 32'sd-0.06738354696335433, 32'sd-0.02364506986249053, 32'sd0.025031202667124088, 32'sd0.06653415791345162, 32'sd0.02640569487418031, 32'sd-0.019501257813055336, 32'sd-0.06817051111298846, 32'sd0.05429108135429429, 32'sd0.018637886216226033, 32'sd-0.01258895479522768, 32'sd-0.07536316049445997, 32'sd-0.11084572002198745, 32'sd0.06774109341273478, 32'sd-0.025347592699649684, 32'sd-0.08756533860884062, 32'sd-0.03294211604143342, 32'sd-0.13229170318050268, 32'sd-0.14917913228700083, 32'sd-0.037413412519570796, 32'sd-0.043617328790656176, 32'sd-0.041161743042532235, 32'sd0.024379272873121794, 32'sd0.14281983348314822, 32'sd0.0961153999773863, 32'sd0.04977959651576008, 32'sd-0.09610426134098018, 32'sd0.07397022079273104, 32'sd0.07214331049040042, 32'sd0.08225273993753901, 32'sd-0.07687755120315715, 32'sd0.057201692276142656, 32'sd0.03665179187145784, 32'sd-0.1168154523161963, 32'sd0.04356443543543017, 32'sd0.07882530120541512, 32'sd0.07515093304388519, 32'sd0.1056952671473795, 32'sd-0.023101185261577978, 32'sd-0.0734380875799757, 32'sd-0.14033167394404836, 32'sd1.7470214270353712e-05, 32'sd0.037550924854793236, 32'sd-0.13691229421727188, 32'sd-0.09065020185669925, 32'sd-0.05250186939859021, 32'sd0.014338495174029015, 32'sd-0.023365479822048875, 32'sd-0.04921968705023174, 32'sd0.08998431755396316, 32'sd0.23734305968510339, 32'sd0.15047781892966453, 32'sd0.0625450539611356, 32'sd0.014679751074884749, 32'sd0.046080972867241596, 32'sd-0.02327202003279821, 32'sd-0.01524964515466627, 32'sd-0.020410345491566426, 32'sd0.025986117664651878, 32'sd-0.00655886673623899, 32'sd-0.0746299925300977, 32'sd0.03853421284531616, 32'sd0.0021610835477227476, 32'sd-0.005954333657690017, 32'sd0.015054975259247285, 32'sd0.10759135826727416, 32'sd0.09670757028307728, 32'sd-0.07632170521823058, 32'sd-0.14462563491454866, 32'sd-0.05084343085579971, 32'sd-0.12067074340705053, 32'sd0.06209988294125824, 32'sd-0.051949466963027165, 32'sd0.057180007637427185, 32'sd-0.041804803192244604, 32'sd-0.08563394555139871, 32'sd-0.0704225937891441, 32'sd0.07837362586223535, 32'sd0.18740920957624158, 32'sd0.09562636163631166, 32'sd0.059602683791713976, 32'sd0.018943077301768734, 32'sd-0.02531476633612427, 32'sd-0.22548020864812848, 32'sd-0.020877855612840085, 32'sd0.00442834831779444, 32'sd-0.05292700422288646, 32'sd-0.04726453475238594, 32'sd-0.009471515510132129, 32'sd-0.06110176836119592, 32'sd-0.07985303535361017, 32'sd0.14032480844197262, 32'sd-0.020340253434414715, 32'sd0.1499386575895223, 32'sd0.07794849370738215, 32'sd0.12937936290399088, 32'sd0.1009864590898579, 32'sd0.030225565306720697, 32'sd0.11268653741603445, 32'sd0.00042143805362293183, 32'sd-0.004382098535075308, 32'sd0.07629839584321155, 32'sd-0.08148002531127944, 32'sd-0.15194175816901545, 32'sd-0.010478406206371077, 32'sd0.16195827389513473, 32'sd0.12639748878526, 32'sd0.014630817894703356, 32'sd0.06163715514437938, 32'sd0.019432919980345645, 32'sd-0.020533709322946948, 32'sd-0.07227720823092533, 32'sd-0.03454753574763215, 32'sd0.1770806150844797, 32'sd-0.028430556206945654, 32'sd-0.0180267001026417, 32'sd-0.037118008743679855, 32'sd0.019977191859203765, 32'sd-0.02497676578627958, 32'sd0.08013318828622767, 32'sd0.1470085571102061, 32'sd0.06708365408795983, 32'sd0.18850361228871343, 32'sd0.14339737999674915, 32'sd0.08393896617407001, 32'sd0.10746768220362177, 32'sd-0.08392038498718626, 32'sd-0.011911681502505904, 32'sd-0.08405499545720672, 32'sd0.027951388153884604, 32'sd-0.10960752176630247, 32'sd-0.02970497261059504, 32'sd0.04605166900987184, 32'sd0.025253452347644582, 32'sd0.06711532279631517, 32'sd0.0724721825296054, 32'sd0.023311135716838145, 32'sd0.00923463995641948, 32'sd-0.08049680583774171, 32'sd0.03684966221987671, 32'sd0.028513926635387366, 32'sd0.13582851145555538, 32'sd-0.03833599243940808, 32'sd-0.04366448157599582, 32'sd-0.06205997395147899, 32'sd-0.032484299546796894, 32'sd-0.04794199282466475, 32'sd0.07148774748312131, 32'sd0.04722221021696175, 32'sd0.04412932449904493, 32'sd0.07464194927430148, 32'sd0.08763382895768312, 32'sd0.031193750927163692, 32'sd-0.0295539868629845, 32'sd-0.04199094577096337, 32'sd0.016218226051622826, 32'sd0.07046828744682211, 32'sd0.011416433513567794, 32'sd-0.0051972030587511394, 32'sd0.00570095785916289, 32'sd0.018433153930847317, 32'sd0.1113954575947818, 32'sd-0.08445571117678162, 32'sd-0.07445616990656813, 32'sd-0.0485068326778576, 32'sd0.00026199982164914196, 32'sd-0.11020400101967864, 32'sd-0.023250376470695517, 32'sd-0.07614832606352956, 32'sd0.03688268394432625, 32'sd-0.02851692811250219, 32'sd2.438017509747254e-115, 32'sd-0.06182885039659732, 32'sd0.008565895619702698, 32'sd-0.02754625122856363, 32'sd0.04423268831082883, 32'sd-0.06578723163039099, 32'sd-0.03083828211678673, 32'sd0.07583742568266856, 32'sd0.09031026902215142, 32'sd0.22189944893552657, 32'sd0.1045678134814338, 32'sd0.0783518013576694, 32'sd-0.03946238995447117, 32'sd-0.04470182188196332, 32'sd-0.07031614806638924, 32'sd0.01731747122475853, 32'sd0.031264266376414065, 32'sd0.030209690996898818, 32'sd-0.04735677210508471, 32'sd-0.027325538592670506, 32'sd0.07212063061901254, 32'sd0.036404654326629295, 32'sd-0.06524624217093952, 32'sd-0.10498636641967975, 32'sd0.04635492788650554, 32'sd0.062416225653382465, 32'sd-0.04298599610672512, 32'sd0.03966144261578505, 32'sd0.06732491860653361, 32'sd0.050749449574184535, 32'sd0.013217636981922742, 32'sd-0.1296948684529789, 32'sd-0.08622362511055685, 32'sd-0.10511867478502744, 32'sd-0.04466246658895829, 32'sd0.04838264686440925, 32'sd0.02023082468152957, 32'sd0.06503087733492946, 32'sd0.12614842028212697, 32'sd0.08734933097249352, 32'sd0.02483790268025606, 32'sd0.01409331747561038, 32'sd0.12176934612766385, 32'sd-0.008646125036302297, 32'sd-0.10767569839334402, 32'sd0.013495567172779182, 32'sd-0.027793587946169065, 32'sd0.03361379898432498, 32'sd0.06867960615703039, 32'sd0.11630269604265832, 32'sd-0.067909763857523, 32'sd-0.032457093626093544, 32'sd0.023173010398703692, 32'sd-0.04590496175676507, 32'sd-0.05154175633012912, 32'sd-0.03124664621531224, 32'sd0.024918537148476135, 32'sd-0.032449532250090986, 32'sd0.014914513412666593, 32'sd0.03914597465785112, 32'sd-0.1391847823393943, 32'sd-0.11013379929378105, 32'sd-0.008243336464805805, 32'sd0.06414526604914267, 32'sd0.05863790821426284, 32'sd-0.07700818693590572, 32'sd-0.03020750025451702, 32'sd0.04984938389100961, 32'sd0.16861070330095498, 32'sd0.1307779672423933, 32'sd0.06838977524555381, 32'sd-0.05244559733630722, 32'sd0.05035430096856537, 32'sd-0.04946766484278561, 32'sd0.09013276295474308, 32'sd0.13214952823702972, 32'sd-0.06313727412746976, 32'sd0.10421574642923084, 32'sd-0.09819620512536341, 32'sd-0.11696073235158166, 32'sd0.04427826043500527, 32'sd-0.0615413756435882, 32'sd-0.030328962400098518, 32'sd-0.06726714420036316, 32'sd1.6326604092089168e-115, 32'sd0.08509425780821604, 32'sd-0.15861082229646054, 32'sd-0.009765215174053172, 32'sd0.03142881474810158, 32'sd0.048044406000351175, 32'sd0.0022096709084606053, 32'sd0.013625858366888415, 32'sd-0.04302574513241162, 32'sd-0.1409071913345994, 32'sd-0.045724889411840025, 32'sd-0.01847422032364559, 32'sd0.10257096878621642, 32'sd0.04110356327841117, 32'sd0.002948139236730817, 32'sd-0.12175087574786324, 32'sd-0.015376318076414121, 32'sd0.022026424999718804, 32'sd0.10503489958660478, 32'sd0.0863978599683425, 32'sd0.010590703929812937, 32'sd0.16279352678367223, 32'sd-0.06725073501668599, 32'sd-0.12611968571040647, 32'sd-0.034885526402533173, 32'sd0.06695887588979561, 32'sd0.059992260135905466, 32'sd-0.038001986220058376, 32'sd0.014228666366125665, 32'sd-0.0756059541107263, 32'sd-0.02688099909030506, 32'sd0.0074924989186788485, 32'sd0.056792677549611204, 32'sd0.060508143457179545, 32'sd0.11680909274603775, 32'sd0.09501381517152278, 32'sd-0.025853550230254714, 32'sd-0.1530686270558844, 32'sd-0.020996014779120237, 32'sd-0.012819516427905452, 32'sd0.06210024027255318, 32'sd-0.06412828279311986, 32'sd0.005036275103189223, 32'sd-0.10205509657272958, 32'sd0.047297854216039124, 32'sd-0.1065062631825506, 32'sd0.020713708834634626, 32'sd0.02972160724308793, 32'sd0.028094182714630975, 32'sd0.04540516121524594, 32'sd0.07446772386165162, 32'sd-0.08350434838118127, 32'sd-0.0543411870309763, 32'sd0.036317716762778195, 32'sd0.10515242296651657, 32'sd-0.04289100375364073, 32'sd0.004194653641322364, 32'sd-0.07890721995604658, 32'sd0.0012257254225378608, 32'sd0.039006489091372706, 32'sd-0.038726247764443424, 32'sd0.08690233197948145, 32'sd0.14341658753694972, 32'sd-0.01052519037524223, 32'sd0.013643547847904228, 32'sd0.057089809706572105, 32'sd-0.004233341593820991, 32'sd0.025041661036296736, 32'sd0.017622694827407283, 32'sd-0.0505087623719526, 32'sd-0.10398643030651533, 32'sd-0.08168955084470553, 32'sd-0.03783573255176861, 32'sd0.01382506239218234, 32'sd0.05382804668169039, 32'sd-0.030723800104016815, 32'sd-0.025794405409555465, 32'sd0.1297517913599361, 32'sd0.055443114911102855, 32'sd-0.08807491432943615, 32'sd-0.040686398327718344, 32'sd-0.04551921103806905, 32'sd0.12269646787323585, 32'sd0.0042977178650537955, 32'sd1.3144593343671997e-122, 32'sd-0.04877651295827338, 32'sd-0.015297626635045481, 32'sd0.019449779999019073, 32'sd-0.12555587850517022, 32'sd-0.09286977994368543, 32'sd0.03438267131489529, 32'sd0.003242202072521796, 32'sd0.053111513740521664, 32'sd-0.023691521015755293, 32'sd-0.06659361137860978, 32'sd0.05894427781517781, 32'sd0.012055938212117716, 32'sd-0.011087327774477615, 32'sd-0.022757046167351736, 32'sd0.04385791727495514, 32'sd-0.043521681452883515, 32'sd-0.07731698610561642, 32'sd-0.08058902243376923, 32'sd-0.04556301924373877, 32'sd0.09775839388352278, 32'sd-0.0029086760666022214, 32'sd0.08056511729796136, 32'sd0.05022853897187481, 32'sd-0.01027050072605342, 32'sd0.022130541058199227, 32'sd-0.027986991530491955, 32'sd1.2712245799304389e-117, 32'sd-6.321378117261921e-122, 32'sd-2.3816904815485267e-124, 32'sd0.006439558599620794, 32'sd0.09105489387140157, 32'sd0.09974788791315238, 32'sd0.017751795095259777, 32'sd-0.03212879632156929, 32'sd-0.01910164883957125, 32'sd0.05830903100455204, 32'sd0.05123474928123325, 32'sd-0.060178946885581494, 32'sd-0.1022359381893097, 32'sd-0.035620874717285145, 32'sd-0.10380063105342868, 32'sd-0.058797229581194155, 32'sd-0.04584173455035559, 32'sd0.02299883241469726, 32'sd-0.05591762862355505, 32'sd-0.01997451129592954, 32'sd0.08642779127188668, 32'sd0.056695035805571135, 32'sd-0.006892015444146369, 32'sd-0.01467318961236662, 32'sd0.02656974905128908, 32'sd0.10329147884017303, 32'sd-0.0342926647487735, 32'sd-0.011376341966764979, 32'sd-1.0128979986024444e-124, 32'sd5.282591977563849e-119, 32'sd1.9071888985990962e-127, 32'sd0.06096439945189483, 32'sd-0.04893240085297974, 32'sd0.005200231569954901, 32'sd0.08562943743941054, 32'sd-0.0030655251376737274, 32'sd0.021815479107444524, 32'sd0.05837214141430516, 32'sd0.010819806290234539, 32'sd-0.045079327620717445, 32'sd-0.033894155760517894, 32'sd-0.11901504907093792, 32'sd-0.20507184428235153, 32'sd-0.04597001869489458, 32'sd-0.08987467366927333, 32'sd-0.14133709455287174, 32'sd-0.176389508905756, 32'sd-0.06586006758814898, 32'sd-0.006676715919913366, 32'sd0.02582735687369698, 32'sd-0.03317917039191212, 32'sd0.04299163762377199, 32'sd-0.035839177587175135, 32'sd0.005372994019964952, 32'sd0.07878926281869014, 32'sd-0.04613323095955438, 32'sd-1.953884655576151e-119, 32'sd-1.0786852350801856e-121, 32'sd-2.491737665194321e-124, 32'sd2.597759052254249e-120, 32'sd0.0003300896243779705, 32'sd-0.007795577618316463, 32'sd0.07839111539725148, 32'sd0.0851043639591451, 32'sd0.05929992959757685, 32'sd0.06444923792765356, 32'sd-0.19734630209377643, 32'sd-0.11157424078936945, 32'sd-0.01886001620232604, 32'sd-0.0014646188076180915, 32'sd0.03811316749062808, 32'sd0.05701009918271594, 32'sd0.0482219090792121, 32'sd-0.010609425767966304, 32'sd-0.06265286302429006, 32'sd-0.06239655077442456, 32'sd0.017218244512019316, 32'sd-0.06936967083201631, 32'sd-0.023763290461659096, 32'sd-0.05545748610060101, 32'sd-0.05936232181586465, 32'sd-0.026486030428115037, 32'sd0.006350915087392301, 32'sd-1.6534944240240803e-125, 32'sd2.9829388243433703e-127, 32'sd3.505400370813364e-116, 32'sd6.696322788346376e-126, 32'sd-1.7834828255420749e-127, 32'sd8.577379605455161e-117, 32'sd-0.05291568543715928, 32'sd-0.05580385323015173, 32'sd-0.006020030445969645, 32'sd-7.939562599339718e-05, 32'sd-0.006259370506886354, 32'sd-0.009523360668803556, 32'sd0.07423529285081829, 32'sd0.08710425113422085, 32'sd-0.060905601367649435, 32'sd-0.11127362938721867, 32'sd-0.07516868912317895, 32'sd-0.014078247081568422, 32'sd-0.010926083112251201, 32'sd0.03266589045568206, 32'sd0.0005193431492018734, 32'sd-0.02380682189769024, 32'sd-0.020654828913131553, 32'sd-0.05476934578285693, 32'sd-0.04543771152764635, 32'sd-0.044065326860477066, 32'sd-9.120186651050562e-121, 32'sd9.701083158905304e-129, 32'sd1.1316590072423455e-127, 32'sd1.8187925070494797e-123},
        '{32'sd5.565710937203271e-122, 32'sd4.6643032370699846e-126, 32'sd6.891486098811294e-117, 32'sd-4.71594895814143e-118, 32'sd-2.700457550823855e-127, 32'sd-1.8032977174440098e-127, 32'sd-3.2362442101932486e-121, 32'sd1.5792903213284028e-123, 32'sd8.812609601243029e-127, 32'sd-3.0528642136066065e-120, 32'sd2.0504583276372675e-116, 32'sd3.4988098492723127e-119, 32'sd0.04755391367108931, 32'sd0.07488101782054099, 32'sd0.011616968335177792, 32'sd0.09846070304496041, 32'sd2.636342947448251e-129, 32'sd-3.168799547601808e-116, 32'sd-2.513062431597721e-124, 32'sd-3.2689730540363925e-120, 32'sd6.77190740347466e-124, 32'sd-3.2637316608124116e-125, 32'sd2.940193304297262e-115, 32'sd-1.1536879468279601e-129, 32'sd-1.6298402198666625e-119, 32'sd-1.5515813881983676e-121, 32'sd6.0424034377278876e-123, 32'sd-1.1402775754501992e-118, 32'sd1.049365766820998e-120, 32'sd1.0864324591679202e-115, 32'sd-1.9357976897075122e-127, 32'sd2.5254782981906772e-126, 32'sd-0.004351493464051609, 32'sd-0.020436034531324806, 32'sd-0.019474294148225928, 32'sd-0.04610193073536578, 32'sd0.020855318320054193, 32'sd0.0024286819865423775, 32'sd0.049894737018089046, 32'sd0.004559499018295905, 32'sd0.019181018878614006, 32'sd-0.021838696417189205, 32'sd-0.07848832773536099, 32'sd0.0071433540506269265, 32'sd-0.031458130508382386, 32'sd0.062401210989563964, 32'sd-0.002177315662928817, 32'sd0.08413953981573702, 32'sd0.05075477461756919, 32'sd0.01671927302156754, 32'sd0.04790535220130596, 32'sd-0.007780512131720433, 32'sd1.1512591472338438e-115, 32'sd6.6843796527573116e-124, 32'sd-1.7362992747142844e-125, 32'sd1.028857261210358e-121, 32'sd3.4296198350668726e-124, 32'sd4.749423451783227e-118, 32'sd0.044769926477589414, 32'sd-0.00534105608233312, 32'sd-0.013239454528428115, 32'sd-0.05861802187723131, 32'sd-0.023882069093534262, 32'sd-0.05694984283381161, 32'sd-0.01492166971906301, 32'sd-0.11620545748797544, 32'sd-0.03395188492436884, 32'sd0.0920959162778808, 32'sd0.09821635873033949, 32'sd0.03303326598822281, 32'sd0.0795247513763288, 32'sd0.05087822311060725, 32'sd0.11738104436252769, 32'sd0.09232692708645138, 32'sd0.019795823474422512, 32'sd0.0971178388201944, 32'sd0.0847317049201358, 32'sd0.12475460028049491, 32'sd0.10080580980315317, 32'sd0.019297836132364486, 32'sd0.057067467721099024, 32'sd-0.015129477698448213, 32'sd1.1059794238347827e-121, 32'sd-7.105549067747331e-124, 32'sd-5.7232542084472526e-120, 32'sd-9.158663539284233e-119, 32'sd0.005374194000605496, 32'sd-0.009435608524251845, 32'sd0.031058600197564866, 32'sd0.05762572266423309, 32'sd0.04739990889239757, 32'sd-0.08963767157340431, 32'sd-0.19591124324845002, 32'sd0.10295802358829301, 32'sd-0.012088505191569615, 32'sd0.041606653308036916, 32'sd-0.03535124674301642, 32'sd0.1119310950368815, 32'sd0.06052040054416766, 32'sd-0.103931871129032, 32'sd-0.010137223310660831, 32'sd-0.11755567121243223, 32'sd-0.039304877849007096, 32'sd-0.07324753211369292, 32'sd0.007016470200730444, 32'sd0.09266961441311754, 32'sd-0.006578900443916656, 32'sd0.06256235924687026, 32'sd0.03206188321980893, 32'sd0.027401326671276045, 32'sd-0.15088194580654757, 32'sd4.728435871527623e-123, 32'sd-1.4605542816435298e-124, 32'sd0.030062368247041532, 32'sd0.009695594915040824, 32'sd0.0177042866531418, 32'sd0.056284303980668735, 32'sd0.0426387182250609, 32'sd0.01899020127888563, 32'sd-0.014069872582621892, 32'sd-0.14361765788856032, 32'sd0.02981788672628184, 32'sd-0.04979840757294212, 32'sd-0.008439440171408866, 32'sd-0.02508888905343641, 32'sd-0.10724795614242437, 32'sd-0.20133583392163032, 32'sd-0.20054464426057694, 32'sd-0.011852468355644677, 32'sd0.01619385815723268, 32'sd0.01017203631797193, 32'sd-0.026122472863255197, 32'sd-0.07743417193883351, 32'sd0.021651062601833793, 32'sd-0.006113752982562886, 32'sd-0.05325745512166499, 32'sd-0.05542502894542169, 32'sd-0.10626494371435274, 32'sd-0.04404445389615285, 32'sd0.050237105731352275, 32'sd3.109664129392095e-119, 32'sd-0.016062050192938073, 32'sd-0.0798174344580319, 32'sd0.025235846617107455, 32'sd0.10054223798354565, 32'sd0.06912218726811671, 32'sd-0.04191222990575897, 32'sd-0.05854380851701721, 32'sd-0.030906516487531215, 32'sd-0.058206723846378094, 32'sd-0.018420692128684326, 32'sd0.026898717411662592, 32'sd-0.11450117994054959, 32'sd-0.09175010042119895, 32'sd-0.026055237716660185, 32'sd-0.055147867995250996, 32'sd-0.07791374358783369, 32'sd0.06368563568858815, 32'sd-0.033094112991306116, 32'sd0.13047382233465682, 32'sd-0.03106499124850653, 32'sd0.0766163507646696, 32'sd-0.0049638010602911994, 32'sd0.029969680138591234, 32'sd0.01279567010327534, 32'sd-0.1571006206182226, 32'sd-0.06292999033760993, 32'sd-0.0016181629687928682, 32'sd1.3690758195661635e-120, 32'sd-0.017740462989170435, 32'sd-0.06450362191593702, 32'sd0.010198395446872954, 32'sd-0.1359563086116962, 32'sd0.0012947289838929953, 32'sd0.08948017427031237, 32'sd0.028031833546594213, 32'sd-0.09161818330958084, 32'sd-0.07822123261788758, 32'sd-0.06617075777078321, 32'sd-0.038990247437793224, 32'sd-0.022511714069353997, 32'sd-0.07043627230896256, 32'sd-0.1614493824526402, 32'sd0.006868338920168354, 32'sd-0.04994361317658127, 32'sd-0.07334054363304235, 32'sd-0.015774589483437955, 32'sd0.0369234867521392, 32'sd0.1905673222942723, 32'sd0.14078922217377693, 32'sd0.055496784804561966, 32'sd-0.02816550816121948, 32'sd-0.057796081755500474, 32'sd-0.01622367225314465, 32'sd-0.04537387931637686, 32'sd0.1056625676727276, 32'sd0.027853761871489982, 32'sd0.016803788649050702, 32'sd0.010303194694086118, 32'sd-0.07940337785775467, 32'sd0.011703940673914243, 32'sd-0.06913917646945376, 32'sd0.0765904191537382, 32'sd-0.02791859791059846, 32'sd0.029816656529993553, 32'sd0.03317695375348238, 32'sd0.032424890540090796, 32'sd-0.006103049418947442, 32'sd0.03350216879062605, 32'sd-0.1049296456515757, 32'sd-0.16231452955078077, 32'sd0.11008413134318383, 32'sd0.07391343580898399, 32'sd0.02296053342620029, 32'sd0.06676345323013105, 32'sd0.010271398502343529, 32'sd0.13233599658673123, 32'sd0.07085056165936689, 32'sd0.0877176060737222, 32'sd0.06740976076541946, 32'sd-0.12867275681875895, 32'sd-0.02816362901076695, 32'sd0.10195345038613977, 32'sd0.0020559885601307767, 32'sd0.04414853398854009, 32'sd0.03688289888447116, 32'sd-0.05370830418052248, 32'sd-0.02140798489010591, 32'sd-0.037965358916702385, 32'sd-0.036196112750863596, 32'sd-0.05785432311278038, 32'sd0.06573874535032273, 32'sd0.04637873007788768, 32'sd0.09751855918815087, 32'sd0.12041919067537642, 32'sd0.18818980991393036, 32'sd0.0923850803724164, 32'sd-0.018307310203214886, 32'sd0.01844922313271295, 32'sd-0.09305191160738835, 32'sd0.04330631849518006, 32'sd0.000727793086589324, 32'sd0.005435955331009228, 32'sd-0.03641393095912062, 32'sd0.03817621787898598, 32'sd0.08900522256941731, 32'sd0.06007835362256074, 32'sd-0.15314595211577042, 32'sd-0.06994486932531059, 32'sd0.10858617676126349, 32'sd0.02675440989212739, 32'sd-0.032822619366692556, 32'sd0.03713251113052646, 32'sd0.037902220303936335, 32'sd-0.12842104850135114, 32'sd-0.020321736506725058, 32'sd-0.018089150225910032, 32'sd-0.13584764495002663, 32'sd-0.12644586998585852, 32'sd-0.09781574775186207, 32'sd-0.11360792762414076, 32'sd-0.13529598273621105, 32'sd0.1396052315236499, 32'sd0.22333419184200462, 32'sd0.03877030257068421, 32'sd0.022962882364246255, 32'sd-0.1489441430567886, 32'sd-0.058760830054931185, 32'sd-0.09843876297002695, 32'sd-0.04027197350044307, 32'sd-0.08499104949451913, 32'sd-0.10401988797306819, 32'sd0.027334115413576943, 32'sd0.019377751192651504, 32'sd-0.10507837897987635, 32'sd-0.08575222117125135, 32'sd-0.06631712515161965, 32'sd0.1747521475040608, 32'sd-0.05468553166381141, 32'sd-0.11287062212055268, 32'sd0.06370830702051207, 32'sd0.0915525631085902, 32'sd-0.00851991343904025, 32'sd-0.10920297580334092, 32'sd-0.014254389124745952, 32'sd-0.1103497098978655, 32'sd-0.1356200847143086, 32'sd-0.15109789988950068, 32'sd-0.11478791936747629, 32'sd-0.14277569180298058, 32'sd0.017270078197834604, 32'sd0.22412864532630578, 32'sd-0.01800872688721493, 32'sd-0.06315660608380913, 32'sd-0.16660364806623257, 32'sd-0.12662561050856147, 32'sd0.06580884779188592, 32'sd-0.02167151519816251, 32'sd-0.14001367758607025, 32'sd-0.1415859497058791, 32'sd-0.09828587968401319, 32'sd-0.127933777045731, 32'sd-0.10407985691235325, 32'sd-0.1965572626781674, 32'sd-0.03051358878910316, 32'sd0.057440796675074214, 32'sd0.03678500377800519, 32'sd-0.1177175799067912, 32'sd0.0849072500422423, 32'sd-0.011559767659573573, 32'sd-0.062328402216135004, 32'sd0.042500729261778177, 32'sd0.04608321619032256, 32'sd-0.1376031811886665, 32'sd-0.0001452012784124731, 32'sd-0.122894729384186, 32'sd-0.05470716150366928, 32'sd-0.12500344217678086, 32'sd-0.02800277918034473, 32'sd0.19446448703969613, 32'sd0.1564827821072261, 32'sd0.05159499427121929, 32'sd-0.1030271907431783, 32'sd-0.09244938345832152, 32'sd0.07456256710777713, 32'sd-0.019953886176576067, 32'sd-0.05063711773513682, 32'sd0.003357295097986841, 32'sd0.05631775430855287, 32'sd-0.036031414316233086, 32'sd-0.03532607457148755, 32'sd-0.07427013124911314, 32'sd-0.06905119226439081, 32'sd-0.02812459729561249, 32'sd0.04305387835409825, 32'sd-0.033827515463760637, 32'sd0.03145427472566038, 32'sd-0.031215179865812688, 32'sd0.06959018076942536, 32'sd0.04162817342612131, 32'sd-0.03298680841990144, 32'sd-0.09776286053193238, 32'sd-0.048024768611471536, 32'sd-0.10674849189312419, 32'sd-0.14224222713113288, 32'sd-0.12365345896281406, 32'sd-0.053592481697103775, 32'sd0.11650140286758137, 32'sd0.1206060816554645, 32'sd-0.09556584740698922, 32'sd-0.14107064792392462, 32'sd-0.0871912137580772, 32'sd-0.03690501371778169, 32'sd0.013285638107785918, 32'sd-0.005301972530870163, 32'sd-0.05893862821921113, 32'sd0.0997501097633388, 32'sd0.041869686498439564, 32'sd0.036777262288770374, 32'sd-0.0838624762542804, 32'sd-0.0699940032081393, 32'sd-0.029215328667106764, 32'sd0.016747686145456547, 32'sd0.0072078808429417544, 32'sd-0.020485799596829318, 32'sd0.0499397238464582, 32'sd-0.03540968325422086, 32'sd-0.05016523115961637, 32'sd0.01818045564556106, 32'sd0.0385761828578263, 32'sd-0.0008489360678477199, 32'sd-0.07383184225340389, 32'sd-0.13691555321081778, 32'sd-0.0889709175536113, 32'sd0.09827811631087083, 32'sd0.010693439398582643, 32'sd-0.057858686194364746, 32'sd-0.1445058983222382, 32'sd-0.1676142870498175, 32'sd-0.019578557848780563, 32'sd0.025480927369503522, 32'sd0.007958196244415754, 32'sd0.05008945647458168, 32'sd0.12905112092952914, 32'sd0.042169858137292036, 32'sd0.059854473247923416, 32'sd0.11212537126031945, 32'sd-0.03434913058201128, 32'sd-0.1831032078368704, 32'sd-0.07092302235272775, 32'sd0.009385769139307111, 32'sd-0.0023693297606807557, 32'sd0.04609352480656233, 32'sd0.04808760190912151, 32'sd0.047850433811532686, 32'sd-0.019479154304231396, 32'sd0.018489530291071147, 32'sd0.004719959598247275, 32'sd-0.12360359181764076, 32'sd0.0011887348086397967, 32'sd-0.13862165898674353, 32'sd0.028615810418909197, 32'sd0.15421083001707048, 32'sd0.09709703608008934, 32'sd-0.02522918781294496, 32'sd-0.007365314797243943, 32'sd-0.07303002922881949, 32'sd0.0949263533881805, 32'sd0.03126936524129188, 32'sd-0.13572699214388026, 32'sd0.10624707660099315, 32'sd0.05534625513990501, 32'sd0.1950833963942204, 32'sd0.20039143260808606, 32'sd0.10234654135693629, 32'sd-0.07297992557255817, 32'sd-0.12050983570550672, 32'sd0.05626362425979907, 32'sd0.03704267530884749, 32'sd0.04293401974294685, 32'sd-0.04299772677303529, 32'sd0.016095348148426437, 32'sd-0.0232138387167823, 32'sd-0.04120161445205658, 32'sd-0.14459504050807775, 32'sd-0.14563565208162343, 32'sd-0.09982976552189866, 32'sd-0.04170340596413905, 32'sd-0.03465308625674628, 32'sd0.034448527203879455, 32'sd0.15824782407286275, 32'sd0.07823943888912907, 32'sd-0.03885971775069717, 32'sd-0.029945879764374232, 32'sd0.06738968591595978, 32'sd0.08671005442511424, 32'sd0.052681444683963324, 32'sd0.0741307444332404, 32'sd0.08158563915674646, 32'sd0.09806020745844621, 32'sd0.045976578677436895, 32'sd0.07079039276267467, 32'sd-0.09474676747975165, 32'sd-0.04515496874988718, 32'sd-0.15610959237986044, 32'sd0.011967994441056635, 32'sd0.02853789080531952, 32'sd-0.034979366075798414, 32'sd-0.0009562170003916229, 32'sd0.02817167783132952, 32'sd-0.13495046260036248, 32'sd-0.09007482376426346, 32'sd-0.0920989007160517, 32'sd-0.014538234132611638, 32'sd-0.09806395993708132, 32'sd-0.10735393833258755, 32'sd0.019624932199902394, 32'sd0.07809846739081477, 32'sd-0.04654967303278388, 32'sd0.02065120937240194, 32'sd-0.02913115875968198, 32'sd-0.0314397662661274, 32'sd-0.03668616589959147, 32'sd0.03173020729566609, 32'sd0.04531265342095835, 32'sd0.011113317337630692, 32'sd0.011914193237952831, 32'sd-0.12042081976664044, 32'sd-0.06307243269397474, 32'sd-0.08911288012618283, 32'sd-0.006535620974258286, 32'sd-0.15780558078754173, 32'sd-0.047269266808292694, 32'sd0.059195026152558616, 32'sd0.07290416149638052, 32'sd0.012604353307405274, 32'sd-9.828849369696489e-123, 32'sd0.028075547603123058, 32'sd-0.0767385957113596, 32'sd0.0060539510494165664, 32'sd0.06692609548928492, 32'sd0.05878854644646393, 32'sd-0.16819582397812655, 32'sd-0.08955278143219678, 32'sd0.06429544861299796, 32'sd-0.016228039125413693, 32'sd0.1201492235156722, 32'sd-0.025835271756959703, 32'sd-0.10821330133175533, 32'sd-0.08184754173904957, 32'sd0.07691664276737865, 32'sd0.001444423619314037, 32'sd0.09573172461356476, 32'sd-0.09189575425773329, 32'sd-0.02696962538268, 32'sd-0.11176520606143729, 32'sd-0.04658502044980673, 32'sd-0.11529715278440017, 32'sd-0.09381758068092924, 32'sd-0.1035291239736415, 32'sd-0.16277018494537848, 32'sd0.028171935308450916, 32'sd-0.05485230696556747, 32'sd-0.02483779377143298, 32'sd-0.03737103513228658, 32'sd0.03778314821627247, 32'sd0.03582975490938023, 32'sd-0.022063021965314848, 32'sd0.01582366263352426, 32'sd-0.13362682616368, 32'sd-0.1242605368338882, 32'sd-0.04126253845954917, 32'sd0.06860224809506472, 32'sd0.04102627008152757, 32'sd0.02067450053823699, 32'sd0.06291223487743865, 32'sd0.023919786050343773, 32'sd0.029648537635435932, 32'sd0.09499317938141873, 32'sd0.12874383209702664, 32'sd-0.04369362109376483, 32'sd-0.03706255368388782, 32'sd-0.0034424276111691254, 32'sd0.0007672529206188427, 32'sd-0.16439419986893156, 32'sd-0.132139158385011, 32'sd-0.05809537343043536, 32'sd-0.049346686747485526, 32'sd-0.08727942377418442, 32'sd-0.10703239851239887, 32'sd-0.1355868735550072, 32'sd0.03838481624728258, 32'sd0.01154130064299484, 32'sd-0.04319616968151127, 32'sd0.03037176108198672, 32'sd-0.05867853498365445, 32'sd0.021508914648879045, 32'sd0.008408950023072905, 32'sd-0.12375711718212891, 32'sd-0.12046618293995173, 32'sd0.06362916965853578, 32'sd0.06023987294055667, 32'sd0.1533085821855024, 32'sd0.08437053107410572, 32'sd0.056496443717004796, 32'sd-0.10448414720936242, 32'sd0.052127747322680835, 32'sd-0.02107326146256157, 32'sd-0.055244605714926044, 32'sd-0.1916124031060607, 32'sd-0.03285168240045358, 32'sd0.08293022079139062, 32'sd-0.020137206406400165, 32'sd-0.10107270072437291, 32'sd-0.02378741355186932, 32'sd0.07370122062047495, 32'sd0.07541518707633982, 32'sd-0.019926384253366607, 32'sd-0.05857070666888435, 32'sd0.09069106464185836, 32'sd-6.114803709022872e-126, 32'sd-0.06932209186088872, 32'sd0.05535056796612322, 32'sd-0.1147834144897355, 32'sd-0.08774477522453818, 32'sd-0.1546435436708715, 32'sd-0.03538187291351178, 32'sd-0.13810057401809012, 32'sd-0.06152563614935572, 32'sd0.04783763452367165, 32'sd0.1436518727197001, 32'sd0.13879768485720542, 32'sd0.05432890772545741, 32'sd-0.15272526040562312, 32'sd-0.060333269060001776, 32'sd-0.14184755404652252, 32'sd-0.12346333780776918, 32'sd-0.12168890939268359, 32'sd-0.0293874134716693, 32'sd-0.04528903954611077, 32'sd-0.10614306119733605, 32'sd-0.0821816761498556, 32'sd-0.028370923601968065, 32'sd0.07001736640474683, 32'sd0.06972883502320233, 32'sd-0.004413544103137574, 32'sd-0.02935092734374403, 32'sd0.051342823286339496, 32'sd-0.010787190259605861, 32'sd0.032843650593019184, 32'sd0.015601371719854734, 32'sd-0.03500358038359586, 32'sd-0.11220131926693105, 32'sd-0.18231195861547145, 32'sd-0.20376073797572195, 32'sd-0.15059881944405984, 32'sd-0.07042145136167334, 32'sd-0.05119553216673852, 32'sd-0.06011023739124114, 32'sd0.02819076700733539, 32'sd0.10209749324860963, 32'sd0.06848484553869948, 32'sd-0.06144543791890609, 32'sd-0.10374494077633195, 32'sd-0.09965021139874256, 32'sd-0.05463387639972374, 32'sd-0.10236509204855912, 32'sd-0.14235232053320665, 32'sd-0.2105262393826825, 32'sd-0.014818048405260943, 32'sd0.1265477626177892, 32'sd0.14410147510268997, 32'sd0.1263647076289817, 32'sd-0.004050169259412346, 32'sd0.0017108020119816333, 32'sd0.031463685073788016, 32'sd-0.05882446438426988, 32'sd-0.00502109099082939, 32'sd0.03418484773905625, 32'sd-0.03483922292387203, 32'sd-0.11108139417131543, 32'sd-0.04363320190938525, 32'sd-0.12786999131445012, 32'sd0.016994524867393803, 32'sd-0.07657749420062764, 32'sd0.023265966463635032, 32'sd-0.04013527892657752, 32'sd-0.06685294794277033, 32'sd0.10693699833594464, 32'sd0.1831430160828288, 32'sd0.0924918070253682, 32'sd0.088378672302302, 32'sd5.384055789619733e-06, 32'sd-0.1169851096193286, 32'sd-0.06703435255894796, 32'sd-0.06182634699247492, 32'sd-0.10746035193884716, 32'sd-0.015179678227096996, 32'sd0.06673829235323066, 32'sd-0.02922339540046644, 32'sd-0.04465541774141134, 32'sd0.0811576811669571, 32'sd0.10507884094670518, 32'sd-0.020530176777283863, 32'sd2.3413942573913317e-124, 32'sd0.051458981118971125, 32'sd-0.024491398762406073, 32'sd0.033656752026515475, 32'sd-0.19196938643512293, 32'sd-0.11932593902001229, 32'sd-0.06473685797987756, 32'sd-0.034797560823716385, 32'sd0.09116023108259622, 32'sd0.11109766310792692, 32'sd-0.008992658745270554, 32'sd-0.07363456390798348, 32'sd0.09296742464781792, 32'sd0.12733470233814212, 32'sd0.0250805126658864, 32'sd-0.1081805674987964, 32'sd0.031624028671327055, 32'sd-0.0330078671473775, 32'sd-0.06919321365664582, 32'sd-0.08259062488401961, 32'sd-0.05507374595705554, 32'sd0.06695273454244766, 32'sd0.08185164170418663, 32'sd0.06054756196019599, 32'sd-0.06560458301834035, 32'sd0.06379014066123144, 32'sd-0.011153479554135686, 32'sd1.3387143906984537e-122, 32'sd-8.923760934687827e-125, 32'sd7.224979890827148e-119, 32'sd-0.0030576261701913236, 32'sd0.03300131003537172, 32'sd-0.11301589844103124, 32'sd-0.11267866034500928, 32'sd-0.04776865718324438, 32'sd-0.06725002683505821, 32'sd-0.1231367449422576, 32'sd-0.1355484314902317, 32'sd-0.036373199198307914, 32'sd-0.0019663333250446286, 32'sd0.11095568201354805, 32'sd0.027141239944090442, 32'sd-0.027164958767035684, 32'sd0.03647600785253713, 32'sd0.11888490805426996, 32'sd-0.004520559717421068, 32'sd-0.15090114569764568, 32'sd-0.10747249100617835, 32'sd-0.09878989957238961, 32'sd-0.02175250307092274, 32'sd-0.05864791739597196, 32'sd-0.09796126480085222, 32'sd-0.04427375397388427, 32'sd-0.038729430221083334, 32'sd0.06845833104509758, 32'sd3.341017787072968e-120, 32'sd1.3835264547336366e-115, 32'sd-4.843653876208434e-119, 32'sd-0.010873397329012368, 32'sd-0.00492391544681011, 32'sd-0.008693923467704928, 32'sd0.058599361956070004, 32'sd-0.03922199990347375, 32'sd0.022169808976239137, 32'sd-0.146136331187676, 32'sd-0.09281922544966223, 32'sd-0.030294086994360387, 32'sd-0.04083230311833815, 32'sd0.09942027690527123, 32'sd-0.030457699984813486, 32'sd0.08840030302198612, 32'sd0.24410548833133203, 32'sd-0.001054506827279657, 32'sd-0.05579592537498781, 32'sd0.009559048121065955, 32'sd-0.0542634108062402, 32'sd-0.0859551104722319, 32'sd-0.11078336663128784, 32'sd-0.08544835129150649, 32'sd0.0313079237470211, 32'sd0.07735848426877433, 32'sd-0.006057360039147915, 32'sd0.01626783691944551, 32'sd3.253393164786763e-126, 32'sd6.043950843776001e-121, 32'sd2.812889668889427e-123, 32'sd5.644545777151549e-127, 32'sd0.02768155417879259, 32'sd-0.07570173105739077, 32'sd-0.10215998703148363, 32'sd0.026682778509701653, 32'sd0.026749683766137188, 32'sd0.11330155005519842, 32'sd0.027898417443610043, 32'sd0.030750804854117023, 32'sd-0.07790536995903186, 32'sd-0.04069246945929762, 32'sd0.11656808615519013, 32'sd-0.056315182711014426, 32'sd-0.03984311588439225, 32'sd-0.02365737999368799, 32'sd-0.03897312228510798, 32'sd0.00933031172532422, 32'sd-0.025509148030733512, 32'sd0.03797542612041807, 32'sd-0.04785474371139358, 32'sd-0.05650161966684992, 32'sd0.011526063897433521, 32'sd0.018628708460034744, 32'sd0.062461288949499795, 32'sd2.9828592057756745e-122, 32'sd2.4513727576401584e-125, 32'sd-3.417556234501449e-124, 32'sd3.8281853691431873e-119, 32'sd-1.0614416870587104e-121, 32'sd-1.563403034717627e-123, 32'sd-0.01719501344454109, 32'sd-0.030146047644983246, 32'sd0.03260330963008868, 32'sd-0.013769774494496958, 32'sd0.02096742197099031, 32'sd0.030619943436078836, 32'sd-0.03829780795970126, 32'sd-0.029173329340390963, 32'sd-0.05456473149665278, 32'sd0.060083640068542374, 32'sd-0.016395625228754266, 32'sd0.012125228119769484, 32'sd-0.03179025185688224, 32'sd0.048399350458994295, 32'sd0.03314841189636385, 32'sd0.03919071782400508, 32'sd-0.014493307180445935, 32'sd-0.010485215025257958, 32'sd-0.0348093046984875, 32'sd-0.015334654718068282, 32'sd7.53213681851393e-127, 32'sd2.3200107565000463e-120, 32'sd-8.61996947369413e-121, 32'sd8.808593674197157e-116},
        '{32'sd2.552740678522959e-122, 32'sd2.8896644952480505e-123, 32'sd6.116281479377847e-115, 32'sd-4.1523789317692275e-115, 32'sd5.241939180215187e-118, 32'sd1.3350993579019754e-122, 32'sd-1.2770585345609418e-115, 32'sd-3.501863447096834e-130, 32'sd4.852975799681466e-122, 32'sd6.999525982796195e-119, 32'sd5.948177528603374e-119, 32'sd-8.78173669562027e-127, 32'sd-0.11501769965621725, 32'sd-0.04404294483631126, 32'sd-0.04587378172494238, 32'sd-0.0036915004449179886, 32'sd-8.909401532960828e-122, 32'sd3.1561802568901057e-125, 32'sd2.7312582757923764e-121, 32'sd2.932988654057601e-121, 32'sd9.873796658734089e-123, 32'sd1.5802803308932992e-116, 32'sd-2.2760210467796144e-118, 32'sd1.529488590972231e-127, 32'sd3.800883974402045e-122, 32'sd-1.8157008618500155e-123, 32'sd2.9173610422950663e-122, 32'sd-1.5258802013055257e-117, 32'sd-1.3858462987408035e-117, 32'sd-5.865706706449106e-125, 32'sd-5.207158317120089e-124, 32'sd1.3725947773710494e-124, 32'sd-0.00010806635730285257, 32'sd0.024222529910665855, 32'sd0.04926010765510998, 32'sd-0.08167439060121559, 32'sd-0.03290129695554694, 32'sd-0.04228842244625906, 32'sd0.019180466476913918, 32'sd0.0711514638314195, 32'sd-0.06552432186372262, 32'sd-0.0554126367751031, 32'sd0.03695060364242104, 32'sd0.10832335239233505, 32'sd-0.012978142872218722, 32'sd-0.004469462512996026, 32'sd0.07520535757940833, 32'sd0.03587903659189075, 32'sd-0.04786944638890066, 32'sd0.05839326469812966, 32'sd0.015647028446962745, 32'sd0.0013672269786700719, 32'sd-2.676354064603722e-124, 32'sd-1.9284329829311183e-129, 32'sd5.072271814720591e-120, 32'sd1.2603682632702723e-125, 32'sd-6.2356344586772e-126, 32'sd2.684134003202732e-119, 32'sd-0.005921783726362852, 32'sd-0.008127905269493722, 32'sd-0.022935061585676698, 32'sd-0.0020202619281715585, 32'sd-0.03706457395254638, 32'sd-0.08652225131226084, 32'sd-0.0348114711071082, 32'sd-0.07520358070180064, 32'sd0.04179515097791124, 32'sd-0.07886911521035643, 32'sd-0.006140724024827924, 32'sd-0.15899317090976442, 32'sd-0.07511796867061571, 32'sd0.1332714608400926, 32'sd0.07830102512449695, 32'sd-0.03572274854439054, 32'sd-0.035414876503801464, 32'sd0.07498428325977259, 32'sd-0.06316975919308244, 32'sd-0.007856986111839222, 32'sd0.014498798766225509, 32'sd0.034500368363687785, 32'sd0.03995658001597759, 32'sd-0.012260296756166062, 32'sd-8.779299073450166e-127, 32'sd8.544827300559477e-117, 32'sd1.4792605259998017e-123, 32'sd8.826392765093993e-127, 32'sd0.052520197708945046, 32'sd-0.002269711706095546, 32'sd0.02980330056999574, 32'sd0.014105120850543804, 32'sd-0.014906016520102322, 32'sd-0.13635629692576784, 32'sd-0.05806979852493247, 32'sd0.05358204363730068, 32'sd0.019480622177947063, 32'sd0.03436737096734149, 32'sd-0.03648208812634099, 32'sd0.011039569539211418, 32'sd0.003724861547777905, 32'sd0.06275899117112864, 32'sd-0.15724634199646237, 32'sd-0.19028935192516727, 32'sd-0.11480168063785033, 32'sd-0.1018107773460773, 32'sd-0.08176890159827657, 32'sd0.0377195935569901, 32'sd0.04631910599025428, 32'sd0.013126017332009519, 32'sd-0.08523540338570275, 32'sd-0.04279819049553057, 32'sd-0.013982339762613458, 32'sd8.566268095033752e-119, 32'sd-8.085544608712277e-117, 32'sd-0.0027402938700745233, 32'sd0.05318769983031721, 32'sd0.06942221033499742, 32'sd-0.03673267703472995, 32'sd-0.03983586714223941, 32'sd-0.1566693437260592, 32'sd0.005921776284739637, 32'sd0.0023020974781168485, 32'sd0.09781250733050391, 32'sd0.0430508267355491, 32'sd0.03800428417284469, 32'sd-0.1525777231792553, 32'sd-0.18490960037721027, 32'sd0.046080767036212014, 32'sd0.03898962304413156, 32'sd0.054618379182124234, 32'sd0.08948977972184667, 32'sd-0.06720972173668141, 32'sd-0.06606796197440669, 32'sd-0.12858675534222502, 32'sd-0.1065480563207159, 32'sd-0.13594670348750648, 32'sd-0.015699985962438302, 32'sd-0.11849520314278869, 32'sd-0.028714830241869747, 32'sd-0.03220706394721016, 32'sd-0.007605824067485099, 32'sd3.6876341731277595e-128, 32'sd-0.010934259526299369, 32'sd-0.0492727690054974, 32'sd-0.03885830907917881, 32'sd-0.07913690834650393, 32'sd-0.04857530113406564, 32'sd0.020743778094599617, 32'sd0.11189613192488286, 32'sd-0.06794753006920637, 32'sd0.02122648183741097, 32'sd0.05534100251257071, 32'sd0.08331062949173175, 32'sd0.10445149487469647, 32'sd0.09608138946713077, 32'sd0.21887287095291647, 32'sd-0.06551980780809778, 32'sd-0.05157897404372139, 32'sd-0.0151048009091822, 32'sd-0.19121386518989253, 32'sd-0.11562205374929628, 32'sd0.03589602238013323, 32'sd0.1318624958979245, 32'sd-0.01821465797807556, 32'sd-0.15572233071296238, 32'sd-0.06453189663598322, 32'sd-0.043273436651879285, 32'sd0.05875823076168885, 32'sd-0.0670070442288195, 32'sd-2.4436414417207012e-116, 32'sd-0.01763713629267993, 32'sd-0.030364479107451815, 32'sd0.0765044016333151, 32'sd-0.06599102019661535, 32'sd0.1245843703960127, 32'sd0.1379403197195924, 32'sd0.0959773817013923, 32'sd0.012804277649303138, 32'sd-0.01411340551957204, 32'sd0.11550999038489519, 32'sd0.08576235495726886, 32'sd0.24085080826995167, 32'sd0.06821509819611939, 32'sd-0.06502197352507746, 32'sd-0.031110389819961257, 32'sd-0.2461606335459254, 32'sd-0.1496750254870536, 32'sd-0.15051760703002606, 32'sd-0.05150381784956872, 32'sd-0.030195186776755773, 32'sd0.03782036348183466, 32'sd-0.08650325349339982, 32'sd-0.009396065224715078, 32'sd-0.033767251407940596, 32'sd0.07508040385473437, 32'sd0.07299643090241335, 32'sd0.012622152365417284, 32'sd-0.007893685178254669, 32'sd0.04114326382605467, 32'sd-0.044345930105205586, 32'sd0.09461509373418274, 32'sd-0.095834331211381, 32'sd0.04108486880881548, 32'sd0.13150773585670564, 32'sd0.05882939324155382, 32'sd0.06758127648817862, 32'sd0.026053372492760473, 32'sd0.04741432793852299, 32'sd0.052342967109028395, 32'sd0.05945471030025652, 32'sd-0.028512531789641887, 32'sd-0.00898482220405344, 32'sd-0.11075221245468751, 32'sd-0.02409329932100451, 32'sd-0.04854576590916811, 32'sd-0.05413458042573443, 32'sd0.07424335447169333, 32'sd0.07521585063998143, 32'sd0.15062433041548995, 32'sd0.07329826610299361, 32'sd-0.0769122586775713, 32'sd-0.08242144434958144, 32'sd0.03976808956062204, 32'sd-0.08879623975836497, 32'sd0.06545543950281832, 32'sd-0.029156299376050274, 32'sd-0.055578448630250424, 32'sd0.007105865716527427, 32'sd-0.06381047663737616, 32'sd0.012245768554218344, 32'sd0.09061300633475536, 32'sd0.1212943725476533, 32'sd0.17573353353899046, 32'sd0.09769166190968505, 32'sd0.03678754060839801, 32'sd0.13603928852371433, 32'sd0.03752376144579149, 32'sd0.10807048753873108, 32'sd0.010087451388874976, 32'sd-0.034031945378227714, 32'sd-0.009305793368937868, 32'sd0.06358711321415915, 32'sd0.0660918456500357, 32'sd0.0494294541073629, 32'sd0.17283558291264692, 32'sd0.1643386884347562, 32'sd0.09431574620772995, 32'sd0.15607484581172001, 32'sd0.13815765957655815, 32'sd0.09091767970993281, 32'sd0.08366061776350629, 32'sd0.04006972143780492, 32'sd0.09821986803527737, 32'sd0.011633401135720844, 32'sd-0.053722509907637224, 32'sd0.03158616486803122, 32'sd-0.0637187493316682, 32'sd0.042720731800250045, 32'sd-0.015424544731375807, 32'sd0.08254949905982654, 32'sd0.07560625593556498, 32'sd-0.02718831850622176, 32'sd-0.02082941493523574, 32'sd0.10943810952469613, 32'sd0.20134833164231686, 32'sd0.07122797815326398, 32'sd0.10702855763418832, 32'sd0.08815769277115885, 32'sd0.12450964924161476, 32'sd0.1047655769954376, 32'sd0.06537593041073603, 32'sd0.17676188482472305, 32'sd0.17159851837315396, 32'sd0.26677174850070384, 32'sd0.1401115224274508, 32'sd0.18638980113633788, 32'sd0.03145049224704434, 32'sd0.11156379517725434, 32'sd0.11866922984612051, 32'sd0.05323900283670991, 32'sd0.07355763829452495, 32'sd-0.02482712307353513, 32'sd-0.038545268391183184, 32'sd0.0234629865602095, 32'sd-0.1422340454971765, 32'sd-0.024182337585156748, 32'sd-0.053300330489549734, 32'sd0.002685013710356654, 32'sd-0.017941523669986702, 32'sd0.00688228987536634, 32'sd-0.1065411198433982, 32'sd0.03671802084805901, 32'sd0.09678881175453191, 32'sd0.05237343642471005, 32'sd0.053212784175461936, 32'sd0.08626281762673808, 32'sd0.17659925518323258, 32'sd-0.00822148179211089, 32'sd0.0058741636876344285, 32'sd0.2555149385426638, 32'sd0.2515388447646015, 32'sd0.1649726142862276, 32'sd0.15107556648316503, 32'sd0.10050885995046208, 32'sd-0.00039069659182154354, 32'sd0.18679014788800016, 32'sd0.10136402964815039, 32'sd-0.028161273639135054, 32'sd0.05512250130100932, 32'sd0.012937503868764914, 32'sd-0.039112236401037156, 32'sd0.015235016866026995, 32'sd-0.08274488506371849, 32'sd-0.059308810075018745, 32'sd0.05719690115761685, 32'sd0.061581852770743156, 32'sd0.08532257720316283, 32'sd-0.08820109061219963, 32'sd-0.11168126390567745, 32'sd-0.06757753242804075, 32'sd0.06165262906531667, 32'sd-0.2107669273773972, 32'sd-0.12201660434204063, 32'sd-0.0743700823855095, 32'sd-0.002479634042863442, 32'sd-0.040192870023936796, 32'sd-0.033023965203939805, 32'sd0.05901748872720132, 32'sd0.05964338539514533, 32'sd0.0712688610212793, 32'sd0.05106715623492289, 32'sd0.03778933849253004, 32'sd-0.06031379071434179, 32'sd0.03210227937023233, 32'sd0.014274813030693759, 32'sd0.0858141435292753, 32'sd0.07709726232331798, 32'sd0.026153175820962618, 32'sd0.03687428100133123, 32'sd0.02858134131610375, 32'sd-0.007151017453685681, 32'sd-0.04646255429007257, 32'sd-0.06724755264229455, 32'sd-0.07081078524384725, 32'sd0.12103128998119149, 32'sd0.12332587695401168, 32'sd0.08061718106256156, 32'sd-0.1342472320543697, 32'sd-0.02060276280897489, 32'sd-0.0930055638914004, 32'sd-0.09192135938333723, 32'sd-0.12107149749045487, 32'sd-0.10404847818885014, 32'sd-0.188520608165323, 32'sd0.003779062278407493, 32'sd-0.11793223730197908, 32'sd-0.0453029065230623, 32'sd-0.09748990239506852, 32'sd0.06772673019024224, 32'sd-0.00671718208703262, 32'sd-0.09225387880309334, 32'sd-0.05094170642225945, 32'sd0.12598109354408066, 32'sd-0.021136016836797757, 32'sd-0.060709849369161524, 32'sd-0.022697884900072567, 32'sd0.07854523870513196, 32'sd0.10100942581593371, 32'sd0.018681126121085, 32'sd-0.06364374725350003, 32'sd-0.12520580045710097, 32'sd-0.07211923022836533, 32'sd0.04484861420570949, 32'sd0.16091400594882413, 32'sd0.02065409526036589, 32'sd0.06673046857846104, 32'sd-0.06237009833006348, 32'sd-0.1115323814887306, 32'sd-0.16907383162360468, 32'sd-0.15924043331721097, 32'sd-0.17524224688608747, 32'sd-0.04387306767796073, 32'sd-0.020089941143022216, 32'sd-0.14419452961037318, 32'sd-0.23862899194200743, 32'sd-0.09120045944541595, 32'sd-0.043359309187912885, 32'sd-0.08248219783302782, 32'sd-0.09618387819720578, 32'sd-0.027743981543489074, 32'sd0.12442648724392778, 32'sd-0.026337777956719845, 32'sd-0.01517436497203564, 32'sd0.11414253265869373, 32'sd0.03767976947155942, 32'sd-0.08081805076468054, 32'sd0.01671769802492036, 32'sd-0.1176794375378392, 32'sd-0.17337380789500062, 32'sd-0.10590355554091481, 32'sd-0.07533240273282185, 32'sd0.033167645728963045, 32'sd0.022687589690569027, 32'sd0.1035493095504078, 32'sd0.004408801813588647, 32'sd-0.08190898407500848, 32'sd-0.1788117939441178, 32'sd-0.1519901676207027, 32'sd-0.1447981851833391, 32'sd-0.14965935796903765, 32'sd-0.04192827676016475, 32'sd-0.18292748276457216, 32'sd-0.23720562603123158, 32'sd-0.11440946236560448, 32'sd-0.025853160621146416, 32'sd-0.07033294408419032, 32'sd0.006947540914222696, 32'sd-0.13506650075437715, 32'sd-0.11751682600546141, 32'sd-0.08447439355926159, 32'sd0.03703076019674506, 32'sd-0.007425241639530506, 32'sd-0.10948395240082404, 32'sd-0.12642428495077626, 32'sd0.016584345400663128, 32'sd0.05652782467050218, 32'sd-0.09923567028353761, 32'sd0.0097844031275062, 32'sd0.02891099070611772, 32'sd-0.011019173432174923, 32'sd0.08913343393029152, 32'sd0.08714796619218208, 32'sd-0.010549091118422787, 32'sd-0.1376713891214605, 32'sd-0.07990620553029948, 32'sd-0.22198276998552077, 32'sd-0.11370618724014132, 32'sd-0.21505059108896915, 32'sd-0.0942370627549099, 32'sd-0.16042243390621574, 32'sd-0.1769269683085386, 32'sd-0.16781756770583492, 32'sd0.056687640857698604, 32'sd-0.1340720052980387, 32'sd0.06392007698734326, 32'sd-0.0915021923448929, 32'sd0.0012943815543280956, 32'sd-0.04214851858908926, 32'sd0.0006109492025431707, 32'sd0.03761731743175346, 32'sd0.02927001490357615, 32'sd-0.10095689584754904, 32'sd0.05348726839869841, 32'sd0.029335772032432796, 32'sd-0.01780784505529805, 32'sd0.04020569357629849, 32'sd-0.011805406763552415, 32'sd0.031166875414948964, 32'sd0.1967134986415525, 32'sd0.03930559570965919, 32'sd-0.07525611717627322, 32'sd-0.2287034257825049, 32'sd-0.1579454808422401, 32'sd-0.06339101821071719, 32'sd-0.051388661712280535, 32'sd-0.095686966194693, 32'sd0.05858785862403154, 32'sd-0.025282583912277067, 32'sd-0.006092640739107278, 32'sd-0.10122713246084016, 32'sd0.040061180961153506, 32'sd-0.010235172088649037, 32'sd0.09613834236946388, 32'sd-0.06056943965992099, 32'sd0.1559219867492713, 32'sd-0.09180595621079023, 32'sd0.00939235749175642, 32'sd7.138162458687607e-123, 32'sd0.056675190864535235, 32'sd0.05529003316318173, 32'sd0.002947119487487144, 32'sd0.0736673037707264, 32'sd0.09363209219734525, 32'sd0.05622074591206842, 32'sd0.11460682678792125, 32'sd0.17592978331822384, 32'sd0.1812161839068107, 32'sd0.06563029260377483, 32'sd-0.057446470091782074, 32'sd-0.09679505102061975, 32'sd-0.09541104128690645, 32'sd-0.0674396120586115, 32'sd0.023737280495628024, 32'sd0.08543091028825234, 32'sd0.03933552860984447, 32'sd0.015359946762275404, 32'sd-0.08440703371934118, 32'sd0.00714322402789603, 32'sd-0.10014421587713208, 32'sd-0.08230254392964875, 32'sd-0.05330860578296453, 32'sd0.0007731334986986969, 32'sd-0.07907273302745581, 32'sd0.00798509433096603, 32'sd0.04173795604950731, 32'sd-0.023555753800061873, 32'sd-0.028530651757441225, 32'sd0.013656597846871883, 32'sd-0.0815413961041519, 32'sd-0.052155106422434004, 32'sd0.03899417264570166, 32'sd0.10524228507792033, 32'sd0.14873982186950976, 32'sd0.07151649073914154, 32'sd-0.015967560568664836, 32'sd0.06187846017369005, 32'sd-0.023556406605761943, 32'sd-0.06404271849767648, 32'sd0.10757219931073497, 32'sd0.0813954326592436, 32'sd0.025408273710204772, 32'sd0.05715516752310008, 32'sd0.01972228896577958, 32'sd-0.016893298426408104, 32'sd-0.07005077347191725, 32'sd-0.03951441561659382, 32'sd0.0454197871814592, 32'sd-0.08215532470589193, 32'sd0.0668730784168808, 32'sd-0.03148179950509151, 32'sd-0.05818840478481364, 32'sd0.02856087486232303, 32'sd0.04383281643544752, 32'sd0.04630581117998421, 32'sd-0.06834751516854065, 32'sd-0.08823309024154204, 32'sd-0.06861882824921871, 32'sd0.09603546286562231, 32'sd-0.030589942961160063, 32'sd0.07304340500740025, 32'sd0.07896149208362828, 32'sd-0.022127660423347996, 32'sd0.022121372479733312, 32'sd-0.1284985576269604, 32'sd-0.07926006519677803, 32'sd0.06956083371648489, 32'sd0.07152226796275957, 32'sd0.027116110457799648, 32'sd0.02257696912819382, 32'sd0.016972422027913544, 32'sd0.001180044650220009, 32'sd0.0020605056910694163, 32'sd-0.021153748193964296, 32'sd-0.09078372727767378, 32'sd-0.025374195145150283, 32'sd-0.03545088201388352, 32'sd-0.06517042419034283, 32'sd0.07466899953072856, 32'sd-0.05478411350167864, 32'sd0.028694255800338138, 32'sd0.109033039134349, 32'sd2.5344027271073623e-128, 32'sd0.003001228111139917, 32'sd0.09923535853366891, 32'sd0.0012503677651584005, 32'sd-0.0574309313047064, 32'sd0.04169157682205978, 32'sd-0.049354378161465276, 32'sd0.06813809975689122, 32'sd-0.0671128668815417, 32'sd-0.12281006023379895, 32'sd0.037336050566116594, 32'sd0.024118569072875084, 32'sd0.12693879958259122, 32'sd0.07985286940716055, 32'sd0.12702659460032054, 32'sd0.14757000743153043, 32'sd0.03500802843600827, 32'sd-0.11457205300725713, 32'sd-0.11933898852882507, 32'sd-0.12271653244877435, 32'sd-0.045056779573633285, 32'sd-0.05042665215440673, 32'sd-0.050763724446451684, 32'sd-0.09653992310349856, 32'sd0.0072261025017472235, 32'sd-0.1435956641502242, 32'sd-0.0992277638258665, 32'sd0.02323928465152545, 32'sd0.03253348299977766, 32'sd-0.06833822136223636, 32'sd0.008502695926099032, 32'sd0.14017469080869938, 32'sd-0.05281792022153421, 32'sd-0.08999430731731044, 32'sd-0.03570258005029995, 32'sd0.02009082758905395, 32'sd0.0436532176481589, 32'sd0.018947017346872215, 32'sd-0.01556258075884042, 32'sd0.09717008562389821, 32'sd0.0028819124591642187, 32'sd0.033753095548801834, 32'sd0.00535129744873888, 32'sd0.09322199317485542, 32'sd0.0034870024892974666, 32'sd-0.06195215938638425, 32'sd-0.11578568134036334, 32'sd-0.06734935300532342, 32'sd-0.07628561872658778, 32'sd0.005821980390388461, 32'sd-0.03241449236251757, 32'sd-0.07049459671639405, 32'sd0.039749279753591264, 32'sd0.0293324097448388, 32'sd-0.017661752939915433, 32'sd0.005756338988737995, 32'sd-0.029530211025762917, 32'sd0.0039960639878569215, 32'sd0.005881929525802034, 32'sd-0.07513581175249434, 32'sd-0.031930376515665354, 32'sd-0.03179398768313039, 32'sd0.08623611670017453, 32'sd0.03969271685495661, 32'sd0.09455468514161305, 32'sd-0.01099471610531946, 32'sd0.07615717727984324, 32'sd0.06533916370157239, 32'sd0.12205659430092014, 32'sd-0.013134813157980933, 32'sd0.036611426353931685, 32'sd0.015491487914276306, 32'sd-0.08214600840374556, 32'sd0.030592980909186104, 32'sd0.045419021812981845, 32'sd-0.052584126115857624, 32'sd0.01825075272818996, 32'sd0.014251574715410446, 32'sd-0.024679975346401515, 32'sd-0.03256602380228932, 32'sd-0.006586111238606835, 32'sd0.058440817850948255, 32'sd-0.038914311397280785, 32'sd0.01825332485314257, 32'sd-4.76582196216264e-123, 32'sd0.0230827969063214, 32'sd0.030358261978173016, 32'sd-0.04531117542705176, 32'sd-0.08496106067407784, 32'sd-0.08072730541159316, 32'sd-0.04482018310430316, 32'sd0.03140904912268471, 32'sd-0.04595377127338848, 32'sd-0.06501811886598187, 32'sd-0.013728810710047765, 32'sd0.11631823477623, 32'sd0.17542133274734176, 32'sd-0.024530236971117204, 32'sd0.009827362954073875, 32'sd0.023195989479082326, 32'sd0.07250662645367205, 32'sd-0.011221004801484068, 32'sd0.006913756381290625, 32'sd0.07498617300851132, 32'sd0.023287960579327034, 32'sd-0.07251933929706361, 32'sd0.026623967708444864, 32'sd0.05983075283417478, 32'sd0.06574628322584676, 32'sd0.04068372194699809, 32'sd0.009571226790720472, 32'sd-1.3093369372239168e-122, 32'sd-8.918336159903426e-123, 32'sd7.393074106087025e-116, 32'sd-0.07370050399498214, 32'sd-0.04192978119212632, 32'sd-0.04343702942758616, 32'sd0.016037504984030226, 32'sd-0.05758551842685317, 32'sd-0.06987118654186456, 32'sd-0.10116947049983172, 32'sd-0.11349217575925005, 32'sd-0.038585363609139445, 32'sd0.015601469641148242, 32'sd-0.008734139869267632, 32'sd-0.06492041728883309, 32'sd-0.03140854943415859, 32'sd0.04666722576425792, 32'sd-0.012108257409098624, 32'sd-0.026357720345029326, 32'sd0.00951026711784202, 32'sd0.006484060852617925, 32'sd0.07857345955263445, 32'sd-0.018988328687831405, 32'sd-0.08979280561486308, 32'sd0.00016709968816322823, 32'sd-0.031156150144918376, 32'sd-0.00588263242681813, 32'sd0.03846212633113025, 32'sd4.9891876782687506e-120, 32'sd-1.7359081546256574e-126, 32'sd3.6680993433255983e-116, 32'sd0.034815711872205446, 32'sd0.04316925682239919, 32'sd0.07426513747460185, 32'sd0.03939393662379666, 32'sd0.09916170285030483, 32'sd0.0904589297841056, 32'sd-0.06480601624905329, 32'sd0.018200604564146503, 32'sd-0.08710913720214701, 32'sd0.09077503866960536, 32'sd-0.0356511801305913, 32'sd0.001040308330362659, 32'sd0.10419897831824514, 32'sd0.018651402798687662, 32'sd0.03021818567295506, 32'sd-0.02167016075448579, 32'sd0.017781718514160466, 32'sd-0.02922905282784756, 32'sd0.0038886978394022825, 32'sd0.07368798141155242, 32'sd0.034020071591916536, 32'sd-0.002343042388101391, 32'sd0.12582169892124687, 32'sd-0.10384761029468008, 32'sd-0.0064980616301435505, 32'sd-7.866348984857232e-126, 32'sd3.1819710071096695e-121, 32'sd-1.878495168232446e-121, 32'sd6.86650858834829e-124, 32'sd0.04611607655054745, 32'sd-0.07365171992480339, 32'sd0.004172292239791596, 32'sd-0.014907723328977742, 32'sd-0.01576075117509697, 32'sd0.0146332955683662, 32'sd-0.0520876332142408, 32'sd0.058194050952267554, 32'sd-0.08168995025530998, 32'sd-0.03448788106797109, 32'sd0.04632703762055219, 32'sd-0.02365928005933701, 32'sd0.04799820121412852, 32'sd0.07125896905820085, 32'sd0.060004844837120375, 32'sd0.08074656116805098, 32'sd0.11886614484555819, 32'sd0.08601514403482913, 32'sd-0.04233658020708198, 32'sd0.06553888160089158, 32'sd-0.06548468998132384, 32'sd-0.03383513907487718, 32'sd0.0003968769662768732, 32'sd4.628515668959625e-122, 32'sd4.82726892281529e-123, 32'sd3.300898488389333e-120, 32'sd-1.3752940531062419e-121, 32'sd2.413522404334943e-114, 32'sd-2.4540331534063484e-123, 32'sd0.05048879172150154, 32'sd-0.030040117297613033, 32'sd0.052957677759686426, 32'sd-0.036733115784170614, 32'sd-0.01825270477266632, 32'sd-0.09579791303908303, 32'sd0.037176596302632654, 32'sd-0.04514849916493554, 32'sd0.08733534524111278, 32'sd0.005263950447249235, 32'sd0.036420538413243206, 32'sd-0.07333665866184444, 32'sd0.06718666315267993, 32'sd0.030361983897286, 32'sd-0.048826567464673246, 32'sd-0.00020812435237275122, 32'sd0.006891092747546788, 32'sd0.024004181791005618, 32'sd-0.028357430086309792, 32'sd-0.020369123118948333, 32'sd-3.636333198226398e-116, 32'sd-2.1430677196562488e-119, 32'sd1.4507368485501342e-122, 32'sd-1.8672090092204964e-117},
        '{32'sd-5.777252681748961e-121, 32'sd-4.294922867055521e-115, 32'sd-1.1385801524370432e-119, 32'sd-1.68576211225833e-121, 32'sd4.821294527889001e-123, 32'sd1.0477500572344878e-120, 32'sd1.6997196137170257e-125, 32'sd9.090982217091904e-121, 32'sd-1.2957884375502378e-122, 32'sd1.5390850721146846e-123, 32'sd2.8510559085477326e-119, 32'sd8.593066964621704e-117, 32'sd-0.02945201299502953, 32'sd0.006129131642870007, 32'sd-0.02652725231347547, 32'sd0.04012479269150715, 32'sd-8.75034537226039e-120, 32'sd-8.005339161800211e-127, 32'sd4.66750767622327e-127, 32'sd3.105310440647812e-120, 32'sd7.785313590193593e-117, 32'sd-4.129310496686819e-125, 32'sd-3.5758799022366063e-119, 32'sd-2.6799321972681007e-114, 32'sd-1.0647195886805783e-124, 32'sd-1.776894074613201e-124, 32'sd3.339095800015602e-114, 32'sd-6.913967320214973e-127, 32'sd8.123804038165086e-119, 32'sd-1.9429272060476848e-124, 32'sd-8.766083096005644e-122, 32'sd2.260433881867402e-121, 32'sd-0.01030452194759564, 32'sd0.02905064094226699, 32'sd-0.05169215710237282, 32'sd-0.04401975984223706, 32'sd0.018858035977443764, 32'sd0.00873035297153687, 32'sd-0.006301292705625039, 32'sd0.01424650332516255, 32'sd0.07993662552723818, 32'sd-0.04896215581124591, 32'sd0.043609428459431186, 32'sd-0.009691264415976224, 32'sd-0.10412163454768195, 32'sd0.07287674148747782, 32'sd0.044021138257907086, 32'sd0.003885316483524509, 32'sd0.038451567634835905, 32'sd0.041243363889942576, 32'sd-0.03755023603115328, 32'sd0.013285353351029129, 32'sd5.913173636210401e-121, 32'sd-7.156033756683209e-116, 32'sd-2.294285973542343e-124, 32'sd-1.6138489260480738e-119, 32'sd2.597324379762619e-126, 32'sd1.1771099372107565e-127, 32'sd0.006441347420112001, 32'sd0.045163565539748485, 32'sd-0.04225684877108037, 32'sd0.08931326998703852, 32'sd0.08340409273266834, 32'sd0.04336314782502058, 32'sd0.08268211797512565, 32'sd-0.015887400273387278, 32'sd-0.00418607311033931, 32'sd0.022044432275909586, 32'sd0.012006400492340091, 32'sd-0.05262100519456, 32'sd-0.14169122181048086, 32'sd0.01809741363941014, 32'sd-0.08234930846471869, 32'sd-0.07309981545303493, 32'sd-0.016812878914294758, 32'sd0.021327018740613397, 32'sd-0.05964402730583028, 32'sd-0.05126210549523878, 32'sd0.005806797272340782, 32'sd0.07089966329074066, 32'sd0.023623683394309182, 32'sd-0.01349403029297998, 32'sd3.255805429343484e-116, 32'sd1.5048901042433409e-120, 32'sd1.758151560462309e-123, 32'sd-3.2438026931358545e-120, 32'sd-0.07368157889008876, 32'sd-0.03848942294319211, 32'sd0.021618533014136927, 32'sd0.0033367919863061543, 32'sd-0.008279461564697034, 32'sd0.052732438515257225, 32'sd0.0681590539517022, 32'sd0.0357456732059416, 32'sd0.12923096081882945, 32'sd0.026150305172407684, 32'sd0.03357693000931598, 32'sd-0.1156156591239752, 32'sd0.026107826914227344, 32'sd0.037990258702548, 32'sd0.05003873106618498, 32'sd-0.011782259032665067, 32'sd-0.007081238865113884, 32'sd0.031072716371634876, 32'sd-0.009885800158031078, 32'sd0.09000490834303197, 32'sd0.06587414107648833, 32'sd-0.0007491271740642403, 32'sd-0.07075920477950462, 32'sd0.07023605757722785, 32'sd0.0761161679436307, 32'sd6.28454980624547e-126, 32'sd-9.592999253320003e-122, 32'sd-0.0022700297177911605, 32'sd0.062274566943803976, 32'sd-0.006223053701502384, 32'sd0.0028751844711621274, 32'sd-0.023836049890480156, 32'sd-0.10499901940153616, 32'sd-0.05583315268583657, 32'sd-0.04024838858640725, 32'sd-0.20468079159314703, 32'sd-0.09470424249538811, 32'sd0.04039191912497773, 32'sd0.023417838579478486, 32'sd0.07761520027457217, 32'sd-0.01142848190133042, 32'sd-0.041071789819591815, 32'sd-0.0577989635198275, 32'sd-0.04783607672097135, 32'sd-0.1185322015549096, 32'sd-0.06942596369403686, 32'sd-0.1293212092429051, 32'sd-0.10051085938036033, 32'sd0.02102171391898535, 32'sd0.10866730009385908, 32'sd-0.012944907501274527, 32'sd-0.02859776994971553, 32'sd0.08087931174525423, 32'sd-0.01746060961192168, 32'sd-7.790164358645108e-121, 32'sd-0.023398601103011812, 32'sd0.04978354836076085, 32'sd-0.041029679815668345, 32'sd-0.02604949144489113, 32'sd-0.01338641258512533, 32'sd0.025264554419136758, 32'sd0.013535776009374568, 32'sd-0.012526693979130697, 32'sd-0.07536211668084306, 32'sd-0.007927924857461884, 32'sd-0.1625499769027353, 32'sd-0.0757812884556228, 32'sd0.04384573122949588, 32'sd0.10264251031791156, 32'sd0.02100739067595912, 32'sd0.060090446309657375, 32'sd-0.17275311873198174, 32'sd-0.23145605685091478, 32'sd-0.18382786616984373, 32'sd-0.043239669137901275, 32'sd0.027659198305571835, 32'sd-0.08521256608983255, 32'sd0.037017694626959516, 32'sd-0.05075407516201629, 32'sd-0.03095139497106388, 32'sd-0.023623995255436122, 32'sd-0.05273320570472005, 32'sd3.641410822665901e-123, 32'sd0.0121811164703602, 32'sd-0.039176518949409614, 32'sd-0.07200169542891888, 32'sd-0.014517555571406689, 32'sd0.05625528051615429, 32'sd-0.052335453199469494, 32'sd0.00916263011030485, 32'sd-0.10618319297014098, 32'sd0.18672087935131626, 32'sd0.1248197016475913, 32'sd-0.033388826082099775, 32'sd0.029602443526692432, 32'sd0.09137594605428252, 32'sd0.08314079646597851, 32'sd0.022165360983241754, 32'sd-0.02075190458224159, 32'sd0.0024487616769557218, 32'sd0.029877936226574708, 32'sd0.052632131972348735, 32'sd0.13057894745258783, 32'sd0.1519665769749868, 32'sd0.17499505160512804, 32'sd0.006193332581402138, 32'sd0.04411433881777352, 32'sd-0.03810975434302393, 32'sd0.015840387788548477, 32'sd0.012574184425207316, 32'sd0.03463571449204617, 32'sd0.023181878633708835, 32'sd-0.005746034597776652, 32'sd0.10212019827821511, 32'sd-0.020226261039073858, 32'sd0.007410449282859347, 32'sd-0.016889949825918543, 32'sd0.08467336724900215, 32'sd0.08312154657582044, 32'sd0.0299015060705884, 32'sd0.14903987173955205, 32'sd0.08997815388671707, 32'sd0.03309449658339582, 32'sd0.03208868577540847, 32'sd0.0479007318264299, 32'sd-0.10335819433374997, 32'sd0.0791273092238912, 32'sd0.09157596575497061, 32'sd0.07005318408716225, 32'sd0.09550371256651842, 32'sd0.0539712297266252, 32'sd0.0888163401764626, 32'sd0.0027164803250791084, 32'sd-0.11047108216905013, 32'sd-0.0015221654634319955, 32'sd-0.0053278983909407, 32'sd-0.051121126274199624, 32'sd0.030958509877816513, 32'sd-0.03817035970050128, 32'sd0.05677598568390001, 32'sd-0.0280059082611854, 32'sd0.11829157409644947, 32'sd0.01636622114475907, 32'sd0.06162008112335901, 32'sd-0.08133979190642822, 32'sd0.11826993415007064, 32'sd0.011243768980165075, 32'sd0.13581078398193952, 32'sd0.22496094354310034, 32'sd0.2128248878870203, 32'sd0.2161064762755343, 32'sd0.2509187034060767, 32'sd0.16890724791156186, 32'sd0.1801601955019494, 32'sd0.1750458424299648, 32'sd0.08166454671776958, 32'sd0.12314541744248521, 32'sd0.031301751054297444, 32'sd0.07692566973855146, 32'sd-0.02047717602263721, 32'sd0.13377301561892765, 32'sd0.10856480865291325, 32'sd0.023023146159938085, 32'sd0.019863078400312227, 32'sd-0.022421773063682968, 32'sd0.05945182884653336, 32'sd0.06241149078404949, 32'sd0.006005097106608354, 32'sd0.007118085768920562, 32'sd-0.1259895551366503, 32'sd-0.0010905234413735852, 32'sd-0.06760988666120074, 32'sd0.04212430038630045, 32'sd0.1394369250838178, 32'sd0.12267199841766901, 32'sd0.13314218993411295, 32'sd0.13513854128720024, 32'sd0.14145882769704424, 32'sd0.17851332227428035, 32'sd0.14774357856231593, 32'sd0.21727354622484452, 32'sd0.12608497034705657, 32'sd0.10451506004567596, 32'sd0.08393320522571933, 32'sd0.04516645593449604, 32'sd-0.13218044398434423, 32'sd-0.031435116347506495, 32'sd0.04387192136799846, 32'sd0.07304714721542975, 32'sd0.12498420851137182, 32'sd0.07057921366897928, 32'sd0.005418021839152477, 32'sd0.011404029578278435, 32'sd0.037827716886599375, 32'sd0.02131897933828741, 32'sd-0.005370163958064953, 32'sd-0.09715579403850344, 32'sd0.02258204519383645, 32'sd-0.04330701160825534, 32'sd-0.025248335398890983, 32'sd0.06047387675245942, 32'sd0.13621555417498551, 32'sd0.1636171525006271, 32'sd0.08611633365768723, 32'sd0.0766734731795985, 32'sd-0.049063106187111745, 32'sd-0.011700227537432523, 32'sd-0.0011338641325004078, 32'sd-0.07232577996615289, 32'sd-0.03739257996515354, 32'sd0.001046443825051059, 32'sd-0.12215430383239695, 32'sd-0.14172295080476374, 32'sd-0.03893749701066054, 32'sd-0.05299922540680246, 32'sd-0.06730635608994785, 32'sd0.1351286328396839, 32'sd0.08673637451013513, 32'sd0.08443669460326496, 32'sd0.025110125884208783, 32'sd0.028867111014166814, 32'sd-0.00796780796683761, 32'sd-0.024172200566275757, 32'sd-0.07989385846257412, 32'sd-0.03905461704447936, 32'sd0.01933442786303493, 32'sd0.0424874453439268, 32'sd-0.01648100922458847, 32'sd0.00884111715467953, 32'sd0.008404247526795696, 32'sd0.2183487767789113, 32'sd-0.01634229266669938, 32'sd-0.12540004441469924, 32'sd-0.12347631468232365, 32'sd-0.14689027970806737, 32'sd-0.24116652523312676, 32'sd-0.26980677653215773, 32'sd-0.1176535071686601, 32'sd-0.09580193917131599, 32'sd-0.18717491518599338, 32'sd-0.04109557574544097, 32'sd-0.15022577095643866, 32'sd-0.09154931734022674, 32'sd0.06664239575857404, 32'sd0.1352791794558271, 32'sd0.03113043101283766, 32'sd0.01537573339222277, 32'sd-0.08112778377924212, 32'sd0.06558856180581189, 32'sd-0.09097082013572827, 32'sd0.06228008734281687, 32'sd-0.07888929687540881, 32'sd0.02695622988713264, 32'sd0.02698330942438557, 32'sd0.01999736217981346, 32'sd0.007849646553422313, 32'sd-0.09515976034048541, 32'sd-0.10811320016097489, 32'sd-0.004516567856639435, 32'sd-0.2117792904567427, 32'sd-0.30866862072455464, 32'sd-0.23951891767676337, 32'sd-0.19039556720529993, 32'sd-0.21717925279644507, 32'sd-0.18176488828401377, 32'sd-0.010040949423049582, 32'sd-0.023962007127388274, 32'sd0.007088755858953536, 32'sd-0.022326019799808628, 32'sd0.011702624446501426, 32'sd-0.029332063682574176, 32'sd-0.053117187708292, 32'sd-0.12519242692535174, 32'sd-0.03881590435835101, 32'sd-0.06983942076023097, 32'sd0.09582717770649789, 32'sd0.044040084789381456, 32'sd0.0563224736382864, 32'sd-0.004354891294833585, 32'sd-0.05708314194995559, 32'sd-0.05683501688637517, 32'sd-0.037529967572949054, 32'sd-0.06759040331603873, 32'sd-0.10078721253015231, 32'sd-0.1840671727712796, 32'sd-0.26441020924952535, 32'sd-0.2572499368910115, 32'sd-0.33370197310426275, 32'sd-0.22313998196187707, 32'sd-0.06417396330360925, 32'sd-0.11754192162188665, 32'sd-0.148466010717273, 32'sd0.002584177495142148, 32'sd-0.11108869881859279, 32'sd-0.03223601902019506, 32'sd-0.06331053868055203, 32'sd0.06416468757954208, 32'sd-0.12163742935360429, 32'sd-0.22754905605989045, 32'sd-0.08452936268900088, 32'sd0.055194990229340546, 32'sd-0.012740773108873315, 32'sd0.13226199682128154, 32'sd0.039081379244705415, 32'sd-0.0018701233068749356, 32'sd0.06886494461757339, 32'sd0.009057726307033836, 32'sd-0.04885655359815759, 32'sd0.0177088291634432, 32'sd-0.010238714976197195, 32'sd-0.12479148955956598, 32'sd-0.22434255762429905, 32'sd-0.23497692751573984, 32'sd-0.25156063445437, 32'sd-0.1792680071903636, 32'sd-0.2667090880664519, 32'sd-0.025149806807621574, 32'sd-0.08012501057921244, 32'sd0.028118543030115833, 32'sd-0.005802349229502697, 32'sd0.030816075388768027, 32'sd0.044473629710206665, 32'sd0.016751390447507654, 32'sd0.17526474046919305, 32'sd0.11141266029859231, 32'sd-0.0036059859143656647, 32'sd-0.06890821165140765, 32'sd0.08058316394921043, 32'sd0.09924522496005186, 32'sd-0.008658977379513226, 32'sd-0.018400484026691723, 32'sd0.002995271907929389, 32'sd-0.011017043830787814, 32'sd0.02309694236825497, 32'sd-0.038680609657203366, 32'sd-0.01489665951828713, 32'sd-0.07688709892974861, 32'sd-0.15032662026679564, 32'sd-0.1711251675569821, 32'sd-0.2606584564496563, 32'sd-0.18591057305441042, 32'sd-0.16947019656175277, 32'sd-0.06878486273436686, 32'sd-0.07185786570044202, 32'sd0.04466740602223471, 32'sd0.08171153059643445, 32'sd0.040751468539902885, 32'sd0.13040787161468517, 32'sd-0.0029483206682498083, 32'sd0.16395055996648264, 32'sd0.07360387890480553, 32'sd0.11557814575590641, 32'sd-0.03742013495336801, 32'sd0.014958385486359459, 32'sd-0.03872956451079317, 32'sd-0.02510793581791386, 32'sd0.05386933226435056, 32'sd0.01223059607866593, 32'sd0.05441059925361039, 32'sd-0.11616510206907806, 32'sd0.012437635869492345, 32'sd-0.047722611846084444, 32'sd0.06463990999755408, 32'sd-0.04971138133051513, 32'sd-0.041577392894393245, 32'sd0.019881063724071925, 32'sd-0.09779389485796634, 32'sd-0.09976913198217374, 32'sd-0.01284997815459708, 32'sd0.023418103759063617, 32'sd0.07694006211766667, 32'sd0.05571604282623754, 32'sd-0.052047722424846836, 32'sd0.10047861067264596, 32'sd0.07750516574859277, 32'sd0.015728948637467415, 32'sd0.18439369362955124, 32'sd0.08160434574209374, 32'sd0.15305001444220734, 32'sd0.1041137561916003, 32'sd0.09432574481216197, 32'sd0.09718499192566696, 32'sd0.009586799449516091, 32'sd0.0605818189246161, 32'sd0.018327054706600024, 32'sd0.09721160205631524, 32'sd0.0033997253874234338, 32'sd-0.001086232107786059, 32'sd0.05348513202400181, 32'sd-0.07124757883476524, 32'sd6.626965688958365e-124, 32'sd0.03904941481071583, 32'sd-0.04014258199660717, 32'sd0.019186470465181765, 32'sd0.057108631639945444, 32'sd-0.06482677582741063, 32'sd-0.09645856397998931, 32'sd-0.006975466553820461, 32'sd0.032571767742159474, 32'sd0.0631076012323187, 32'sd0.02571791640135876, 32'sd0.014342483525716192, 32'sd-0.008086451853940987, 32'sd0.029778139139323315, 32'sd0.17466410930204318, 32'sd0.14944965285010298, 32'sd0.08965702488600989, 32'sd0.02235502742021841, 32'sd-0.01735236124783183, 32'sd0.08178427298620965, 32'sd0.020525426368840485, 32'sd-0.028213469865911646, 32'sd-0.12198866512888265, 32'sd-0.16436541884159475, 32'sd0.014279072661296202, 32'sd-0.06761408595759273, 32'sd-0.07401312831259749, 32'sd0.06202700681335876, 32'sd0.007240588413625962, 32'sd0.08063434832606857, 32'sd-0.03550110984681509, 32'sd-0.09223984353305953, 32'sd-0.03424057306267452, 32'sd-0.042953865575820316, 32'sd0.027373788645501388, 32'sd-0.0317078374976762, 32'sd-0.015148131827731007, 32'sd0.008195778616769187, 32'sd0.0664654962453377, 32'sd-0.0169419983580536, 32'sd0.056420559984252966, 32'sd0.08374011842357494, 32'sd0.10527103474339196, 32'sd0.16709801831330306, 32'sd0.049540088732038905, 32'sd0.010035427033674387, 32'sd-0.043389410122068865, 32'sd0.08650791626544586, 32'sd0.07736785097189038, 32'sd-0.1428559362961152, 32'sd-0.1775785999412992, 32'sd0.012395519699672536, 32'sd-0.09805243386640741, 32'sd-0.03333894793790772, 32'sd-0.1074396712425578, 32'sd0.06345035848967023, 32'sd-0.022897244853889987, 32'sd-0.01957741856188311, 32'sd0.024430353791388627, 32'sd0.02128221661217445, 32'sd0.05426076485722151, 32'sd0.006894500270169923, 32'sd0.030586882337771546, 32'sd0.04144644856884912, 32'sd0.02167346652712145, 32'sd-0.020682031100259297, 32'sd-0.07982631818548691, 32'sd0.020925886768930105, 32'sd-0.011219229888082766, 32'sd0.16964125273013406, 32'sd0.07960123054218166, 32'sd0.012246893608375572, 32'sd-0.01401295156676257, 32'sd-0.08623877619254831, 32'sd-0.16897287917972195, 32'sd-0.00998385805240783, 32'sd-0.03474587734504118, 32'sd-0.1361401930400099, 32'sd-0.03704220920621562, 32'sd-0.0213913012345726, 32'sd0.03012832229727964, 32'sd-0.07182126533011103, 32'sd-0.06438883385315512, 32'sd0.038318616931459853, 32'sd-1.3050716171538662e-123, 32'sd-0.06453198896905435, 32'sd0.07726731627262162, 32'sd0.10138543241118562, 32'sd0.04918185075451206, 32'sd0.06534630219674804, 32'sd0.07325366274358498, 32'sd0.08054316084947011, 32'sd0.0943387172845139, 32'sd0.03361153649454552, 32'sd0.006798551274071676, 32'sd-0.04578532643262065, 32'sd0.1057274589707174, 32'sd0.02951110517825085, 32'sd0.08600897343862868, 32'sd0.10185480572097963, 32'sd-0.016937038196306195, 32'sd-0.14158045797671018, 32'sd-0.08882397602767386, 32'sd-0.10316640949203554, 32'sd-0.07650165501622483, 32'sd-0.007283488227724265, 32'sd-0.008854329681873817, 32'sd-0.005956895811615611, 32'sd-0.036170477931501, 32'sd-0.014114250425419595, 32'sd-0.05412181576314467, 32'sd-0.03523984691042827, 32'sd0.033948056213040964, 32'sd0.007905059270497226, 32'sd0.05236669761386177, 32'sd-0.03769495324912605, 32'sd0.07862451107695481, 32'sd0.008773961902544014, 32'sd0.09234292753794439, 32'sd0.03940226226473104, 32'sd-0.04152382721309503, 32'sd-0.04749818586542015, 32'sd0.08438759217609791, 32'sd0.059607953492099415, 32'sd0.16819919021272273, 32'sd0.032143467691147926, 32'sd-0.017690907493672962, 32'sd-0.011070372549957465, 32'sd-0.058835537932630605, 32'sd-0.09607091117882048, 32'sd-0.03201516783098798, 32'sd0.0654046120128912, 32'sd-0.041278175894164375, 32'sd0.013782937305348679, 32'sd0.024870262177520676, 32'sd0.048607987996569055, 32'sd0.04917480900833347, 32'sd-0.0322884288250209, 32'sd-0.026454558986520292, 32'sd0.01573430618847344, 32'sd-0.0043061753768157945, 32'sd-0.03557412155384854, 32'sd0.003388519011081888, 32'sd-0.07203311856680197, 32'sd0.10560842870536688, 32'sd-0.007088013344249035, 32'sd-0.005866345901680479, 32'sd-0.08035638774353213, 32'sd0.058045099430748356, 32'sd0.006058079652972642, 32'sd0.15763256295793268, 32'sd0.14701376318709858, 32'sd0.03752418670826512, 32'sd-8.276784226768335e-05, 32'sd-0.05052077805665498, 32'sd0.010611472875254376, 32'sd-0.027227017800657397, 32'sd0.04356000487294996, 32'sd0.027840176404483264, 32'sd-0.05140580823569933, 32'sd-0.06120318130939533, 32'sd-0.040453198430643426, 32'sd0.08627578890129564, 32'sd-0.02014057320992546, 32'sd0.032872751688072424, 32'sd-0.09988325821666963, 32'sd-0.004871244152404758, 32'sd-0.0006364103320365207, 32'sd7.475048625451173e-117, 32'sd0.03226789491853631, 32'sd-0.09553022214851016, 32'sd-0.15786359638602815, 32'sd0.05324513571971087, 32'sd0.008258931367803892, 32'sd0.08571187372359028, 32'sd0.05883417895781278, 32'sd-0.01270515430322682, 32'sd0.01687049094350141, 32'sd0.002207976879973554, 32'sd0.04678110034947461, 32'sd0.016417339697731143, 32'sd-0.060760364648663634, 32'sd0.0900913187178823, 32'sd0.0738250681771286, 32'sd0.10441311638805921, 32'sd0.053955642945360836, 32'sd0.07333843654258894, 32'sd-0.06342701950758006, 32'sd-0.10101302122018434, 32'sd0.002482650491830974, 32'sd0.048659921029339505, 32'sd0.07836329541547316, 32'sd0.066522581271269, 32'sd-0.06382518288559319, 32'sd0.06439833915911888, 32'sd-6.0733210832814256e-124, 32'sd-2.639712251770394e-119, 32'sd-2.1324964825091545e-126, 32'sd0.09373380641059251, 32'sd-0.05102366628531745, 32'sd-0.04007419560765741, 32'sd0.02104032646864399, 32'sd0.05487378591070402, 32'sd-0.0026732621380732655, 32'sd-0.011376722336037929, 32'sd0.07547198994258826, 32'sd0.04797883485281983, 32'sd-0.04351294676733322, 32'sd-0.07695514631330014, 32'sd0.04109474449743666, 32'sd0.05653866417910092, 32'sd0.047401520913396555, 32'sd-0.013993387155523838, 32'sd-0.0036009594752343427, 32'sd-0.06690906993639649, 32'sd-0.18241540140608217, 32'sd0.029086608148831718, 32'sd-0.006224869406158044, 32'sd0.05451806361826151, 32'sd-0.043418822837357214, 32'sd0.045746294806777256, 32'sd-0.004515177834456466, 32'sd0.010000986477031144, 32'sd1.1260527854062808e-122, 32'sd-2.594649431289391e-125, 32'sd2.0892555396388452e-120, 32'sd0.04764689326977457, 32'sd0.10467436112289764, 32'sd0.08756448434110572, 32'sd0.04178216738409824, 32'sd0.06456076507765204, 32'sd0.08556093294259463, 32'sd0.03428458837380706, 32'sd0.11116986437443277, 32'sd0.13685739108010425, 32'sd-0.0451073900433792, 32'sd0.06763943577004845, 32'sd-0.023761328993707084, 32'sd-0.03192208008491599, 32'sd0.12977710026145228, 32'sd0.015242366091547077, 32'sd0.03219676424319891, 32'sd-0.14694786531273346, 32'sd0.04659750996734227, 32'sd-0.00470687483474536, 32'sd-0.007031626507552878, 32'sd0.016594747799711013, 32'sd0.04404598030586864, 32'sd0.02915561160457302, 32'sd0.07274207466754812, 32'sd-0.032957663407508504, 32'sd2.4382665278089692e-123, 32'sd9.451398604791183e-117, 32'sd7.858180625108788e-127, 32'sd-1.5834609524778823e-119, 32'sd-0.0050448462492758035, 32'sd-0.035732135973490384, 32'sd-0.10436056425444182, 32'sd0.01278210349182061, 32'sd0.09317413001002839, 32'sd-0.013113755437183836, 32'sd0.09152182845339434, 32'sd-0.10857304051006625, 32'sd-0.13880075114773432, 32'sd-0.08078063701429573, 32'sd0.07030355030763416, 32'sd0.007059183825780026, 32'sd0.05076044673650524, 32'sd-0.17201414453736458, 32'sd-0.0436789768757682, 32'sd-0.052056582501190087, 32'sd-0.044014161675874616, 32'sd-0.09498976758352654, 32'sd-0.09965424492388253, 32'sd-0.018415500560478488, 32'sd-0.042366879188865496, 32'sd-0.06364624757152394, 32'sd-0.034561757649887746, 32'sd1.899950040547777e-125, 32'sd-5.702383327901063e-121, 32'sd-1.6274459644763553e-117, 32'sd-6.81285018437699e-116, 32'sd-3.286573925571041e-120, 32'sd-6.022009329239473e-125, 32'sd0.00032369520454854947, 32'sd-0.0374229767263665, 32'sd0.05016122925240149, 32'sd-0.04765802672404152, 32'sd0.020306799780870154, 32'sd-0.027760326725819805, 32'sd0.08634829682330263, 32'sd0.04085488218629259, 32'sd-0.06595329711638734, 32'sd0.036463090747544946, 32'sd0.15067326957260596, 32'sd0.0898734317768421, 32'sd0.08720120813972082, 32'sd0.09370654838301871, 32'sd0.0652541561953173, 32'sd-0.09163281240688194, 32'sd-0.012661093774874429, 32'sd0.03030626837114725, 32'sd-0.052525143975345, 32'sd0.011417969607362884, 32'sd5.706478467236997e-115, 32'sd-1.1140939179134611e-122, 32'sd-2.388184571744847e-126, 32'sd4.182606555064941e-124},
        '{32'sd-2.1173058200926795e-117, 32'sd-1.5780861406841234e-125, 32'sd6.426346840356496e-120, 32'sd-1.7367509976363077e-125, 32'sd-1.8127671049198667e-128, 32'sd-2.365570885178276e-125, 32'sd3.6127714128882125e-116, 32'sd-1.4302629621846415e-118, 32'sd-4.375857034383688e-118, 32'sd5.674473482759995e-124, 32'sd-6.183160080752597e-122, 32'sd3.56551632964381e-119, 32'sd0.11838491477491644, 32'sd0.07851946699152237, 32'sd0.1425756791341308, 32'sd0.1414014073972393, 32'sd-8.031487669772406e-127, 32'sd2.053409930256114e-117, 32'sd-3.333982346220388e-119, 32'sd2.625365247324116e-123, 32'sd1.6069337435692875e-127, 32'sd2.538493270271351e-117, 32'sd-3.3920884403620476e-120, 32'sd7.215187609785813e-115, 32'sd4.081796951643977e-115, 32'sd6.840646975781812e-126, 32'sd-1.2583784080773863e-117, 32'sd3.3125088264930957e-116, 32'sd-1.2728406974212615e-117, 32'sd1.7673695634040167e-123, 32'sd-4.27712830057443e-123, 32'sd8.111375136086607e-127, 32'sd0.018331097454263447, 32'sd0.04454340187235606, 32'sd0.055413089395201745, 32'sd-0.046556164672744337, 32'sd-0.05384366930314438, 32'sd0.11091896946137013, 32'sd0.007103225080420004, 32'sd0.10949241990675317, 32'sd0.07711428570066096, 32'sd0.013541578018400334, 32'sd-0.05175611822037795, 32'sd0.05635630372133148, 32'sd0.08199272534879781, 32'sd0.06412901922462075, 32'sd-0.025711050044542366, 32'sd0.06131842864600418, 32'sd-0.0060338068538152755, 32'sd0.04412871195423533, 32'sd-0.020615261759461774, 32'sd0.048067106605271276, 32'sd2.1668617061431323e-127, 32'sd1.2128302991182785e-116, 32'sd-3.720336480444959e-119, 32'sd9.290932015737213e-123, 32'sd5.582069670550535e-119, 32'sd-6.854639542710473e-123, 32'sd0.1295924141590221, 32'sd-0.06069461440646114, 32'sd0.03941107720608704, 32'sd-0.02152287150385274, 32'sd0.11720414729221436, 32'sd0.053635137635770005, 32'sd0.05440305630954434, 32'sd0.015147526918835107, 32'sd0.16522631196282825, 32'sd0.022036834802279987, 32'sd0.05842037789681234, 32'sd-0.09089471505503129, 32'sd0.058268030653724885, 32'sd-0.02949343916706464, 32'sd0.09519905406617384, 32'sd0.16072141288845126, 32'sd-0.023238802373425273, 32'sd0.0901558960875871, 32'sd-0.03693891398985438, 32'sd0.09781480574386751, 32'sd-0.04111022436954896, 32'sd0.023303133915524615, 32'sd0.07079014970900589, 32'sd0.16791268936364687, 32'sd-5.706557161033672e-127, 32'sd1.921995712210805e-117, 32'sd-4.047882927141253e-125, 32'sd7.592314014645604e-119, 32'sd0.15501178162863366, 32'sd0.05475823112468289, 32'sd0.016281787851929203, 32'sd-0.04068684181124055, 32'sd0.003729388050867638, 32'sd-0.08538790840394135, 32'sd-0.020585393892389364, 32'sd-0.05058738517726795, 32'sd0.04574687749324813, 32'sd0.0945628075576822, 32'sd0.03501556066786646, 32'sd0.08206263258575971, 32'sd0.06407360530655926, 32'sd0.14341353019265218, 32'sd0.1410921094558669, 32'sd0.07788104702420927, 32'sd-0.09250795219005124, 32'sd-0.08287015527507545, 32'sd-0.09845386389234863, 32'sd0.06698293775323443, 32'sd0.13248985854212267, 32'sd-0.0043774448452708805, 32'sd-0.02101281178520966, 32'sd-0.03337361337772207, 32'sd-0.0832837722935253, 32'sd3.532497823143468e-116, 32'sd2.0810118614063412e-117, 32'sd0.05502568842231646, 32'sd0.03608049056879013, 32'sd-0.006264708871475887, 32'sd-0.10120907616724535, 32'sd-0.08384812454143721, 32'sd-0.04672383979419047, 32'sd-0.007166766699703753, 32'sd-0.02164649179399189, 32'sd-0.054227855671815026, 32'sd0.06801432362345922, 32'sd-0.020302305854560606, 32'sd0.025297015655518142, 32'sd0.11582622255600945, 32'sd0.04010140880991051, 32'sd-0.07208082232590347, 32'sd-0.09948423035878484, 32'sd-0.014912863738329528, 32'sd-0.038325952530709605, 32'sd-0.03765242155684217, 32'sd-0.12568583781987602, 32'sd-0.07374818200571796, 32'sd0.07873367432298717, 32'sd0.03846790065832179, 32'sd-0.10422365569362561, 32'sd-0.03070415075081913, 32'sd0.09542574419925758, 32'sd-0.04079530553654545, 32'sd-3.093064541479147e-122, 32'sd0.07443232700845258, 32'sd0.03427692741924148, 32'sd0.026828649852197618, 32'sd0.03848394639762665, 32'sd0.0005167682689449343, 32'sd0.0248480063483081, 32'sd-0.12465731495665507, 32'sd0.07491245675514255, 32'sd0.10924631963159308, 32'sd0.017060970212381833, 32'sd0.18527789886634527, 32'sd0.0844142286929311, 32'sd0.11175081035148414, 32'sd-0.07601789610346255, 32'sd-0.10401276562446063, 32'sd-0.15748612517039182, 32'sd-0.15180850121384892, 32'sd-0.09723436382776748, 32'sd-0.07853023214549637, 32'sd-0.04857338285386949, 32'sd0.00931103205798207, 32'sd-0.0194865345386476, 32'sd-0.011826750722032691, 32'sd0.041958679020993164, 32'sd0.14712435104602967, 32'sd0.11770257558123004, 32'sd0.06850245127271717, 32'sd-9.852971860029304e-120, 32'sd0.06801552221923422, 32'sd-0.006367484872636274, 32'sd-0.01575299978227523, 32'sd-0.05329622958677089, 32'sd-0.03919150715291369, 32'sd-0.15869286168968919, 32'sd-0.036566170485506394, 32'sd-0.02027147306216964, 32'sd-0.0400114372926209, 32'sd0.11530612139124106, 32'sd0.13810713939818914, 32'sd0.14842238262745996, 32'sd0.009744655045953253, 32'sd0.05295510030784483, 32'sd-0.06840945703994893, 32'sd-0.11698195675604123, 32'sd-0.007290044325105719, 32'sd-0.1457060872595807, 32'sd-0.05603985276402065, 32'sd0.005241385647412722, 32'sd0.11342475864786673, 32'sd0.07835853878845699, 32'sd-0.07923514483963683, 32'sd0.05107717695373922, 32'sd0.15229340209347014, 32'sd0.04817965230732198, 32'sd-0.0184776638737269, 32'sd0.1184715348543221, 32'sd0.05219214870387198, 32'sd0.02850337340524744, 32'sd-0.03584642924185124, 32'sd0.013637106465186021, 32'sd-0.03368033122878086, 32'sd-0.09089294239131154, 32'sd-0.12382228966766388, 32'sd-0.08454446955676019, 32'sd-0.0577897513064587, 32'sd0.013169541053445146, 32'sd0.08527359875771152, 32'sd0.12231333377387828, 32'sd0.05708273327184974, 32'sd-0.005192468101431761, 32'sd0.027897854711079636, 32'sd0.10439072677497159, 32'sd0.0734766899695814, 32'sd0.11421601117877571, 32'sd0.09976474550228114, 32'sd0.1210281037779462, 32'sd0.11491150421652226, 32'sd0.08304778375521137, 32'sd0.07783484465977629, 32'sd0.0016864192956083026, 32'sd0.030312511884126012, 32'sd0.09975306222802245, 32'sd-0.06817495442251664, 32'sd0.020085826167449267, 32'sd0.022579070729442246, 32'sd0.04917108170800635, 32'sd-0.006094146187179689, 32'sd0.10393718616867129, 32'sd-0.05862424572436207, 32'sd-0.0032258198001464135, 32'sd-0.06547649602827717, 32'sd-0.07384695762703194, 32'sd0.030584069100894614, 32'sd0.01988452159127983, 32'sd0.06361945891250742, 32'sd0.10582606433950752, 32'sd0.1634606062521756, 32'sd0.09559996217760262, 32'sd0.09654540549064117, 32'sd0.02990727485321227, 32'sd0.17303382866772213, 32'sd0.12590207225952577, 32'sd0.24626590293165235, 32'sd0.2573152940812804, 32'sd0.19542973048472156, 32'sd0.12863633294778337, 32'sd0.18238794531265087, 32'sd0.15286457047972768, 32'sd0.11117334741864288, 32'sd0.08720981646305845, 32'sd-0.03949610169828042, 32'sd0.10042124081725096, 32'sd0.02255331772121353, 32'sd0.09584241096803943, 32'sd0.11681246967391691, 32'sd0.12416328337782115, 32'sd0.0335365034913696, 32'sd-0.04745900302252787, 32'sd-0.12253746606939461, 32'sd-0.12574968804468178, 32'sd-0.04294778201603878, 32'sd-0.07602424809376039, 32'sd0.06748853523009755, 32'sd0.06305517840215176, 32'sd0.17523725562861048, 32'sd0.10341180008720303, 32'sd-0.04652305213382201, 32'sd0.19108793930563417, 32'sd-0.0358642484652476, 32'sd0.11019427965511018, 32'sd0.11842713657157411, 32'sd0.09910320713453716, 32'sd0.05759865206708964, 32'sd0.10072646360706569, 32'sd0.013852908800599806, 32'sd0.10790191037739143, 32'sd-0.05718058756977316, 32'sd0.03603900553667202, 32'sd0.08167560258389951, 32'sd0.06069104871796071, 32'sd-0.028916549303382152, 32'sd0.10431480760742913, 32'sd0.03950980599795387, 32'sd0.03198978996701783, 32'sd0.01287059397135467, 32'sd-0.009653686277713293, 32'sd-0.051412698675175554, 32'sd-0.05286531437427678, 32'sd-0.059181536718205224, 32'sd0.1256266329624475, 32'sd0.010658020074228421, 32'sd0.11253363644923156, 32'sd0.09416440676960212, 32'sd-0.057678380015334006, 32'sd0.07484238371089799, 32'sd0.09881825894764541, 32'sd-0.07482952028512425, 32'sd0.015182317629099589, 32'sd-0.06931178622865777, 32'sd0.04781548169052161, 32'sd0.0638275322450022, 32'sd-0.03220387289906915, 32'sd-0.025890267092167796, 32'sd-0.05422691249276527, 32'sd-0.08224434905388464, 32'sd-0.0076634436570415685, 32'sd0.0719621716337039, 32'sd0.07824968259198901, 32'sd0.03164745724463229, 32'sd-0.025275813716834097, 32'sd0.0603667855528797, 32'sd-0.005595573877139011, 32'sd-0.11629653774625567, 32'sd0.0313662265307814, 32'sd-0.055650526195346946, 32'sd-0.05792979851836748, 32'sd0.03574211752811353, 32'sd0.02781496923675316, 32'sd0.03120698703976183, 32'sd0.125599104599326, 32'sd-0.001896675057333867, 32'sd-0.0032028781410729035, 32'sd0.006078092192280709, 32'sd-0.08268918398472269, 32'sd-0.12017968354792906, 32'sd-0.13802086100041738, 32'sd-0.17339303642530962, 32'sd-0.15794282684496186, 32'sd0.043359986069811694, 32'sd-0.0973109663595645, 32'sd-0.03655931566590101, 32'sd-0.09897153899009557, 32'sd-0.07209391731476203, 32'sd0.008949978037270734, 32'sd0.07352241047173243, 32'sd0.0880195812389781, 32'sd0.06267054594617752, 32'sd-0.039960610060885936, 32'sd0.011148897082379962, 32'sd-0.028006278753497364, 32'sd-0.04876944904024207, 32'sd-0.1002037060317406, 32'sd-0.07362958795396109, 32'sd-0.05886830833290523, 32'sd0.007002793941741202, 32'sd-0.08616898450801164, 32'sd-0.0015180042487014484, 32'sd0.07306475973783587, 32'sd-0.060154138406084884, 32'sd-0.09867270319572016, 32'sd-0.04571832805602994, 32'sd-0.10175942123499271, 32'sd-0.048352745790120694, 32'sd-0.1361689833655951, 32'sd-0.16598171572931927, 32'sd-0.05141686363445472, 32'sd0.015599755931292566, 32'sd0.07262747061652847, 32'sd-0.04216617518499283, 32'sd-0.007660798000010573, 32'sd-0.08472955977060231, 32'sd-0.13150342562698425, 32'sd0.06319617592217341, 32'sd0.06026044135935052, 32'sd0.05543804181846357, 32'sd0.04279694006582831, 32'sd0.06699035473626248, 32'sd-0.14088798566051, 32'sd0.08204137290271986, 32'sd-0.010941035976969885, 32'sd0.0059351358060164665, 32'sd-0.14491218448231766, 32'sd-0.050954996720812974, 32'sd-0.06024431576201542, 32'sd-0.13148946645573314, 32'sd0.04596219017137139, 32'sd0.04485149749136859, 32'sd0.02061141760639572, 32'sd-0.02468150708107644, 32'sd0.012869620162771562, 32'sd-0.004815913542298116, 32'sd-0.02595591319466989, 32'sd-0.11926722104492804, 32'sd-0.13179728970205798, 32'sd-0.13887945712754415, 32'sd-0.05946864526831502, 32'sd-0.11074490021555242, 32'sd-0.18095366868794557, 32'sd-0.06809811032030741, 32'sd0.039432556194799816, 32'sd0.03923671395473358, 32'sd0.1382857174961445, 32'sd0.06055906772295195, 32'sd-0.0804703445245811, 32'sd-0.05637151989888669, 32'sd-0.09222915994847099, 32'sd0.05417954423340419, 32'sd-0.18023956974886945, 32'sd-0.029488928142648904, 32'sd-0.16214152523987113, 32'sd-0.15236474370015388, 32'sd-0.10264344453037279, 32'sd-0.09609431103931737, 32'sd0.10308155900488837, 32'sd0.18498630878794406, 32'sd0.09417803045186819, 32'sd0.03628374086212572, 32'sd0.10189031945633761, 32'sd0.04336195884808798, 32'sd-0.08661973286181603, 32'sd0.017298927285683042, 32'sd-0.17452434415111834, 32'sd-0.08864148273753589, 32'sd-0.1156363047791847, 32'sd-0.059477276793750956, 32'sd-0.12282398897134178, 32'sd0.032137297795078686, 32'sd0.016020461085669496, 32'sd0.08640306790166855, 32'sd-0.0014090728765365583, 32'sd0.005894174282210164, 32'sd-0.039644936462007854, 32'sd-0.08854487902247417, 32'sd0.0059974513652004515, 32'sd-0.08458593299540479, 32'sd-0.20320026358271973, 32'sd-0.13143614299193646, 32'sd-0.10454815363027564, 32'sd-0.17414728264629875, 32'sd-0.06122182419240001, 32'sd0.04053538866905847, 32'sd0.11212597523125264, 32'sd0.17880258809341487, 32'sd0.08945926493191687, 32'sd-0.08330332154078027, 32'sd-0.03600877915607983, 32'sd-0.009988438302169361, 32'sd-0.015871349820034634, 32'sd-0.13908740903676436, 32'sd-0.07738273403463675, 32'sd-0.02918371809873486, 32'sd-0.10470739997453352, 32'sd-0.14871626012016212, 32'sd-0.08742557981298398, 32'sd0.08683603295071592, 32'sd0.09718564074190308, 32'sd0.0753765013115248, 32'sd0.03674486715274053, 32'sd0.0229548941188597, 32'sd0.007583832803045861, 32'sd-0.10881703338959724, 32'sd0.07440034599952842, 32'sd-0.0707602156190703, 32'sd-0.0690935507208325, 32'sd-0.1187522320709116, 32'sd-0.15683849805445546, 32'sd-0.16196814879266194, 32'sd0.052938955773470686, 32'sd0.19014655936241134, 32'sd0.15752206737808058, 32'sd0.18593219475090922, 32'sd0.03921931317963868, 32'sd-0.11278472877798967, 32'sd-0.11524559626051245, 32'sd-0.026100513924252205, 32'sd-0.15019614013832924, 32'sd-0.14301576732236385, 32'sd-0.12083589183561155, 32'sd0.0036702864344160054, 32'sd0.13196505758419, 32'sd0.028135408181965874, 32'sd0.061234840998672116, 32'sd0.12009868774349375, 32'sd0.07389839337361198, 32'sd0.09296344231126151, 32'sd8.864793639655381e-122, 32'sd0.022785211874638587, 32'sd-0.011963500551444963, 32'sd-0.06678014915285395, 32'sd-0.018652405163286145, 32'sd0.010445658716742872, 32'sd0.022834544627473755, 32'sd0.06546983354808002, 32'sd-0.07434768754032345, 32'sd-0.054970344918845226, 32'sd0.13521571990761524, 32'sd0.3219273181368047, 32'sd0.33835086456056845, 32'sd0.12136252783815357, 32'sd-0.0971872761710908, 32'sd-0.1567415874550466, 32'sd-0.12977875205775127, 32'sd-0.03209725720370662, 32'sd-0.059447766969209906, 32'sd-0.08917650999024468, 32'sd0.0341814800185984, 32'sd0.0648951785609256, 32'sd0.18765162428213802, 32'sd0.0942700849687731, 32'sd0.004711220985202482, 32'sd0.14750969230553695, 32'sd0.07225614118423142, 32'sd0.024927511720016553, 32'sd0.005901993044214922, 32'sd-0.013900242847808546, 32'sd-0.014595874559099786, 32'sd0.023699299726133216, 32'sd-0.039726040988924766, 32'sd-0.12784300817911173, 32'sd0.023198594597360678, 32'sd0.08169080623530303, 32'sd0.04385823300539996, 32'sd0.11401641816713, 32'sd0.15211224989798888, 32'sd0.22860886941299574, 32'sd0.2539335113405784, 32'sd-0.02996147674304768, 32'sd-0.262005386384858, 32'sd-0.3379021939324299, 32'sd-0.12687997345018406, 32'sd0.03793923716907628, 32'sd-0.0984247740747627, 32'sd-0.013443619085089955, 32'sd0.052321439018550665, 32'sd-0.024364868170448147, 32'sd0.07824237606373344, 32'sd0.01194904583561666, 32'sd0.11442635625872119, 32'sd0.1206268318346796, 32'sd0.19434554045118335, 32'sd0.05758554959754736, 32'sd0.008475547590157272, 32'sd0.043970370132598594, 32'sd-0.04492901373878275, 32'sd0.013053367371517268, 32'sd-0.09907749006180969, 32'sd-0.09339625624207905, 32'sd-0.034265200754586306, 32'sd-0.000253503401036233, 32'sd0.06308177069544413, 32'sd0.037401998370581904, 32'sd0.2058682248417044, 32'sd0.26856379391317353, 32'sd0.1736827428633523, 32'sd-0.11933035726742472, 32'sd-0.22405543586027418, 32'sd-0.23057031496404376, 32'sd-0.06769130608440925, 32'sd-0.06305027342349012, 32'sd-0.07561536927368534, 32'sd-0.002024580638572797, 32'sd0.08713777978571682, 32'sd-0.011263287139404641, 32'sd-0.09082082837706397, 32'sd-0.0013836183539702998, 32'sd0.05796933908804433, 32'sd0.14606090880576464, 32'sd0.1506278859984733, 32'sd-0.007191327974343512, 32'sd-1.616704504016549e-126, 32'sd-0.0038246103845715213, 32'sd0.01260133936062703, 32'sd-0.01586723293903681, 32'sd-0.12597129318346012, 32'sd0.05995086292411027, 32'sd0.002582480124604568, 32'sd0.0071499142706846755, 32'sd0.09229237789123167, 32'sd0.03764217145971333, 32'sd0.1960144255834863, 32'sd0.2599286714031828, 32'sd0.0020111223425033254, 32'sd-0.19870433301877777, 32'sd-0.2881677531152238, 32'sd-0.14746644094946032, 32'sd-0.023199618792982702, 32'sd-0.047177726741487465, 32'sd0.014157961057770042, 32'sd-0.010419774564231758, 32'sd0.011111960702198472, 32'sd-0.08642658874275513, 32'sd-0.011077106458640037, 32'sd-0.02263718371668288, 32'sd0.009318853484019906, 32'sd0.05819516753320684, 32'sd0.04299668495759055, 32'sd0.14756697504707594, 32'sd0.04045906034213314, 32'sd0.06177831000564999, 32'sd0.09232089698172546, 32'sd0.08520783488346012, 32'sd0.09580341265101192, 32'sd0.03553829306114906, 32'sd-0.020864863255311207, 32'sd0.07906743378566182, 32'sd0.03526055820936917, 32'sd0.22034695117104838, 32'sd0.12884378618655715, 32'sd0.051720742660590506, 32'sd0.07871826926380343, 32'sd-0.08784178001064058, 32'sd-0.14013762793351522, 32'sd-0.18863134937298448, 32'sd-0.07822835859667467, 32'sd-0.004563776877127489, 32'sd-0.13393638627410454, 32'sd-0.06223160076046355, 32'sd0.06415553326702819, 32'sd0.05796744755870994, 32'sd0.0036648986015648966, 32'sd0.0058819252615522274, 32'sd0.028567823609871156, 32'sd0.11240958422264319, 32'sd-0.03569321430336791, 32'sd0.08526478089674837, 32'sd-0.03742852224721462, 32'sd-0.04937686639717146, 32'sd0.009068844812503366, 32'sd-0.05668341887205333, 32'sd-0.0590869854240778, 32'sd0.08603677542574063, 32'sd-0.010204981396766805, 32'sd0.001972648562688707, 32'sd0.14720684637631376, 32'sd0.17201680621118706, 32'sd0.0301798152690365, 32'sd-0.0579060614017741, 32'sd-0.1294143018322949, 32'sd-0.0270352284260977, 32'sd-0.12094778502285863, 32'sd-0.0665286598362569, 32'sd-0.1862623402477532, 32'sd-0.07789598190072884, 32'sd0.011051706118783582, 32'sd-0.06814897925519978, 32'sd0.07550309693818993, 32'sd0.018764618197079367, 32'sd0.019122840945243167, 32'sd-0.03538803815133033, 32'sd-0.012300326934876408, 32'sd0.0983682567993839, 32'sd-0.010256218803985724, 32'sd0.06613368841137902, 32'sd1.5956873214521122e-123, 32'sd-0.04988180206226369, 32'sd0.025572572486313113, 32'sd-0.015357559862256209, 32'sd-0.04625611096664706, 32'sd0.06946360576086759, 32'sd0.14700316354742338, 32'sd-0.05145326935215154, 32'sd0.010658322002048241, 32'sd0.08526864642441921, 32'sd0.12548457583528752, 32'sd0.04354135622244846, 32'sd0.014986302374580672, 32'sd-0.08589915253893408, 32'sd0.011131437218814752, 32'sd0.037624798898016516, 32'sd0.011301601944352228, 32'sd-0.022392827731887825, 32'sd-0.11416513417006137, 32'sd0.1275547356563554, 32'sd-0.03605512516221941, 32'sd-0.11721889310476151, 32'sd-0.09264409728711183, 32'sd-0.14747828088871898, 32'sd0.06930317152868982, 32'sd0.043359899873467535, 32'sd0.006544100086734173, 32'sd1.0270759794263956e-124, 32'sd4.697162671452009e-123, 32'sd1.7576587198901527e-122, 32'sd0.003177536793317326, 32'sd-0.09879518176869993, 32'sd-0.13948912253202594, 32'sd-0.11547864749762793, 32'sd-0.012586911098096447, 32'sd-0.01292665132468446, 32'sd0.04169135004711109, 32'sd-0.03228108092598809, 32'sd0.019058213908418997, 32'sd0.07417626932554741, 32'sd0.20188941169271216, 32'sd0.12146860125888714, 32'sd0.04947067350391924, 32'sd-0.07459667230017199, 32'sd0.028806683515630673, 32'sd-0.08721049108570655, 32'sd0.03529910041690135, 32'sd0.055390730645594057, 32'sd-0.11648520919028839, 32'sd-0.009954093796348672, 32'sd0.009877470268876356, 32'sd-0.008161536885656859, 32'sd0.05488113035262143, 32'sd0.022920317861028643, 32'sd0.03386527827457903, 32'sd-2.1849898926429955e-126, 32'sd9.12901841596749e-121, 32'sd-3.929373493053841e-119, 32'sd-0.0056954275346893365, 32'sd0.05175789238812598, 32'sd0.10755620489111418, 32'sd-0.06391956660868527, 32'sd-0.10271568860382894, 32'sd0.04479177246657562, 32'sd0.031001802222983762, 32'sd0.05150626189289034, 32'sd-0.08843282948240158, 32'sd0.018867559212376386, 32'sd0.008453942747128785, 32'sd0.05529048459481812, 32'sd-0.0711951441587253, 32'sd-0.06714185845266746, 32'sd-0.08824481834017665, 32'sd0.06031344052250871, 32'sd-0.04615884788996943, 32'sd-0.18854341924190765, 32'sd-0.13340517619993736, 32'sd-0.1108167538517803, 32'sd-0.07027322926788365, 32'sd0.03884106188695352, 32'sd-0.03701842521254726, 32'sd0.00922574049672671, 32'sd0.02174527925104437, 32'sd-3.0185654006379613e-118, 32'sd1.6568544250202222e-127, 32'sd1.0841473626971732e-115, 32'sd1.7387724385513882e-125, 32'sd0.13098482470710165, 32'sd-0.004643472895489277, 32'sd0.09723318044938, 32'sd0.01632749283455561, 32'sd0.024153724611262143, 32'sd0.05386428099536598, 32'sd-0.029443933633611554, 32'sd0.06319466027993996, 32'sd0.04408248343975603, 32'sd-0.1054601215809334, 32'sd-0.038332970061236336, 32'sd-0.09894837088579582, 32'sd-0.08420046405437043, 32'sd0.026502863990658376, 32'sd0.07558648378778147, 32'sd-0.054603811865253704, 32'sd0.0858908174288098, 32'sd0.03366659614134603, 32'sd0.00805959129409697, 32'sd0.07642899412714553, 32'sd-0.05490894898327263, 32'sd0.07400100768819998, 32'sd0.09379810416696942, 32'sd6.547379773215907e-115, 32'sd4.9145912416963395e-124, 32'sd-2.642435966482919e-123, 32'sd-2.714060548035409e-118, 32'sd-3.044154519068758e-126, 32'sd-6.44613512924026e-115, 32'sd0.12710326532216762, 32'sd0.07652877823475453, 32'sd0.08219063375906335, 32'sd0.06496701516768245, 32'sd0.005140687928563876, 32'sd-0.08454867986654184, 32'sd0.03297199555024873, 32'sd0.057000692677166155, 32'sd-0.04455100518636819, 32'sd0.10848211405507037, 32'sd0.13295306246942773, 32'sd0.08625066846755511, 32'sd0.09301621369995229, 32'sd0.04330200601381949, 32'sd0.016703106604565223, 32'sd0.1376296663437826, 32'sd0.09107230651050671, 32'sd0.05504267660118679, 32'sd-0.06328745643092212, 32'sd0.06292015698379415, 32'sd9.417160299120035e-117, 32'sd3.0381228936086844e-123, 32'sd-1.5776958611011189e-121, 32'sd-9.333578743719252e-117},
        '{32'sd1.51685690272491e-126, 32'sd9.299777356930232e-125, 32'sd-5.192933114637386e-118, 32'sd7.956229560937905e-122, 32'sd1.4065502679762945e-123, 32'sd1.5604035946145572e-121, 32'sd4.33269072505107e-124, 32'sd8.642931306022299e-117, 32'sd1.3614451075779646e-125, 32'sd-5.244348746930323e-119, 32'sd-1.2622121835251898e-116, 32'sd2.563127430759761e-120, 32'sd0.005525489573701383, 32'sd0.014907005360560843, 32'sd0.016230932872843756, 32'sd0.1024806042857457, 32'sd6.852833785526406e-115, 32'sd-1.0647206365038067e-117, 32'sd4.08046926855558e-123, 32'sd5.358078255234176e-124, 32'sd-3.0690545248130993e-121, 32'sd1.6225023614865048e-121, 32'sd5.344338271006819e-120, 32'sd-6.674076978791344e-126, 32'sd-4.8200689774615165e-120, 32'sd1.8257665245690956e-117, 32'sd5.5635082764419836e-120, 32'sd6.695926339804085e-126, 32'sd-2.8159959302205247e-122, 32'sd-3.6089739712249586e-122, 32'sd1.1369350119918606e-126, 32'sd1.727442812853062e-123, 32'sd0.030548174965372363, 32'sd-0.040296103261533704, 32'sd0.028918353404049628, 32'sd0.05322730988831027, 32'sd-0.014114558771548576, 32'sd-0.01730010006235759, 32'sd0.13978508282096688, 32'sd0.133532209427974, 32'sd0.062145650332192146, 32'sd0.02465706652853584, 32'sd-0.06487442018442482, 32'sd0.01173191936649052, 32'sd-0.03736873795463041, 32'sd-0.01213586232285079, 32'sd-0.03632474854127667, 32'sd-0.010958040525519236, 32'sd0.1046129552367646, 32'sd0.039699746102010186, 32'sd0.08707572294507532, 32'sd0.04445606485440228, 32'sd3.2766647773170693e-121, 32'sd-2.0342586172003545e-120, 32'sd1.705657316770133e-125, 32'sd-2.5772668368036076e-126, 32'sd-5.1024091051386753e-126, 32'sd-1.4251339954709451e-128, 32'sd0.08814583772363023, 32'sd0.07178336264475693, 32'sd0.026633043605485487, 32'sd0.004904084829667863, 32'sd0.11300502524540733, 32'sd0.09313314261227335, 32'sd0.10175331444852247, 32'sd0.08318756117334712, 32'sd0.004845866950990963, 32'sd0.053592543938223366, 32'sd-0.0360974040447247, 32'sd-0.10509977057598338, 32'sd-0.039610549686371864, 32'sd-0.049175820102903965, 32'sd0.0033306122863986896, 32'sd0.0687951763197355, 32'sd0.09763688350778273, 32'sd0.1069964923110662, 32'sd0.04505919234832111, 32'sd0.126642986712308, 32'sd0.09518371192463837, 32'sd-0.012031569708924161, 32'sd0.04018151580067562, 32'sd0.03303517220821313, 32'sd1.4205599020160156e-118, 32'sd7.345361516864911e-125, 32'sd-1.0860487146575508e-124, 32'sd2.1177991126048107e-127, 32'sd0.010147342237654537, 32'sd0.043930649974372016, 32'sd0.07241071581677445, 32'sd0.044548148713416884, 32'sd0.0711908218622183, 32'sd-0.06859055165035535, 32'sd-0.010187885524184658, 32'sd0.030651729600272164, 32'sd-0.11784234059411078, 32'sd-0.09780159915313873, 32'sd-0.014806547215498105, 32'sd-0.1487668589482998, 32'sd-0.030262100864690614, 32'sd-0.11349961170697244, 32'sd-0.015324620110225734, 32'sd-0.008264217699727969, 32'sd0.11287671122978908, 32'sd0.08741398277857024, 32'sd0.07760133395823958, 32'sd0.08511617271461275, 32'sd-0.005699774053763447, 32'sd-0.06094094058952591, 32'sd0.0030626219198562287, 32'sd-0.15311360800848733, 32'sd0.07549269037723019, 32'sd-6.988316929224385e-117, 32'sd-6.704054613722329e-115, 32'sd-0.002984191087497015, 32'sd0.009591306414806435, 32'sd0.024612551949222166, 32'sd0.005137236524606395, 32'sd-0.03816278170966586, 32'sd-0.07286241091421747, 32'sd-0.0999960565814527, 32'sd0.01710319507403807, 32'sd-0.1323411866278002, 32'sd-0.1243018512864199, 32'sd0.11682319159464939, 32'sd-0.053204116304745135, 32'sd0.05526271234488113, 32'sd-0.05742453205834766, 32'sd0.048218080337410575, 32'sd-0.00277270686738516, 32'sd-0.09163369994125536, 32'sd-0.0730799707213078, 32'sd-0.127159272198394, 32'sd-0.10584548629551424, 32'sd0.029453833765403586, 32'sd-0.026400945983362525, 32'sd-0.0006106286887605221, 32'sd-0.04018572494907329, 32'sd0.018543108140831998, 32'sd0.07535145432840092, 32'sd-0.04465837452937871, 32'sd3.505464047195044e-117, 32'sd0.05155590849768711, 32'sd-0.07150614951772245, 32'sd-0.10275618799214896, 32'sd0.004638573242451751, 32'sd0.017941819414815093, 32'sd-0.12395489204741282, 32'sd0.025083664014425362, 32'sd-0.1340317735294578, 32'sd-0.15833024515940042, 32'sd-0.15603998695089777, 32'sd-0.11506154195987421, 32'sd-0.15843968988476342, 32'sd-0.10993006961356297, 32'sd-0.17804893956435772, 32'sd-0.11790653302991917, 32'sd-0.10598046197633297, 32'sd-0.12142840221136879, 32'sd-0.029488598012308805, 32'sd-0.09191721344638885, 32'sd0.09186558605264598, 32'sd-0.040342735646964153, 32'sd0.032553410353239824, 32'sd0.052519541051548824, 32'sd0.05570029961058879, 32'sd-0.024201593825398427, 32'sd-0.05709620780506723, 32'sd-0.038574909317065066, 32'sd3.897275008461251e-119, 32'sd0.04091932071353586, 32'sd0.055368931137400865, 32'sd0.059911155691072714, 32'sd0.06346910234925394, 32'sd0.02513243690862799, 32'sd0.12400049620066267, 32'sd0.046114120972585715, 32'sd-0.003489135369306035, 32'sd-0.12003024523955809, 32'sd-0.22428263027850556, 32'sd-0.2013986001888323, 32'sd-0.23314791839911234, 32'sd-0.11260944476816723, 32'sd-0.05184003551577618, 32'sd-0.1862272866062075, 32'sd-0.11673866701904112, 32'sd0.040357947214173955, 32'sd0.003548942346964422, 32'sd0.07374637631835519, 32'sd0.006661209383682139, 32'sd0.05536214103806614, 32'sd0.06510654599667837, 32'sd-0.062014635646056984, 32'sd-0.03209654800613921, 32'sd0.09246304453521445, 32'sd0.08868672221045845, 32'sd-0.005314840831916021, 32'sd0.03529176678457177, 32'sd0.017558154360254156, 32'sd-0.12660855684099773, 32'sd0.027851422681601193, 32'sd0.06344487951963963, 32'sd-0.027063129466522774, 32'sd-0.06561109821715704, 32'sd0.060624327054981386, 32'sd0.0901973940679305, 32'sd-0.13934980563264637, 32'sd-0.1787070465656759, 32'sd-0.10853459597940068, 32'sd-0.1242411464708272, 32'sd-0.11430505948472, 32'sd-0.04406752726214257, 32'sd0.13378248218961658, 32'sd0.07820994661962016, 32'sd-0.017220781160801706, 32'sd0.06944838233987435, 32'sd0.08063279255398788, 32'sd0.056376389497411764, 32'sd0.11810040650225491, 32'sd0.14471688253779333, 32'sd0.09088057947923123, 32'sd0.01724722913430014, 32'sd0.0099189624989787, 32'sd0.10719368015455907, 32'sd0.039588391988895126, 32'sd0.048065114760780306, 32'sd-0.07742425121303166, 32'sd-0.07816476213337316, 32'sd-0.1303630873063355, 32'sd-0.048652754701196115, 32'sd-0.06606724030733993, 32'sd-0.13744619475499073, 32'sd-0.15478643543941878, 32'sd-0.08503576829730165, 32'sd-0.1298531797686598, 32'sd-0.10240966762518715, 32'sd-0.10237001360556115, 32'sd-0.1354966657600505, 32'sd0.014777599515886653, 32'sd-0.01788318518610813, 32'sd-0.01695591642734948, 32'sd0.07365445320297014, 32'sd0.0828451424035828, 32'sd0.0019749088795485317, 32'sd0.03581721144308893, 32'sd0.16324662297263057, 32'sd0.10113118421082953, 32'sd0.008650173063178796, 32'sd0.05134793435501701, 32'sd0.09308093030340804, 32'sd0.015561131054686353, 32'sd0.05199913313349687, 32'sd0.044051990628082835, 32'sd-0.013765431722525047, 32'sd0.014433494095561756, 32'sd0.015873978364121362, 32'sd0.0776254685617909, 32'sd-0.13165702314413885, 32'sd-0.11568580269493241, 32'sd-0.2441467393842104, 32'sd-0.13078729415041843, 32'sd-0.05966090071998916, 32'sd-0.004231765871110082, 32'sd-0.10660005081477708, 32'sd-0.1160170856849655, 32'sd0.08641485243876504, 32'sd0.1961826214986819, 32'sd0.0018814435471452852, 32'sd6.92432137347602e-05, 32'sd-0.02173135792430417, 32'sd0.07948922923574248, 32'sd-0.09203281409139909, 32'sd0.004146783953037365, 32'sd0.04294390759690763, 32'sd0.04395839236586247, 32'sd0.11035950190860638, 32'sd-0.0032386067759488392, 32'sd0.00532081027667774, 32'sd0.09935089565222902, 32'sd-0.04827300930021953, 32'sd-0.0162440717426082, 32'sd0.018202743929334114, 32'sd-0.012081199934375614, 32'sd0.05946430610960405, 32'sd0.03226840021143182, 32'sd0.042511405354983885, 32'sd-0.13577987338100972, 32'sd-0.17303433363252252, 32'sd-0.06093606116479907, 32'sd-0.05518923769556337, 32'sd-0.038837155163300746, 32'sd-0.06365731167012538, 32'sd-0.03885112292305976, 32'sd0.12827874132869935, 32'sd0.0249662168344735, 32'sd0.11128126961884989, 32'sd0.1038575282785892, 32'sd0.014664838142823492, 32'sd-0.04029389144868514, 32'sd-0.13269439037150763, 32'sd-0.09524728034606361, 32'sd-0.08968162720612952, 32'sd0.008522032683012581, 32'sd0.12386846128042495, 32'sd0.11126150674137454, 32'sd0.04222336108609481, 32'sd0.05817150293826219, 32'sd-0.00024616484854851715, 32'sd-0.0629957457082253, 32'sd-0.0021499111658095957, 32'sd-0.09803074873375862, 32'sd0.06654310561179964, 32'sd-0.012465335016400927, 32'sd-0.0018318978657832915, 32'sd-0.033964345028699015, 32'sd-0.0557083464006511, 32'sd0.0312927280631541, 32'sd-0.01582118211162683, 32'sd-0.18157788477943335, 32'sd-0.02526881906774847, 32'sd0.11268160079947358, 32'sd0.014903020169796579, 32'sd0.1123328425990131, 32'sd-0.029894837449190907, 32'sd-0.003616652391035702, 32'sd0.07152260017636608, 32'sd-0.14052457435771215, 32'sd-0.12397098342656906, 32'sd-0.12596479334052327, 32'sd-0.12864161791277318, 32'sd-0.09687198196860737, 32'sd-0.06403643158780714, 32'sd0.03258923469628231, 32'sd0.10115909410681849, 32'sd0.05119275864707581, 32'sd0.07775262159703342, 32'sd-0.002351324187596205, 32'sd0.03489398400744897, 32'sd0.014724579264446787, 32'sd0.04369687538533748, 32'sd0.006678198765792538, 32'sd-0.029381235391799227, 32'sd-0.09628716785771001, 32'sd-0.028491775934677218, 32'sd0.003991006859514433, 32'sd0.08045692234345053, 32'sd-0.015004714665958936, 32'sd-0.11821143374840591, 32'sd-0.03111331978335522, 32'sd0.0975710235531829, 32'sd0.10188933165591274, 32'sd0.13763682952008763, 32'sd0.018564301920659238, 32'sd-0.018182702639906952, 32'sd-0.10958370007314829, 32'sd-0.09112431557977292, 32'sd-0.16429713210733288, 32'sd-0.19108667531852133, 32'sd-0.13784799870749362, 32'sd-0.04975473992264369, 32'sd-0.049848982163944844, 32'sd0.04744123478519686, 32'sd-0.08789535668883035, 32'sd0.06732818399250348, 32'sd0.03742284665744786, 32'sd-0.005390547707272964, 32'sd-0.00836856424884894, 32'sd-0.021982021824622847, 32'sd0.1281866495212041, 32'sd-0.07140783887611563, 32'sd-0.11973384428180578, 32'sd0.014193830334795104, 32'sd0.011966763697301144, 32'sd0.0013472593952990077, 32'sd0.0003812750384409616, 32'sd-0.06951151248131578, 32'sd0.04365877056537717, 32'sd0.14238949161682674, 32'sd0.1574643669360101, 32'sd0.2571269597232091, 32'sd-0.04956881193663322, 32'sd-0.021474493299402604, 32'sd0.009009278902542077, 32'sd-0.19843911242777143, 32'sd-0.10808039141273475, 32'sd-0.1265312851782534, 32'sd-0.015227425789442273, 32'sd-0.06053331892869154, 32'sd-0.022967778574862225, 32'sd-0.10972764549030585, 32'sd-0.05054182578757964, 32'sd0.07217587897232643, 32'sd-0.07547293643019454, 32'sd0.14920093309753413, 32'sd0.05515584010355549, 32'sd0.022591541189251156, 32'sd0.044525201305919165, 32'sd-0.07558995628409895, 32'sd0.008623421069436338, 32'sd0.05198020881092431, 32'sd-0.00717121758062524, 32'sd-0.05178984520387974, 32'sd-0.03937067291516721, 32'sd0.02464404305670797, 32'sd-0.03056800457346769, 32'sd0.02581451119484407, 32'sd0.021101885490800897, 32'sd0.038099355205606866, 32'sd-0.1258522638526947, 32'sd-0.004063265394880823, 32'sd-0.17691620045573966, 32'sd-0.11252484019037433, 32'sd-0.015916608557157503, 32'sd0.014740693681453438, 32'sd-0.03588469644603085, 32'sd-0.15945773477098624, 32'sd-0.011380628431425031, 32'sd0.06276855415402958, 32'sd-0.06762275728437937, 32'sd0.02243955854803341, 32'sd0.06277270278728402, 32'sd0.10891668125693264, 32'sd0.09152725029620784, 32'sd-0.11256760504949113, 32'sd0.04558341977683551, 32'sd-0.03067438608944676, 32'sd0.15791177172678686, 32'sd0.03712322485278549, 32'sd-0.02418581344770785, 32'sd-0.09309658667503963, 32'sd0.005249396103983119, 32'sd0.04247551330007323, 32'sd-0.040709465246092195, 32'sd0.07096629007676135, 32'sd0.035228929204666005, 32'sd-0.019637290266649236, 32'sd-0.1856754443045087, 32'sd-0.0975553994121553, 32'sd-0.05116505205067204, 32'sd0.002276768030981138, 32'sd-0.03449857302731682, 32'sd0.02750716927013113, 32'sd-0.1268856086018892, 32'sd-0.1464702485542585, 32'sd0.015557158115866554, 32'sd-0.05121506823684685, 32'sd-0.06311004410844359, 32'sd-0.0629047244914415, 32'sd0.047615151488737545, 32'sd0.06517238308942642, 32'sd0.02301776078138719, 32'sd0.001769355386944472, 32'sd-0.008898672698055452, 32'sd0.09505205579965445, 32'sd0.03273136041888178, 32'sd-0.075820931262847, 32'sd-0.04711626393114394, 32'sd-0.09529672792716894, 32'sd-0.14391592331385214, 32'sd0.03276017724853998, 32'sd0.034086977412071236, 32'sd0.04238810990051544, 32'sd-0.07877336930675993, 32'sd0.0019418329386364903, 32'sd-0.0684600494761205, 32'sd-0.03286023648483285, 32'sd-0.11102850642224754, 32'sd-0.06050024704569323, 32'sd0.02078093846321252, 32'sd-0.08293675891019046, 32'sd-0.07754239003820257, 32'sd-0.026245665156102067, 32'sd-0.044997107038068945, 32'sd-0.06947727593952428, 32'sd-0.11631714559699853, 32'sd-0.03608647272549438, 32'sd-0.049819524851728185, 32'sd-1.4473879059830444e-118, 32'sd0.02823016588819855, 32'sd-0.04232495180318291, 32'sd0.015882017987741838, 32'sd0.0853822492574637, 32'sd0.11630254806498784, 32'sd0.083199282762385, 32'sd0.07192413468236399, 32'sd-0.057040065870848464, 32'sd-0.09251022893980256, 32'sd-0.07716420546725025, 32'sd-0.03250566981658217, 32'sd-0.20111164354239508, 32'sd-0.11876732123624181, 32'sd0.05661182858284434, 32'sd0.06382177812910379, 32'sd-0.03509571824743463, 32'sd0.07407749458725099, 32'sd-0.022723155691767374, 32'sd0.014697893773076905, 32'sd-0.02681405499363281, 32'sd-0.07304917221181839, 32'sd0.07223736928138602, 32'sd-0.07296230407837394, 32'sd-0.032201809087406316, 32'sd-0.0410711239835908, 32'sd-0.138470270728271, 32'sd0.027352305622014822, 32'sd0.0019367933306098778, 32'sd0.07655408062228188, 32'sd-0.021732229895795582, 32'sd0.11881886488871526, 32'sd0.09475766562428853, 32'sd-0.002687976939679576, 32'sd0.06450125662480777, 32'sd0.1495415642574159, 32'sd-0.03516314815423709, 32'sd0.008393481556557702, 32'sd-0.0029002429355669814, 32'sd-0.0970465737607389, 32'sd-0.16550857488451873, 32'sd0.04151458804967703, 32'sd0.12254588198476211, 32'sd0.16070065881319892, 32'sd0.08807822062754546, 32'sd0.0947579768818477, 32'sd0.018541296446233597, 32'sd-0.05020383848241865, 32'sd-0.03139853033340578, 32'sd0.029389747974760145, 32'sd-0.0775087817434077, 32'sd-0.05130061332674683, 32'sd-0.08679595514319106, 32'sd-0.004188888074805703, 32'sd-0.08648341984571832, 32'sd0.0402856767782077, 32'sd0.051503087153500875, 32'sd0.017485098300579996, 32'sd-0.05362525388934133, 32'sd-0.07457318030164402, 32'sd-0.06046887339975177, 32'sd0.14184638154674448, 32'sd0.0970874592626744, 32'sd0.08081569320038579, 32'sd0.03058987662384134, 32'sd0.04680544232989517, 32'sd0.12867846931999133, 32'sd0.10783058836965237, 32'sd0.09041985230787118, 32'sd0.10171480958076948, 32'sd0.1764322670779482, 32'sd0.15841436498011727, 32'sd0.10658758121250235, 32'sd-0.03906547435005339, 32'sd-0.07420940112127411, 32'sd-0.04119843918260694, 32'sd-0.045383448832844876, 32'sd-0.02166048031223406, 32'sd0.04480144738565534, 32'sd0.010048093110581417, 32'sd0.02120032319525028, 32'sd0.006064088078211689, 32'sd-0.08870258632984264, 32'sd0.025643675870351632, 32'sd-7.056576230298974e-127, 32'sd0.005772512573003992, 32'sd0.09386248667845747, 32'sd-0.0835667861449366, 32'sd0.009106863049289255, 32'sd0.05177867853636577, 32'sd0.05306100320384507, 32'sd-0.04369637179490876, 32'sd0.06795010965345154, 32'sd0.03453892251959223, 32'sd0.16381747821582357, 32'sd0.13737229932996348, 32'sd0.03345337269232083, 32'sd0.13433119046187955, 32'sd0.18409285729167205, 32'sd0.05805542391531023, 32'sd0.09376303702536598, 32'sd0.029924786637115453, 32'sd-0.14193313626270124, 32'sd-0.0016090406890895011, 32'sd-0.0522815944976671, 32'sd-0.10679108380236917, 32'sd-0.00803987691809616, 32'sd0.003468993321302173, 32'sd0.08559993193315221, 32'sd0.0017025655260636664, 32'sd-0.044422428699055806, 32'sd0.052531695005801037, 32'sd0.029428840278601157, 32'sd-0.016084072429186653, 32'sd-0.030091734267221205, 32'sd0.09323879831494825, 32'sd-0.03115728334774892, 32'sd-0.008822911950524545, 32'sd0.004618652612372045, 32'sd-0.008839799131126964, 32'sd-0.02823517663617284, 32'sd0.0411010119603656, 32'sd0.15237306453819058, 32'sd0.12702222565909518, 32'sd0.11605458269077588, 32'sd0.12200335934283986, 32'sd-0.04910822370459934, 32'sd0.013938178087736727, 32'sd0.03200426993866665, 32'sd0.005008484310797897, 32'sd-0.11049836781483234, 32'sd-0.04580776085706595, 32'sd-0.10060832624555385, 32'sd-0.05615277769216279, 32'sd0.011992645383606077, 32'sd0.03721639197398034, 32'sd0.07382295042595201, 32'sd-0.03209708184181579, 32'sd-0.0665811975616587, 32'sd0.03495341709614431, 32'sd0.00504058300772057, 32'sd0.023072369391978823, 32'sd0.07431607765535787, 32'sd0.03918645961194888, 32'sd-0.039240326144160606, 32'sd-0.10885466160710214, 32'sd0.0024794242746196808, 32'sd0.03417675530765938, 32'sd-0.08919877112561521, 32'sd0.06235569420860159, 32'sd0.01766184165208322, 32'sd0.08425604354851571, 32'sd0.10805717978443749, 32'sd0.003855763540887928, 32'sd-0.07887990729310133, 32'sd-0.03126627582961521, 32'sd-0.1136499613568829, 32'sd-0.06559882507986939, 32'sd-0.13384335146177662, 32'sd-0.06763982081209341, 32'sd-0.056588825479235626, 32'sd-0.12022417303009805, 32'sd-0.0022587576978160676, 32'sd-0.016773061287021187, 32'sd0.14366500905274038, 32'sd0.03155998242578702, 32'sd0.03572915760345083, 32'sd0.04804076533723673, 32'sd3.28251427708557e-117, 32'sd0.07471823296608415, 32'sd-0.011718516501541286, 32'sd-0.06334070820205495, 32'sd-0.09398836043319314, 32'sd0.04757929490449806, 32'sd-0.034264926526683594, 32'sd-0.018727567466920673, 32'sd0.011771370388167786, 32'sd-0.049123120924190064, 32'sd0.02005284004762965, 32'sd-0.10351815819337652, 32'sd-0.06836475842631505, 32'sd-0.10072209064951834, 32'sd-0.020786609469905556, 32'sd-0.07257331839735143, 32'sd-0.13421328500542984, 32'sd-0.06603553673672738, 32'sd-0.02750733960637849, 32'sd-0.060196387310223316, 32'sd-0.05050439608934748, 32'sd-0.06371194620859683, 32'sd-0.009061746387075496, 32'sd0.10795185672451729, 32'sd-0.013133374751676318, 32'sd0.04935293703388303, 32'sd0.06013870243861404, 32'sd-3.882679277241187e-117, 32'sd8.126088377197979e-122, 32'sd-2.4616192413163733e-126, 32'sd0.05228823326306302, 32'sd-0.08032802189120901, 32'sd0.023425845916209307, 32'sd-0.06503388066385604, 32'sd-0.0235107532513661, 32'sd-0.0776261051157397, 32'sd0.013769212700840482, 32'sd-0.06801752537619819, 32'sd-0.1425116944025395, 32'sd-0.15377729927173253, 32'sd-0.07197427198474217, 32'sd-0.1813998590612236, 32'sd-0.20283328543289716, 32'sd-0.10692353430013153, 32'sd-0.10120769154815996, 32'sd-0.12225197766015544, 32'sd-0.09985825130308289, 32'sd0.010466577075019053, 32'sd0.03793097906243945, 32'sd-0.06699182387693528, 32'sd-0.04952093702746529, 32'sd0.07828860333904596, 32'sd-0.032604004232778816, 32'sd0.007421120287856163, 32'sd-0.018921772324554043, 32'sd-2.815103571382206e-116, 32'sd-3.7300080169309546e-125, 32'sd-1.918045383437931e-117, 32'sd0.03098765399373237, 32'sd-0.05397024433729654, 32'sd0.028248157462845733, 32'sd0.04554033920305324, 32'sd0.04680531788064774, 32'sd0.030454333996823183, 32'sd-0.056110656018455676, 32'sd-0.11539742551929248, 32'sd-0.09159979032965804, 32'sd-0.10973839309362761, 32'sd-0.03606402307719468, 32'sd0.006177515553144524, 32'sd-0.035004259204894736, 32'sd0.10872185486082167, 32'sd0.10978921406758725, 32'sd0.06582931551327405, 32'sd0.008876998876945751, 32'sd0.032355033516991205, 32'sd0.05442988828061477, 32'sd0.05746454680929158, 32'sd0.05775656265270082, 32'sd0.12127937634219844, 32'sd0.04725281927587404, 32'sd-0.06851807734266299, 32'sd0.04990997388031718, 32'sd1.3377427154086586e-124, 32'sd-4.078812983313182e-127, 32'sd-6.947920629345714e-124, 32'sd-3.3322007096936515e-125, 32'sd0.06376135336945699, 32'sd-0.07870430361909574, 32'sd-0.027694092654986853, 32'sd-0.07111312840688705, 32'sd0.021784982551809454, 32'sd-0.0836166111750216, 32'sd0.0015337541527387939, 32'sd0.09322124398562871, 32'sd0.13434109494410928, 32'sd0.07515042892061298, 32'sd-0.007255955838767349, 32'sd0.012668713448367395, 32'sd0.06248150093753211, 32'sd-0.04385189973629942, 32'sd0.015089630878052531, 32'sd0.07620970927924108, 32'sd0.023154180499722333, 32'sd-0.052716029327984956, 32'sd0.05334374221707966, 32'sd-0.02933620988487679, 32'sd-0.0034946523356657777, 32'sd0.0932661530313548, 32'sd0.03445485729583586, 32'sd-6.4911410939951e-116, 32'sd1.0652952002962766e-122, 32'sd-9.897961525592639e-124, 32'sd-7.671974489702012e-127, 32'sd-3.358811002317301e-121, 32'sd4.8702304337648855e-123, 32'sd0.13145992057631614, 32'sd0.09609230505582989, 32'sd0.03699231869131599, 32'sd0.12114051382990669, 32'sd-0.04573359279466512, 32'sd-0.0066878093308640274, 32'sd0.012758672926552953, 32'sd0.06252329824684989, 32'sd0.023162797671434626, 32'sd-0.028010705542555546, 32'sd0.0892768162959857, 32'sd0.03413391476642537, 32'sd-0.023796041820152825, 32'sd-0.029858815230591796, 32'sd0.0634102508290772, 32'sd-0.0072789506781662325, 32'sd-0.012914618944902256, 32'sd0.015448267299122324, 32'sd-0.008017818861084743, 32'sd0.12032247750653152, 32'sd4.522842448022875e-124, 32'sd-2.511928854488254e-116, 32'sd7.3782685172654604e-121, 32'sd-9.374185785449393e-124},
        '{32'sd-3.477242692619497e-117, 32'sd-2.0185124873674316e-126, 32'sd-4.873775820688689e-123, 32'sd2.6169295299208375e-126, 32'sd1.3739400429997796e-121, 32'sd-1.1741558212969823e-122, 32'sd1.0457188749101122e-120, 32'sd-4.219962038897147e-125, 32'sd-3.520535512346625e-116, 32'sd2.699611540182885e-124, 32'sd7.525730271904759e-115, 32'sd-4.223801535953506e-123, 32'sd-0.03648142897605203, 32'sd-0.01657365460388617, 32'sd0.03411457011348185, 32'sd0.02875579503433629, 32'sd1.3437958723168475e-118, 32'sd-7.411054310301624e-123, 32'sd-1.2095266540717311e-118, 32'sd-2.662852995287583e-124, 32'sd1.965665818764761e-116, 32'sd6.144255179514171e-124, 32'sd1.1976884630041019e-116, 32'sd4.0105404098089937e-115, 32'sd-2.2412558823545156e-116, 32'sd-3.8954991297566486e-118, 32'sd3.267333589212258e-119, 32'sd-2.3822336001598457e-126, 32'sd-1.8711938244041266e-126, 32'sd3.7957834244567364e-117, 32'sd-3.199046956449724e-126, 32'sd-4.4947026741471705e-127, 32'sd0.026520166189877143, 32'sd0.05299394004436601, 32'sd-0.017869038099700443, 32'sd0.11472714939349735, 32'sd0.09746975950429537, 32'sd-0.018854074168197874, 32'sd0.04165749134648312, 32'sd-0.0052399196404485805, 32'sd0.0019612142309696568, 32'sd0.07307578875767874, 32'sd0.028354033420078906, 32'sd0.054343509472563396, 32'sd0.030163435727838233, 32'sd0.03940897685706942, 32'sd0.012966659741555562, 32'sd0.06727572158888552, 32'sd0.03614631090116725, 32'sd0.10126349978824647, 32'sd-0.033429029092832074, 32'sd0.02037083206817058, 32'sd1.548469529126592e-127, 32'sd-7.122938301220088e-119, 32'sd2.0423511759742894e-116, 32'sd-1.081657637866519e-121, 32'sd1.7479144036335238e-129, 32'sd-2.0720975785080325e-117, 32'sd0.026026622394072132, 32'sd0.045523358189893746, 32'sd0.03747785215106296, 32'sd0.0754815314948131, 32'sd-0.022581241200460893, 32'sd-0.007220484716775989, 32'sd-0.07492424940995696, 32'sd-0.05069460148273562, 32'sd0.029642561544984916, 32'sd-0.027214155825560967, 32'sd-0.014574122693638442, 32'sd0.02767457581830204, 32'sd0.02687608821365534, 32'sd0.15635930580618132, 32'sd0.02197165465807004, 32'sd0.024788199282363598, 32'sd0.026516238036568874, 32'sd0.05333188771531977, 32'sd0.05471753703750015, 32'sd0.033583870199315066, 32'sd0.06895377970197247, 32'sd-0.006481990931554424, 32'sd-0.00815327546880138, 32'sd0.023567308957369727, 32'sd2.4869533818398363e-114, 32'sd-1.999104032082814e-126, 32'sd-7.461364696959232e-115, 32'sd-2.714600787641247e-124, 32'sd0.05735002097717001, 32'sd-0.034779170817957956, 32'sd0.030824655897125425, 32'sd-0.04901794180638279, 32'sd-0.028587348710541135, 32'sd0.07556680330119198, 32'sd-0.0030210482772530987, 32'sd-0.04232507816316782, 32'sd0.05145276691878036, 32'sd-0.05140479912150212, 32'sd-0.048833954102080225, 32'sd-0.026996097863932516, 32'sd0.009493320647281138, 32'sd0.20467841776304704, 32'sd0.13378105548849123, 32'sd-0.11412539046893953, 32'sd0.027207435999891217, 32'sd-0.09212422185878603, 32'sd-0.004613465635829686, 32'sd-0.004097977527765474, 32'sd-0.04399961233935355, 32'sd-0.002407089976130908, 32'sd0.07504601478149245, 32'sd-0.06414671438080859, 32'sd0.018104134874687476, 32'sd3.33361892677762e-119, 32'sd-6.715729536986545e-118, 32'sd0.06058375880989931, 32'sd0.0003189436047792421, 32'sd0.08089289107940495, 32'sd0.019611973977625957, 32'sd0.013338760559601922, 32'sd0.07739484162062656, 32'sd0.03648377966507605, 32'sd0.007762669381266766, 32'sd0.13440256407831278, 32'sd0.12963389650858004, 32'sd0.03433363280605942, 32'sd0.0777600367488986, 32'sd0.02535015031525976, 32'sd-0.03871416361720597, 32'sd0.08130730766730672, 32'sd0.07697052646299796, 32'sd0.04923312388230753, 32'sd0.1053665476318021, 32'sd0.08008439654664427, 32'sd-0.014871572225222205, 32'sd-0.04398121497749119, 32'sd-0.13655947242979777, 32'sd-0.09352134907137306, 32'sd-0.05871639830381244, 32'sd-0.03512224559533553, 32'sd-0.012258491193488099, 32'sd0.06195546396611099, 32'sd-7.546812372083381e-121, 32'sd0.02110949231471161, 32'sd-0.018212772816154344, 32'sd-0.004214810372791463, 32'sd0.008726476755563796, 32'sd0.038114078039292724, 32'sd-0.015927639667880158, 32'sd-0.010990151527358487, 32'sd0.05623082151429045, 32'sd0.04988342643313723, 32'sd0.06024215898210148, 32'sd-0.020181504291306215, 32'sd0.009981055548525589, 32'sd0.07612822434069433, 32'sd0.06271427194642244, 32'sd0.0004946759950528454, 32'sd0.04682627972364607, 32'sd-0.008761257974321819, 32'sd-0.005874321924282766, 32'sd-0.046598901456881975, 32'sd0.019264330271392113, 32'sd0.046927616796142, 32'sd-0.09327819154862402, 32'sd-0.015506984156895274, 32'sd0.06023930753307117, 32'sd0.03643727663858913, 32'sd-0.07793437400788568, 32'sd0.009067657096028286, 32'sd7.887502541178245e-122, 32'sd0.07100101852614284, 32'sd-0.04580926297555348, 32'sd0.009147260028611166, 32'sd0.03621159661185009, 32'sd0.006857531978022209, 32'sd-0.028446985238508447, 32'sd-0.01970550272767355, 32'sd0.07638949266095513, 32'sd0.02130715302989626, 32'sd-0.06373744958879922, 32'sd-0.051691006580240964, 32'sd-0.03312012359026648, 32'sd-0.034918320283348854, 32'sd0.06006426647340255, 32'sd0.03229147951022178, 32'sd0.15615328886077862, 32'sd0.1492929697804066, 32'sd-0.07285133263229625, 32'sd0.039805696958249426, 32'sd-0.06105398280797435, 32'sd-0.07239543904066084, 32'sd0.057013323139607865, 32'sd0.08521716307961781, 32'sd0.01888172409682543, 32'sd-0.02152421260865043, 32'sd0.03472643105274356, 32'sd-0.03535402387237869, 32'sd0.035410625515264874, 32'sd0.0028675979525765102, 32'sd0.04896091038844017, 32'sd0.04035343797684026, 32'sd0.005204703975676596, 32'sd0.044538257025210706, 32'sd0.07599452479840592, 32'sd0.015733921567902178, 32'sd0.02871208308998989, 32'sd0.07277836649629828, 32'sd0.0036584215017914216, 32'sd-0.044644985242288375, 32'sd0.03720794289421648, 32'sd-0.07860163893425591, 32'sd0.01403584382959981, 32'sd0.058914083927021105, 32'sd0.12417581404019529, 32'sd0.1491218625292986, 32'sd0.011602647334951323, 32'sd0.05614008486418909, 32'sd0.003050023673529745, 32'sd0.06943355895118876, 32'sd-0.046199703321215785, 32'sd0.053830235780594725, 32'sd0.05768693491149622, 32'sd0.052125864333133605, 32'sd0.08138942225188313, 32'sd-0.011132184377990422, 32'sd0.037990712566146834, 32'sd-0.0023238583173797946, 32'sd0.08638095434675647, 32'sd0.13386649561501401, 32'sd-0.019129272201725833, 32'sd0.09265701266309155, 32'sd-0.05099760839745371, 32'sd0.003590154517022547, 32'sd0.11662083181119644, 32'sd0.11006578961332132, 32'sd0.10196578332325985, 32'sd-0.03562870618318139, 32'sd-0.11172761412669166, 32'sd-0.02257037199200132, 32'sd-0.0182769125006313, 32'sd0.11230362023689615, 32'sd-0.07691156665618155, 32'sd0.025571932929296128, 32'sd0.016404512888721568, 32'sd-0.044063081336106605, 32'sd-0.07759471653914556, 32'sd-0.004452346670554568, 32'sd0.08037292142241124, 32'sd0.13710922950593737, 32'sd0.1318558631465259, 32'sd0.01057893217897168, 32'sd0.09031224469598627, 32'sd-0.0030283450986779933, 32'sd0.08761909467226629, 32'sd0.021897989591643883, 32'sd-0.005891760200467447, 32'sd-0.07320097299042631, 32'sd0.027057579035351196, 32'sd0.03441898758433214, 32'sd0.052085239665055065, 32'sd-0.00043138033430278807, 32'sd0.1974276666820939, 32'sd0.07072685098465584, 32'sd0.1210195373720733, 32'sd-0.03423379684034479, 32'sd0.029737802180379694, 32'sd-0.01415840165742089, 32'sd-0.09503520694317004, 32'sd-0.11792322233058856, 32'sd-0.1809444659626263, 32'sd-0.009428768564116147, 32'sd-0.14130007853560655, 32'sd-0.07965992397316266, 32'sd-0.0432905558065728, 32'sd-0.0427504020718195, 32'sd0.05811996822736475, 32'sd0.014354741748244653, 32'sd0.07123729830199471, 32'sd0.05248118161930433, 32'sd-0.012104051921171241, 32'sd-0.06824878355762215, 32'sd0.09512365088953137, 32'sd0.06005760571109896, 32'sd-0.06989504939214748, 32'sd0.07226913296800676, 32'sd0.06083386460401492, 32'sd-0.0028567974741223585, 32'sd-0.029183139353550054, 32'sd0.022927574873215846, 32'sd0.10927598304901256, 32'sd0.15620604762629955, 32'sd-0.017942207410257097, 32'sd0.00847335438743463, 32'sd-0.02029656881674052, 32'sd-0.10074288658802269, 32'sd-0.041459462208671555, 32'sd-0.10176875259734038, 32'sd-0.10443950742425949, 32'sd-0.11040792439046661, 32'sd-0.016565288600978816, 32'sd-0.05125679634398477, 32'sd0.03611976280311306, 32'sd-0.043903152520281236, 32'sd-0.08357162234187258, 32'sd-0.08043594856734443, 32'sd-0.07099635286550156, 32'sd-0.03550986955030134, 32'sd0.03715662489547382, 32'sd0.040805318920623807, 32'sd0.0059587223132348864, 32'sd0.030143341005737297, 32'sd-0.015314626817745352, 32'sd-0.01765081840281666, 32'sd0.08119544144898194, 32'sd0.029520569904632036, 32'sd-0.0032085415463062017, 32'sd0.014050076401743425, 32'sd0.047919577375390425, 32'sd0.0630026767559998, 32'sd0.16096945490922107, 32'sd0.0967642096187233, 32'sd0.13615724061711681, 32'sd0.14708745348169783, 32'sd0.11107472157844744, 32'sd0.13111440295956378, 32'sd-0.019738565142625265, 32'sd-0.033351566706019194, 32'sd0.056428018676609966, 32'sd0.03185875327387227, 32'sd-0.04920696547981458, 32'sd-0.11312451111882028, 32'sd-0.16171266903180698, 32'sd-0.19085949156653836, 32'sd-0.045015220460918146, 32'sd-0.10735929000115771, 32'sd-0.023251185035798285, 32'sd-0.020764590376697107, 32'sd0.014423394382868394, 32'sd0.05681079131034717, 32'sd-0.037006247414525156, 32'sd-0.09220125500501435, 32'sd-0.05624308847190595, 32'sd0.050023688722357317, 32'sd0.00405455381955783, 32'sd-0.034061750819904396, 32'sd0.08615155429978315, 32'sd0.016291842907029154, 32'sd0.19376101871101384, 32'sd0.2237732172982304, 32'sd0.1980963970019457, 32'sd0.2569308266259759, 32'sd0.24713318511042898, 32'sd0.14406072757647811, 32'sd0.06759450594832767, 32'sd0.1242562047812734, 32'sd0.16031034630872434, 32'sd0.058492551296822015, 32'sd-0.023760100560635274, 32'sd-0.07657480944263328, 32'sd-0.057185059140231594, 32'sd-0.07719554560656768, 32'sd-0.23502716134104212, 32'sd-0.12644885684810994, 32'sd-0.06316325886212606, 32'sd-0.013638933994331347, 32'sd0.005949864366082809, 32'sd-0.06238004006098422, 32'sd-0.1405271917403722, 32'sd-0.007775833764648512, 32'sd-0.038037786232006, 32'sd-0.059303409925355, 32'sd-0.07434865930493252, 32'sd0.011507056514847139, 32'sd0.0591603306207715, 32'sd0.03180231573775952, 32'sd0.07811479356754529, 32'sd0.19077073500612424, 32'sd0.23571219493652001, 32'sd0.2994164553876432, 32'sd0.32697747826274326, 32'sd0.1699104657401061, 32'sd0.10322290343030924, 32'sd0.08821092582559358, 32'sd0.17017523053582598, 32'sd-0.028594738511522055, 32'sd0.025640976273879977, 32'sd-0.0030338254874056306, 32'sd0.06572601377270224, 32'sd0.00798255096358161, 32'sd-0.09326522533463077, 32'sd-0.005125351219593003, 32'sd-0.044077876531979664, 32'sd0.037573196565635666, 32'sd0.12570376576721315, 32'sd0.03150049966000265, 32'sd0.01772510669902862, 32'sd-0.08946150425691447, 32'sd-0.1438395510828036, 32'sd-0.15190644541975637, 32'sd-0.22078099616703573, 32'sd-0.027539377675696655, 32'sd-0.008622293040959765, 32'sd-0.11402079490642271, 32'sd0.0643731185341548, 32'sd0.028390263537467684, 32'sd0.1408280689532854, 32'sd0.124922573237702, 32'sd0.14791901187918963, 32'sd0.09525950310182422, 32'sd0.06736616017452604, 32'sd0.06221939116854706, 32'sd-0.008966624582280692, 32'sd-0.09326780059538149, 32'sd-0.07762153117281273, 32'sd-0.013172633163123695, 32'sd0.06259622898454158, 32'sd0.03613866043190199, 32'sd0.08357551658760831, 32'sd0.0016441400279855838, 32'sd-0.03504277745607134, 32'sd0.009660091491643725, 32'sd0.09627913691481796, 32'sd0.017159483155808515, 32'sd0.03945690274509654, 32'sd-0.02312203814249892, 32'sd-0.13589064154554334, 32'sd-0.22059684092468754, 32'sd-0.24836440169276075, 32'sd-0.23996354101834566, 32'sd-0.11314054140606689, 32'sd-0.2081581560041711, 32'sd-0.17385991796980008, 32'sd-0.0162835193768688, 32'sd0.043017784396461194, 32'sd0.05873447926619883, 32'sd0.023901831778662844, 32'sd0.05695810878214592, 32'sd0.04545814730554842, 32'sd0.023595810569981744, 32'sd0.037140231604799664, 32'sd0.0028250772287623876, 32'sd-0.018731492956980216, 32'sd-0.008940800948168327, 32'sd0.019634298304239566, 32'sd0.12314575475814353, 32'sd0.11271338765242862, 32'sd0.03132939693162863, 32'sd-0.02856333832808757, 32'sd0.05696851547060807, 32'sd0.006365821277852312, 32'sd-0.03495918334370396, 32'sd-0.039546392002790504, 32'sd0.12335219405902784, 32'sd-0.02820991062021229, 32'sd-0.12156272990446985, 32'sd-0.15169266419754876, 32'sd-0.20548635985261887, 32'sd-0.2512660573138938, 32'sd-0.3482517117841147, 32'sd-0.35082350962587083, 32'sd-0.3024915742081012, 32'sd-0.169121845679589, 32'sd-0.10878076851788464, 32'sd-0.06380666069056273, 32'sd-0.029160337634271307, 32'sd-0.045828664949766756, 32'sd0.09668283166597354, 32'sd0.03653521065887391, 32'sd0.0527550029151544, 32'sd0.047931143953145815, 32'sd-0.01037613665865112, 32'sd0.0039140475833630535, 32'sd0.04954307744124245, 32'sd0.06926755628575183, 32'sd-0.027400343370405374, 32'sd0.014813451610770823, 32'sd0.03688020715276546, 32'sd-3.1402892888690865e-125, 32'sd0.06618729495706244, 32'sd-0.06396484390402374, 32'sd0.04579343976404223, 32'sd-0.06400686684775965, 32'sd-0.06244991883177602, 32'sd0.03326127269443515, 32'sd-0.0004541357882051851, 32'sd-0.08966441284973319, 32'sd-0.2494011398836781, 32'sd-0.3558351994736395, 32'sd-0.3419683945456833, 32'sd-0.43892912846271037, 32'sd-0.300826490430584, 32'sd-0.17291642958023934, 32'sd-0.1472278735286963, 32'sd-0.08141708642757696, 32'sd-0.04805972228816878, 32'sd-0.08383466198745615, 32'sd0.05627928763682477, 32'sd-0.026211897459341806, 32'sd-0.016033342731406594, 32'sd-0.060194715548882866, 32'sd0.10218695676459225, 32'sd0.021086623750061442, 32'sd0.0387011892185021, 32'sd0.032121422611364414, 32'sd-0.01223715201132818, 32'sd0.005818567278949022, 32'sd-0.035828200271352945, 32'sd0.06900180742673537, 32'sd0.14765869341604856, 32'sd0.09470913166121066, 32'sd0.04813717841760039, 32'sd0.08554851179648491, 32'sd0.04412124471423637, 32'sd-0.05948147057193002, 32'sd-0.09864395181862776, 32'sd-0.1751072006196919, 32'sd-0.19175529770894834, 32'sd-0.2917235581496368, 32'sd-0.27851768569648877, 32'sd-0.17996604431733285, 32'sd-0.18220829498439564, 32'sd0.06475101648666118, 32'sd0.023685564040665366, 32'sd-0.035134144705381336, 32'sd0.08517714579171858, 32'sd0.005081554700450875, 32'sd0.09701241718171742, 32'sd-0.07876829744318897, 32'sd-0.006546218077482004, 32'sd0.04579604157017356, 32'sd-0.04527423335338605, 32'sd-0.034246184562825736, 32'sd0.026622761747820172, 32'sd0.050237680338732674, 32'sd0.023726142282805868, 32'sd0.04668946625569503, 32'sd0.029529229190090423, 32'sd0.10000570687564879, 32'sd0.14041109940747898, 32'sd0.12131846895048361, 32'sd0.0864574992029198, 32'sd0.07728809277121443, 32'sd0.03052310337486688, 32'sd0.14646767117754664, 32'sd0.021692720947221297, 32'sd-0.10845524672094173, 32'sd-0.1982656542002885, 32'sd-0.09463356591574913, 32'sd-0.10987519594906225, 32'sd-0.05368886267947701, 32'sd-0.06051936941980772, 32'sd-0.0985595904829608, 32'sd0.08305476785852826, 32'sd-0.08575051727673423, 32'sd0.027116365139294763, 32'sd0.0057626559089970514, 32'sd0.028705346249510842, 32'sd0.08765343562683853, 32'sd-0.037036358225220736, 32'sd-0.11813944587152224, 32'sd-0.1550189008991575, 32'sd2.9064866306693084e-114, 32'sd-0.026387213969299002, 32'sd-0.006786365633438644, 32'sd0.08509929902200679, 32'sd0.06547603036145942, 32'sd0.06102503802656112, 32'sd0.017901563720942235, 32'sd-0.0036844955601666113, 32'sd0.024435071300022308, 32'sd0.07423968249038543, 32'sd0.18288436417791312, 32'sd0.11864184840956489, 32'sd0.03146535795506582, 32'sd-0.09267538161237981, 32'sd-0.045630451868057996, 32'sd0.0021417450675088948, 32'sd-0.035178049049025814, 32'sd-0.001124469598253854, 32'sd-0.049265671839367725, 32'sd0.05417398213473842, 32'sd-0.09647104863437346, 32'sd0.018457266562591997, 32'sd0.053834254322259016, 32'sd0.009047968004925354, 32'sd0.039463196313359775, 32'sd-0.07004919677589733, 32'sd-0.032212338428825045, 32'sd0.04668054199687487, 32'sd0.07371476109643552, 32'sd0.03434206384157841, 32'sd0.027962866322340074, 32'sd-0.08207378272098098, 32'sd0.04898063331432199, 32'sd0.16373393043314202, 32'sd0.07484737034132481, 32'sd0.058205643597262394, 32'sd0.026794832487325865, 32'sd0.028944337285051566, 32'sd0.05199870908542038, 32'sd0.1122997616175464, 32'sd0.08374056554398913, 32'sd0.11799200792863081, 32'sd0.1143329759982561, 32'sd0.07186264086253423, 32'sd-0.03228699499391349, 32'sd0.0037913737280412083, 32'sd-0.07425379449296032, 32'sd0.01776214138657098, 32'sd0.0719241339489808, 32'sd0.05942179086436773, 32'sd-0.10355249718075993, 32'sd-0.08936019837891301, 32'sd0.021939147365192226, 32'sd-0.18372387842474497, 32'sd-0.04609335335108103, 32'sd0.019248761831143796, 32'sd0.11595584641760213, 32'sd0.11594896470597425, 32'sd0.028516301996037663, 32'sd0.06642692959870461, 32'sd0.0004996046986259475, 32'sd-0.06814691778510355, 32'sd0.06765738875196718, 32'sd-0.03198647075282659, 32'sd0.0780952983448219, 32'sd-0.08271482994479931, 32'sd0.11346558383944087, 32'sd0.07290524117493549, 32'sd-0.08779458556285484, 32'sd-0.0416423574430474, 32'sd0.10817729129109732, 32'sd-0.05237384017562029, 32'sd0.06615131791008519, 32'sd0.0941953373832362, 32'sd0.0066273377779726686, 32'sd-0.027438334937606286, 32'sd-0.005996611984887435, 32'sd0.002811480725359037, 32'sd-0.22904617427606316, 32'sd-0.0671512235588067, 32'sd-0.01879659183331042, 32'sd-0.03375454979789127, 32'sd0.05250202945060339, 32'sd0.0056312568224511856, 32'sd-1.3201975123513495e-127, 32'sd0.05974662875142926, 32'sd-0.08267639183355949, 32'sd-0.010773510447949221, 32'sd0.01201109901716502, 32'sd-0.11289086261945466, 32'sd-0.016684183720763954, 32'sd-0.06237613927036503, 32'sd-0.026696780978693067, 32'sd-0.08404886412814325, 32'sd0.11553636425140612, 32'sd-0.036924989812056934, 32'sd-0.048801988723373345, 32'sd0.02353498547431077, 32'sd-0.039452256771390415, 32'sd0.061769773058257926, 32'sd0.09216668916648137, 32'sd-0.01351482282959261, 32'sd-0.028960368571953287, 32'sd-0.016538585821391935, 32'sd-0.05954022999718739, 32'sd-0.04315649410809082, 32'sd-0.05828863599415801, 32'sd0.010931594265618957, 32'sd0.08722990607406207, 32'sd-0.10354776533639183, 32'sd-0.01984462641991149, 32'sd-3.447301265198121e-127, 32'sd3.6622157513252956e-116, 32'sd3.3672648459077895e-120, 32'sd0.025263679681478003, 32'sd-0.052940606988583286, 32'sd0.09880960844345421, 32'sd-0.08532701004556492, 32'sd-0.06394650369221122, 32'sd0.06789289643428614, 32'sd-0.04590006529877315, 32'sd0.008995592637630867, 32'sd0.03472526797785859, 32'sd-0.006209139372187869, 32'sd0.03786330152437081, 32'sd-0.035708816042111256, 32'sd-0.19508977952835324, 32'sd-0.13860942871315723, 32'sd-0.0781462494599276, 32'sd-0.0837106931885282, 32'sd-0.10957612477429186, 32'sd-0.0054662131641575636, 32'sd-0.022157251833657205, 32'sd-0.009061314047759889, 32'sd-0.06480119843838898, 32'sd-0.05859376905643204, 32'sd-0.029827019347181603, 32'sd0.030425412421556088, 32'sd0.04458202573339144, 32'sd8.345998510458716e-125, 32'sd1.0442009025415857e-118, 32'sd8.150631249057142e-122, 32'sd0.090192766510919, 32'sd0.010100912808287548, 32'sd0.02447036957506849, 32'sd0.024507796623843038, 32'sd0.024854619304705564, 32'sd0.06940051670315793, 32'sd-0.04120828724050143, 32'sd-0.07033206949621638, 32'sd0.08428403710070331, 32'sd0.010336756907988093, 32'sd-0.006256937201430679, 32'sd0.025036884213221627, 32'sd-0.05006120774067598, 32'sd0.003545495274661686, 32'sd-0.0006711191402803267, 32'sd-0.05357892840665055, 32'sd-0.11217325085145727, 32'sd-0.14275791389039397, 32'sd0.009114682611073892, 32'sd0.004745344149592349, 32'sd-0.04755354776492167, 32'sd-0.08441197449577612, 32'sd-0.0460996013403341, 32'sd0.03379416305539226, 32'sd0.05549811943423623, 32'sd8.445526238840428e-118, 32'sd-1.07172663232117e-124, 32'sd-5.886806102922042e-126, 32'sd-1.2254397992870769e-120, 32'sd0.020667014507004318, 32'sd-0.006924701476749723, 32'sd0.0015293394669371634, 32'sd-0.00026905282861521007, 32'sd-0.007871019615567285, 32'sd0.031194483765748106, 32'sd0.03471644895991704, 32'sd0.050306034584244784, 32'sd0.0351310469166218, 32'sd0.021487493158558538, 32'sd0.06993148739953589, 32'sd0.06523177227445699, 32'sd0.0773175866418861, 32'sd-0.07036849863479958, 32'sd0.02992632974656536, 32'sd0.011401608450851648, 32'sd-0.02798886650663126, 32'sd-0.0728364287343483, 32'sd-0.004727014541143725, 32'sd-0.0595093833053073, 32'sd-0.009773268047910231, 32'sd0.04405871888428915, 32'sd0.032386067423875786, 32'sd1.254370818666142e-117, 32'sd1.5702685678795054e-115, 32'sd5.22837388735086e-118, 32'sd9.605532891759007e-117, 32'sd2.3130852324648422e-116, 32'sd1.078101401789441e-124, 32'sd0.07156015123384092, 32'sd0.06873043965362136, 32'sd-0.032658627891903075, 32'sd0.044589179998784326, 32'sd-0.01278170303442059, 32'sd0.04036464104589306, 32'sd-0.07440453837191448, 32'sd-0.059642213478470464, 32'sd-0.08106778037750076, 32'sd-0.018636351308788095, 32'sd0.04304440963296295, 32'sd0.00842489473875775, 32'sd0.012678007395769192, 32'sd-0.018646760865046894, 32'sd0.03429336103675363, 32'sd0.05927684011759005, 32'sd-0.03253018363072109, 32'sd-0.11172201231042356, 32'sd-0.06206295282274195, 32'sd0.03747227300998327, 32'sd-1.584146652668533e-116, 32'sd2.962292953990268e-119, 32'sd-3.6605998123080713e-121, 32'sd2.862858885081884e-118},
        '{32'sd-1.3419947652016758e-122, 32'sd1.0050187121834812e-121, 32'sd3.878231080613774e-126, 32'sd2.3363136256367065e-126, 32'sd2.779349193947822e-118, 32'sd-8.362772630876036e-125, 32'sd-6.278178803478572e-121, 32'sd-3.1758935892227785e-120, 32'sd2.1140303926551802e-117, 32'sd3.9918303421227577e-119, 32'sd3.1036068412683006e-121, 32'sd-3.9612267534364424e-126, 32'sd0.027795984415942786, 32'sd0.015662578701695865, 32'sd0.09619648011589811, 32'sd0.08423139249376625, 32'sd1.2060130601259977e-122, 32'sd-2.421936077295073e-126, 32'sd-7.490161261533612e-125, 32'sd6.452202541601295e-126, 32'sd-2.9355529527705965e-130, 32'sd-1.510498630184925e-122, 32'sd-7.688719753661087e-121, 32'sd-4.84973787285158e-121, 32'sd-6.950774221823396e-124, 32'sd-1.9322070871934572e-126, 32'sd-1.162214352406956e-127, 32'sd-3.640436271922309e-116, 32'sd7.256489121717295e-117, 32'sd7.952654726432286e-127, 32'sd-4.526215943943083e-126, 32'sd1.2086119688186003e-122, 32'sd-0.004456415181654508, 32'sd-0.04636526034801871, 32'sd-0.009933106695360861, 32'sd-0.024964609452115972, 32'sd-0.08588714868347193, 32'sd0.0820164633677558, 32'sd0.09786085524095324, 32'sd-0.02322009443653721, 32'sd0.02391697791765199, 32'sd-0.031020526708695893, 32'sd0.04832045233971031, 32'sd-0.04559865359418065, 32'sd0.09292490925847913, 32'sd0.01762784813360713, 32'sd0.05775784524688551, 32'sd-0.03158735284445378, 32'sd0.004162765153744838, 32'sd0.0834608870855051, 32'sd0.06401354653002127, 32'sd0.06400448994042054, 32'sd-6.676372495297107e-115, 32'sd-2.8800127491534197e-127, 32'sd-1.1907029022157518e-122, 32'sd1.5483544813718301e-117, 32'sd-3.776456953642889e-119, 32'sd1.6786432896778465e-125, 32'sd0.04503756790685395, 32'sd-0.04751229830981349, 32'sd0.021332409726793528, 32'sd0.0627601425527849, 32'sd-0.008126517849405402, 32'sd-0.037540771895822674, 32'sd-0.007077204000210168, 32'sd0.0032168442702137563, 32'sd0.028991295985164253, 32'sd0.048579780171348175, 32'sd0.0779373219459736, 32'sd0.02620421086356817, 32'sd0.0017819406597253107, 32'sd-0.032467124237580774, 32'sd-0.03633775167455115, 32'sd0.0312669283102657, 32'sd-0.055322437196293824, 32'sd-0.0687357853574719, 32'sd0.03726421420676468, 32'sd-0.031684067902264225, 32'sd0.033138616292573315, 32'sd0.03767364701301535, 32'sd0.01703442700336189, 32'sd0.005804520565030522, 32'sd-1.195762825945955e-118, 32'sd1.0934844011544629e-116, 32'sd-1.2431323241644055e-121, 32'sd2.7208547981459155e-120, 32'sd0.006992501631980674, 32'sd-0.02910952049800568, 32'sd0.09732173124515894, 32'sd-0.013221736861187152, 32'sd0.01232387867672972, 32'sd-0.06346254847724346, 32'sd0.03621662349181246, 32'sd0.004081550349779069, 32'sd0.04303118719699069, 32'sd0.06783349149055103, 32'sd-0.020712449333781267, 32'sd0.11508748906503179, 32'sd-0.05618697998007979, 32'sd-0.062066784359042976, 32'sd0.09016414728545925, 32'sd0.022968862060595233, 32'sd-0.025672902148927753, 32'sd-0.004518166780331907, 32'sd-0.004265897361623669, 32'sd-0.025102989269875326, 32'sd-0.1376862055850369, 32'sd-0.017135479202262882, 32'sd0.03547182188718926, 32'sd0.04418309783181567, 32'sd0.07308927655770668, 32'sd-2.7114097586143954e-127, 32'sd-2.4760509880053985e-126, 32'sd0.04350130377885425, 32'sd0.03590482050108953, 32'sd-0.12200810098649871, 32'sd-0.006625206688588051, 32'sd0.004004498106256888, 32'sd0.08734350886064024, 32'sd0.1226217105409828, 32'sd0.027125622740042318, 32'sd0.056749849979037176, 32'sd-0.1392857037068215, 32'sd0.030035256428256097, 32'sd0.04404715683855134, 32'sd0.12963185619968287, 32'sd0.1254975762023525, 32'sd0.07917748609733237, 32'sd0.013022836199900877, 32'sd-0.009299156979927474, 32'sd0.06025864164477023, 32'sd0.08300119438539857, 32'sd-0.01970458872191762, 32'sd-0.03268776805076343, 32'sd-0.0380563669713052, 32'sd-0.018052835090084846, 32'sd0.03536170700539967, 32'sd-0.09947029464260781, 32'sd0.03865058258944713, 32'sd0.025481398794388276, 32'sd-1.068790933158732e-124, 32'sd0.055688032998657655, 32'sd-0.033472449727533216, 32'sd0.08321630403027089, 32'sd0.07161241436960492, 32'sd0.004388193522394649, 32'sd0.09993419885075802, 32'sd-0.013861652220409441, 32'sd0.03691259312679272, 32'sd-0.03558539888731841, 32'sd-0.046000591230872516, 32'sd-0.012154132191176727, 32'sd0.12252063151307199, 32'sd0.11691597842017941, 32'sd0.10128653230551707, 32'sd0.08400315762821561, 32'sd0.112100739457109, 32'sd-0.09552923843767529, 32'sd-0.06830247929427921, 32'sd-0.11029350162280045, 32'sd-0.04119658677779408, 32'sd-0.03638305738088785, 32'sd0.0036146460239594156, 32'sd-0.11050604110805684, 32'sd-0.060030477313543766, 32'sd-0.0003970574617476147, 32'sd0.0033729836738857883, 32'sd0.0347369316896328, 32'sd-3.3153849242909805e-120, 32'sd0.0073475321728557665, 32'sd-0.02282592995804063, 32'sd0.08059208826960745, 32'sd-0.04988447282336696, 32'sd-0.08435315864453283, 32'sd0.023278579225864984, 32'sd-0.0849819383275474, 32'sd-0.02788144201697946, 32'sd0.03975868920694631, 32'sd0.12434464757062764, 32'sd0.017590201972190824, 32'sd0.07685170980862562, 32'sd0.11807827993079516, 32'sd0.016881298952578942, 32'sd0.1543063429815887, 32'sd0.12314036601817653, 32'sd0.008675488731425965, 32'sd-0.013372377364876864, 32'sd-0.04055626119254971, 32'sd-0.02867629004088023, 32'sd0.10702959251395606, 32'sd0.022603746110433517, 32'sd-0.06313549369471688, 32'sd0.031397183551716876, 32'sd0.0033438993263256965, 32'sd-0.014571896488774636, 32'sd-0.03738444734481455, 32'sd0.07774403394330001, 32'sd0.013777206408152633, 32'sd0.0047508377684596335, 32'sd0.10745677727972316, 32'sd0.11309745076410546, 32'sd0.03377078992671206, 32'sd0.009573443503955201, 32'sd0.03494482249536596, 32'sd-0.039928267209327406, 32'sd0.06618437309494216, 32'sd0.07395048553118287, 32'sd0.14002940918220338, 32'sd0.07472397152915067, 32'sd0.12876536660979473, 32'sd0.10164992659890254, 32'sd0.05947708019124364, 32'sd0.18276440756075416, 32'sd0.04946142446767393, 32'sd-0.01924264873218031, 32'sd-0.002297408423491768, 32'sd-0.02343582130240775, 32'sd-0.05829075481169398, 32'sd-0.06317112581609302, 32'sd-0.05191356412050623, 32'sd-0.0014132313311884656, 32'sd0.06239453349694722, 32'sd0.06080673626371456, 32'sd-0.0019238550164045287, 32'sd0.06193726563764709, 32'sd-0.05154982589249265, 32'sd0.07549882573988231, 32'sd0.052931084091832774, 32'sd-0.08409871798478408, 32'sd-0.012021936875772762, 32'sd-0.03325002400707797, 32'sd0.03802871219366381, 32'sd-0.08409296596364647, 32'sd-0.02194708392611308, 32'sd0.04313163384500568, 32'sd0.09101828814914273, 32'sd0.02424883930230694, 32'sd0.06366259219973136, 32'sd0.16495976559089956, 32'sd0.04782519520649796, 32'sd0.1470829753987045, 32'sd0.19488926886056746, 32'sd-0.04265829336089936, 32'sd0.03923383114954115, 32'sd-0.017255233727938805, 32'sd0.020163388569891513, 32'sd-0.04232613169781721, 32'sd0.04352573970144394, 32'sd0.01914043687374044, 32'sd-0.00023124377602465953, 32'sd0.0953978995758277, 32'sd0.05375847333544114, 32'sd0.048415366199983184, 32'sd-0.11907168374261064, 32'sd0.07385189976662572, 32'sd-0.006238404165774049, 32'sd0.003992996109986929, 32'sd0.08300134829873268, 32'sd-0.05696215614652349, 32'sd0.004868795358057076, 32'sd-0.05585050288289539, 32'sd0.006198741035884341, 32'sd0.03588416288892444, 32'sd-0.15000008689711622, 32'sd-0.03796263262599589, 32'sd-0.08082394323234601, 32'sd-0.03392131491139033, 32'sd0.06552243821426564, 32'sd0.08945590889113868, 32'sd0.11777313224051729, 32'sd0.16143125544101264, 32'sd0.06526198651069105, 32'sd-0.047841174770473956, 32'sd-0.10233015362595538, 32'sd-0.03279974488015856, 32'sd0.07105698449944979, 32'sd-0.0731907786744982, 32'sd0.044305536408049996, 32'sd-0.05542611430942461, 32'sd0.06350677460639799, 32'sd-0.054373076349461986, 32'sd0.010264648997444838, 32'sd0.08714171708881685, 32'sd0.15198887985321885, 32'sd0.04699394746093852, 32'sd0.11197885171086205, 32'sd0.03751311581163699, 32'sd0.05644793990147233, 32'sd-0.004397102683663251, 32'sd-0.08189405827297469, 32'sd-0.056563091533410846, 32'sd-0.09040631185249642, 32'sd-0.09723939234262578, 32'sd-0.13458110534918108, 32'sd-0.21224993101662498, 32'sd-0.18634871995952837, 32'sd0.0957934093030019, 32'sd0.19363128992131476, 32'sd0.1007300112433236, 32'sd-0.055880877145492044, 32'sd-0.09551257747827752, 32'sd0.04110620940327627, 32'sd-0.07445110578561007, 32'sd0.033034919844108834, 32'sd0.002984690407137853, 32'sd0.028963763417632387, 32'sd-0.07141876287335472, 32'sd-0.09827251143788324, 32'sd-0.07675476278977962, 32'sd-0.017033523308116184, 32'sd-0.026703441447137072, 32'sd0.02915594380827704, 32'sd0.04747875045324987, 32'sd-0.018583878416487367, 32'sd-0.05120972035911011, 32'sd0.06951440259966572, 32'sd-0.024001126006311185, 32'sd-0.033887371664656794, 32'sd-0.07188277118120767, 32'sd-0.11303510480658137, 32'sd-0.07220947526252268, 32'sd-0.15799944432277585, 32'sd-0.3031794138152739, 32'sd-0.057404572020484344, 32'sd-0.024466221167464938, 32'sd0.1321784848352404, 32'sd0.09784417474324673, 32'sd-0.028116699455009192, 32'sd-0.03289073664688484, 32'sd-0.024218079165347264, 32'sd-0.09446229408568116, 32'sd-0.022430608702108484, 32'sd-0.10311759192997437, 32'sd-0.07513244166134225, 32'sd-0.04026031664707133, 32'sd-0.0030701793835453232, 32'sd0.06351706246585875, 32'sd0.03487734601821379, 32'sd0.022639118837499903, 32'sd-0.08173644924199992, 32'sd-0.08818375903764789, 32'sd-0.07369785300106493, 32'sd0.0029407417252393275, 32'sd0.030311752765325727, 32'sd0.018937442145368754, 32'sd-0.019821507808873512, 32'sd-0.04896347180993664, 32'sd-0.09898844482664602, 32'sd-0.06519578043292246, 32'sd-0.251751903016299, 32'sd-0.2954989726879383, 32'sd-0.17655731568350436, 32'sd-0.07953527389968294, 32'sd0.10750190122791753, 32'sd0.07164205018030105, 32'sd-0.0907129804962335, 32'sd-0.05419365424245946, 32'sd-0.05595288991959553, 32'sd-0.1303469548364578, 32'sd0.032483052443791634, 32'sd-0.07701117829779602, 32'sd-0.015122708665514894, 32'sd-0.0663376147310489, 32'sd-0.020711843074783392, 32'sd0.0291379404336848, 32'sd0.054172902653007796, 32'sd-0.10164367035979072, 32'sd0.012264515493233081, 32'sd-0.14871114559752383, 32'sd-0.05325336928921896, 32'sd-0.04375266308608985, 32'sd-0.09601592133690895, 32'sd-0.057847911253936915, 32'sd0.014353957588851107, 32'sd0.022099582150890393, 32'sd-0.02239271348599609, 32'sd-0.1044981578905944, 32'sd-0.13173058556976353, 32'sd-0.2467159368723631, 32'sd-0.1833631685054037, 32'sd0.03221005255271337, 32'sd0.10403259473973678, 32'sd-0.023443696836123063, 32'sd-0.037497459174879406, 32'sd-0.009753566098723259, 32'sd-0.07455387341349676, 32'sd-0.15547119373432242, 32'sd-0.02563555697201052, 32'sd0.030000150605959792, 32'sd-0.05346026860429057, 32'sd0.027396340157813476, 32'sd0.1069055516085615, 32'sd0.06488028939589242, 32'sd-0.05323966417080367, 32'sd0.02301199177260504, 32'sd-0.05541909500225654, 32'sd-0.034552878003985016, 32'sd-0.03397200422898551, 32'sd-0.05029142749328376, 32'sd-0.015569211445724937, 32'sd-0.09386207169703534, 32'sd-0.05599325137407301, 32'sd-0.02884912083401597, 32'sd-0.15768135532773503, 32'sd-0.07792012945510118, 32'sd-0.17968876859202107, 32'sd-0.08448116120987109, 32'sd-0.08301076354581806, 32'sd0.026570644001700797, 32'sd0.06418727619888992, 32'sd0.0794115234155312, 32'sd-0.13352470844656808, 32'sd-0.04727826459639839, 32'sd-0.11375564100040317, 32'sd-0.0485591263458659, 32'sd-0.0954779286857958, 32'sd0.004559771114188889, 32'sd-0.012207836020927761, 32'sd0.053763801158632635, 32'sd0.1529269986950181, 32'sd0.030736545022008545, 32'sd0.044007330890736315, 32'sd-0.023526664001365757, 32'sd0.06058160130325854, 32'sd-0.10362266664556413, 32'sd0.0010917957440890478, 32'sd-0.08449426686319399, 32'sd-0.053966512212269745, 32'sd-0.06782643124169586, 32'sd0.02887334536671423, 32'sd-0.048881201302010846, 32'sd-0.06820225596165996, 32'sd-0.07225148526192521, 32'sd-0.12512189175492994, 32'sd-0.12288060096254047, 32'sd-0.06189051643679756, 32'sd-0.11685025053405627, 32'sd-0.0353578897922024, 32'sd-0.11493098279798981, 32'sd-0.11541187704640411, 32'sd-0.07736975508998738, 32'sd-0.010312135475799806, 32'sd-0.08725195287456365, 32'sd-0.07901029531205597, 32'sd-0.03554855449207593, 32'sd0.020605070439737937, 32'sd0.06986800744904845, 32'sd-0.002232766055821526, 32'sd0.053831209298330754, 32'sd0.05406001612994242, 32'sd0.03493821254743159, 32'sd-0.13046779901448832, 32'sd-0.05223577507291415, 32'sd-0.05072785331965583, 32'sd0.03413735302199179, 32'sd-0.12591537530855978, 32'sd-0.06810602720969561, 32'sd-0.022985323543062333, 32'sd0.018622540347255617, 32'sd0.043546416714134575, 32'sd0.13257356934077957, 32'sd-0.1000774205126313, 32'sd-0.20531191128611057, 32'sd-0.13942259264396817, 32'sd-0.038901055661869494, 32'sd-0.07747806102712099, 32'sd-0.04334423968340817, 32'sd-0.026389125178144703, 32'sd0.011843541830928074, 32'sd0.025891827285294423, 32'sd0.0046564198895548675, 32'sd-0.06868608706677283, 32'sd0.015140482192904956, 32'sd-0.08642607754989369, 32'sd-0.0956990821546494, 32'sd0.013212885753528822, 32'sd-4.192383356090541e-124, 32'sd-0.04234300361699652, 32'sd0.008160952202780498, 32'sd-0.06493006318060496, 32'sd0.02008663938737588, 32'sd-0.11139065452308317, 32'sd-0.07731638104870754, 32'sd-0.025268757301189246, 32'sd-0.05605224585895927, 32'sd-0.01900013876923792, 32'sd0.13719167774665356, 32'sd0.04611650956680938, 32'sd-0.03629917265413576, 32'sd-0.1632745728341349, 32'sd-0.09346157853412493, 32'sd-0.14441934587538593, 32'sd-0.07906301408779173, 32'sd-0.04048729052182599, 32'sd-0.047248165911629836, 32'sd0.0382124560695194, 32'sd-0.0856622253916548, 32'sd-0.11989214859220455, 32'sd-0.09547609171946911, 32'sd-0.0841409413803729, 32'sd-0.08633648387393211, 32'sd0.08816955658339322, 32'sd-0.007685971072606079, 32'sd0.03415012727773575, 32'sd0.0017855813365911972, 32'sd0.0012721246855385464, 32'sd-0.04941246896865366, 32'sd-0.12693540678827728, 32'sd-0.05189891428723624, 32'sd-0.0537678161785788, 32'sd0.0025177901755041366, 32'sd0.003449268812921221, 32'sd-0.02040826133797719, 32'sd0.011016516643398595, 32'sd0.11295450104675663, 32'sd0.059326059057329156, 32'sd0.1277089534042418, 32'sd0.006203211404658901, 32'sd-0.14793953506984342, 32'sd-0.12099214470274304, 32'sd-0.0940889669700356, 32'sd-0.024555723049254456, 32'sd-0.11723628930673073, 32'sd0.0021014380540428693, 32'sd-0.003957409188457061, 32'sd-0.12089748152713695, 32'sd-0.09382731719350706, 32'sd-0.07544228492856134, 32'sd-0.0013419644304736552, 32'sd-0.006381209939359237, 32'sd0.05943245315554029, 32'sd-0.008805611562220757, 32'sd0.01719141278842474, 32'sd-0.0074981411535102625, 32'sd0.07374792736237629, 32'sd-0.05814028451207002, 32'sd-0.0098863338244557, 32'sd-0.11676988514513932, 32'sd0.05200322729758571, 32'sd0.15392622067617573, 32'sd0.016763814696147586, 32'sd-0.010991736759165562, 32'sd0.019445532568728264, 32'sd0.0751491868007437, 32'sd-0.03571483005510675, 32'sd0.014933308040874201, 32'sd-0.16850024221513726, 32'sd-0.007686881044741913, 32'sd-0.005324691435641076, 32'sd-0.024782216375503978, 32'sd-0.09206503236970714, 32'sd-0.02783256835607372, 32'sd0.16232440115539964, 32'sd-0.01323269744990057, 32'sd0.0002771776205647352, 32'sd-0.09334906108166244, 32'sd-0.06342895748951494, 32'sd0.10220761941156986, 32'sd0.09158561996032358, 32'sd0.055977527646753, 32'sd6.893690048212946e-126, 32'sd-0.02601290938691207, 32'sd-0.04710699153898181, 32'sd0.072507085738783, 32'sd-0.06779248375791777, 32'sd0.05055453524159249, 32'sd0.08718805117843793, 32'sd0.04104534024473176, 32'sd0.14640078302527704, 32'sd-0.06385148204393726, 32'sd0.14056966778449237, 32'sd0.18797227255339763, 32'sd0.16844697568021297, 32'sd0.11821597994769066, 32'sd0.12437189364526897, 32'sd0.12679737116921125, 32'sd0.055924619111919406, 32'sd-0.044717216008400215, 32'sd-0.009433685962183701, 32'sd-0.021541168507070576, 32'sd0.12883562880032232, 32'sd0.06425983383587715, 32'sd-0.07110669962116058, 32'sd0.025675667206886677, 32'sd-0.03840741695329596, 32'sd-0.039489112006710465, 32'sd-0.05382050346386405, 32'sd-0.02494146852206704, 32'sd0.007922505337565482, 32'sd-0.0899661079095102, 32'sd-0.0497436475614546, 32'sd-0.025849768356861275, 32'sd-0.06999542776147478, 32'sd0.07983191833322091, 32'sd0.003796942397567409, 32'sd-0.04539158032163903, 32'sd0.06925214677967274, 32'sd0.05672149363151623, 32'sd0.05167988032912503, 32'sd0.15801031246397032, 32'sd0.1351736936559389, 32'sd0.09535758019307297, 32'sd0.16095753231449406, 32'sd0.20288757697532459, 32'sd0.07314757421771129, 32'sd0.02772999109832738, 32'sd0.05806996294233741, 32'sd0.027482806989218535, 32'sd0.021517987871328224, 32'sd-0.004107243847620566, 32'sd-0.06299595120892242, 32'sd0.07494212602759048, 32'sd-0.11286396716057509, 32'sd-0.026014310459780067, 32'sd0.028895610704728184, 32'sd0.031168651532199197, 32'sd0.019036761822761154, 32'sd-0.014515012067724107, 32'sd0.03824396839268055, 32'sd0.01993200742502811, 32'sd-0.04537484305709162, 32'sd0.0839265016850264, 32'sd-0.014870871170324967, 32'sd0.015558039015592958, 32'sd0.015531989920193858, 32'sd0.05652733353866809, 32'sd-0.046070157322364656, 32'sd0.05800281102730785, 32'sd-0.020048040482276888, 32'sd0.08741104550587192, 32'sd0.14726984312934374, 32'sd0.07827917038392466, 32'sd0.06683062453116433, 32'sd0.0822421634700082, 32'sd0.08741188884038778, 32'sd-0.006660429732524272, 32'sd-0.044742310155296415, 32'sd-0.024875690958339195, 32'sd0.08203090708592299, 32'sd0.08030347543486402, 32'sd0.04049753255420578, 32'sd0.004353392970635165, 32'sd-0.07125145922974284, 32'sd0.04120276695062269, 32'sd-1.75880873257844e-117, 32'sd0.022066015705314673, 32'sd-0.0491944718373099, 32'sd-0.08886574477981703, 32'sd0.008028030653927347, 32'sd0.006173437950996164, 32'sd-0.03526138814848193, 32'sd0.035408785230982606, 32'sd0.0639223692128965, 32'sd0.10265243465395098, 32'sd-0.04175834230169298, 32'sd0.047454203376116534, 32'sd0.030593667193074298, 32'sd-0.026667854882639355, 32'sd0.12415615093705086, 32'sd0.04695788350417374, 32'sd0.009031753302998638, 32'sd-0.017770192900271792, 32'sd-0.007844458112037125, 32'sd-0.00450204303913157, 32'sd-0.038554649659228696, 32'sd-0.11099462844130756, 32'sd0.09079649353228186, 32'sd0.09780214296695905, 32'sd0.0699798002695545, 32'sd0.1020314108494461, 32'sd-0.15132817855716277, 32'sd-2.8755353645741343e-124, 32'sd9.454256082108085e-123, 32'sd-1.186432246722735e-121, 32'sd0.012341434742857704, 32'sd0.02225831009733327, 32'sd0.04271621041294458, 32'sd-0.0561701699505041, 32'sd-0.09212424072800814, 32'sd-0.0405200123951211, 32'sd0.02483942479443649, 32'sd-0.00721994612461249, 32'sd-0.011423468124745035, 32'sd0.023316319505008908, 32'sd-0.02002772978959948, 32'sd-0.06098423212156371, 32'sd0.06292346183223886, 32'sd-0.024525256431111447, 32'sd-0.08930793184213318, 32'sd0.015541255362249087, 32'sd0.06883436768554863, 32'sd0.08797537764116213, 32'sd-0.031975406641678014, 32'sd-0.03306538685353049, 32'sd0.012367211160463524, 32'sd-0.01495947133530379, 32'sd-0.01601288314477707, 32'sd-0.010827482285286518, 32'sd0.039000853728658774, 32'sd-1.856925913106287e-116, 32'sd-1.8410357320080665e-124, 32'sd3.256635465995761e-123, 32'sd0.040583503996053136, 32'sd0.044398217063767245, 32'sd0.11484504877629875, 32'sd-0.009376911679644093, 32'sd0.09280713349780247, 32'sd0.05382938593929052, 32'sd0.11248563997185648, 32'sd0.048593545880478664, 32'sd0.14239738360265788, 32'sd0.01471007370283632, 32'sd0.06688250248105931, 32'sd0.013143304593651371, 32'sd0.0317408827128506, 32'sd-0.003021072801916912, 32'sd-0.025265562981385777, 32'sd0.03432215706502356, 32'sd0.1279608502941492, 32'sd0.03646381047610832, 32'sd0.08067241690263936, 32'sd0.10277741467668486, 32'sd0.07974953106926917, 32'sd0.008329290494233308, 32'sd0.020001250037535705, 32'sd0.025621138578744526, 32'sd0.05573160962859252, 32'sd9.799981315382298e-117, 32'sd2.6262065652310683e-121, 32'sd1.1919985560137306e-118, 32'sd-8.666728698982349e-125, 32'sd0.06165478939785956, 32'sd0.013267072798064761, 32'sd-0.059060400824449945, 32'sd0.059523092258043746, 32'sd-0.0042531233549472705, 32'sd0.0798398932621041, 32'sd-0.030720458453330966, 32'sd-0.1082285584218032, 32'sd-0.11367849634896306, 32'sd0.03153668153674727, 32'sd-0.00228764935889068, 32'sd0.03767742143128723, 32'sd-0.021008247987313468, 32'sd0.03786147309151438, 32'sd0.058082579265879127, 32'sd0.048036453396028155, 32'sd-0.0448178710614027, 32'sd-0.09130596279747409, 32'sd-0.12282965884777299, 32'sd0.036945383823725954, 32'sd-0.0746319568861678, 32'sd0.002067842504986628, 32'sd0.0017472416073253342, 32'sd-2.5837710384768392e-114, 32'sd-1.2577703063534593e-127, 32'sd1.343188847849663e-118, 32'sd2.444781151843264e-125, 32'sd1.327487600019706e-127, 32'sd1.298473364923974e-122, 32'sd0.04582824339388617, 32'sd0.03714662417744397, 32'sd0.011605786593643815, 32'sd0.0463970959229609, 32'sd-0.029434715021637716, 32'sd0.06995754598513024, 32'sd0.0304975237757438, 32'sd0.08782497959158592, 32'sd0.049247961352045164, 32'sd0.07214153179915248, 32'sd0.11384525029183906, 32'sd0.02299708571631324, 32'sd0.08401209678853323, 32'sd-0.01928202660643926, 32'sd-0.03437938973270604, 32'sd0.052253629324054134, 32'sd0.005043245726012367, 32'sd-0.07982689168619192, 32'sd-0.03709871671191033, 32'sd0.04396752753397737, 32'sd1.385797183497224e-119, 32'sd7.717058787322122e-117, 32'sd1.011018183073033e-124, 32'sd-1.7669379691441002e-123},
        '{32'sd-4.793499259065451e-123, 32'sd1.7817851241907142e-123, 32'sd3.8045895631331606e-119, 32'sd-1.7523678124010233e-127, 32'sd-7.107017596273172e-115, 32'sd-4.175290833688581e-125, 32'sd2.877549900241929e-124, 32'sd-2.0619181042352864e-120, 32'sd3.1045372373897795e-120, 32'sd8.661654598869252e-120, 32'sd1.6962587420368327e-124, 32'sd-4.652280710680983e-118, 32'sd0.022272524007886377, 32'sd0.023143942785065298, 32'sd-0.010213772308689353, 32'sd-0.043137974779601095, 32'sd-3.259977651930767e-120, 32'sd2.8627833064227808e-126, 32'sd2.994127376374434e-122, 32'sd1.6325006829976367e-115, 32'sd2.38868336715659e-125, 32'sd-1.0093126770571849e-119, 32'sd-3.6264979227868416e-129, 32'sd-1.2159684472439975e-126, 32'sd3.668730595767696e-118, 32'sd2.748171820428347e-120, 32'sd9.055343941293622e-120, 32'sd4.474449874837384e-127, 32'sd-8.579180644639844e-118, 32'sd-9.786229665326292e-123, 32'sd-2.4028142506891993e-119, 32'sd4.246857836534226e-125, 32'sd0.09100339700747585, 32'sd0.10332219497642943, 32'sd0.02198358134600085, 32'sd-0.010022290817804713, 32'sd0.04189911427243061, 32'sd0.06532234091689805, 32'sd-0.06647009947441433, 32'sd-0.007145393385583712, 32'sd-0.027929607144625664, 32'sd0.032745075510115546, 32'sd-0.08439919551061392, 32'sd-0.05211431418744306, 32'sd0.08111456328923652, 32'sd-0.007877767158165145, 32'sd0.01940629713141744, 32'sd0.08949125802972002, 32'sd0.02566411968474057, 32'sd0.08615315751264441, 32'sd0.0636628343052672, 32'sd0.023020661982865773, 32'sd3.841872643988583e-120, 32'sd2.8750007265334687e-121, 32'sd-2.2558628424679505e-124, 32'sd-1.6822935091725549e-125, 32'sd-3.3312179360322126e-120, 32'sd4.874253033314461e-123, 32'sd0.0885831819789811, 32'sd0.06482278411709658, 32'sd0.07319794022893082, 32'sd0.10890156897155703, 32'sd0.0004765900427699302, 32'sd0.0023834582793966527, 32'sd-0.06431689163936964, 32'sd0.026308608699120193, 32'sd-0.0021659738425115933, 32'sd-0.0782691084754845, 32'sd0.06485693729411973, 32'sd0.026139602717001456, 32'sd-0.08473578153938673, 32'sd-0.0769070909784514, 32'sd-0.011740983919554734, 32'sd-0.08824445246946805, 32'sd0.0729703848580459, 32'sd-0.014120543929567408, 32'sd0.10614383253389433, 32'sd0.05541146881289805, 32'sd0.03474574577195961, 32'sd0.0575470257041089, 32'sd-0.029252653304101806, 32'sd0.08871252723083556, 32'sd-3.9644807471323695e-122, 32'sd-2.717534741325302e-118, 32'sd-2.5160473606226436e-130, 32'sd-1.04733370243519e-120, 32'sd0.01586266694684782, 32'sd0.015618628079495666, 32'sd0.034538102609922544, 32'sd-0.0849401633629166, 32'sd0.008293422815982995, 32'sd0.02208959701909569, 32'sd0.032376320982823406, 32'sd-0.039544711370446156, 32'sd-0.15591265937890747, 32'sd0.028603528260788602, 32'sd0.035653842209660655, 32'sd0.007411818350074638, 32'sd-0.05258746778418529, 32'sd-0.09937844208871295, 32'sd-0.040189679260908474, 32'sd-0.025893028922360707, 32'sd0.0828839872908801, 32'sd-0.01363143068852608, 32'sd-0.03476626891494513, 32'sd-0.08530943942814198, 32'sd-0.022081897369928688, 32'sd-0.10898659996931, 32'sd-0.0002097298441627111, 32'sd-0.057555131346490665, 32'sd0.03637977460317933, 32'sd-3.7363443528278696e-125, 32'sd-3.8176897512129294e-126, 32'sd0.032205605303053275, 32'sd-0.0013701124744585514, 32'sd0.08137758624658409, 32'sd-0.004841288853713028, 32'sd0.017450893495523916, 32'sd0.012693444793359227, 32'sd0.06062547207083541, 32'sd-0.12508887704980576, 32'sd0.002741121410155196, 32'sd-0.087451590369288, 32'sd-0.040846056157482886, 32'sd-0.03554030377621925, 32'sd-0.06903035919472598, 32'sd-0.08044361719398947, 32'sd-0.10210390651478642, 32'sd-0.1161283220423743, 32'sd-0.10679013325962639, 32'sd0.048157790700228624, 32'sd-0.0727018536721353, 32'sd-0.13572286671636802, 32'sd-0.1054195328828396, 32'sd-0.0737211590793884, 32'sd-0.11396714918620829, 32'sd-0.0555122635628963, 32'sd-0.1396304100868482, 32'sd0.047976100034264, 32'sd0.06618340122161126, 32'sd-1.0968613571440987e-117, 32'sd0.0008742986071108623, 32'sd0.029111446243990546, 32'sd-0.05542027649672575, 32'sd-0.027147100652055965, 32'sd0.05352242014306704, 32'sd-0.024405805559406142, 32'sd0.04067397122810817, 32'sd-0.02417686136110164, 32'sd0.011748028455624861, 32'sd-0.0705811194562619, 32'sd-0.08433167684639498, 32'sd-0.1484506580928558, 32'sd-0.18732938657864096, 32'sd-0.24041560976040263, 32'sd-0.24160360047649995, 32'sd-0.23203251172488734, 32'sd-0.19589174021879643, 32'sd-0.0356202304166319, 32'sd0.10405032488133656, 32'sd0.16577617672999212, 32'sd-0.11268724470296317, 32'sd-0.07918980502635381, 32'sd-0.10104946297559346, 32'sd-0.105600903492147, 32'sd-0.01043721788008349, 32'sd0.10461974894430104, 32'sd0.02139151261297617, 32'sd4.734911204882914e-117, 32'sd0.06873123027118977, 32'sd-0.026771443240290953, 32'sd-0.07572020478558728, 32'sd-0.006477581910073623, 32'sd-0.0603215276731235, 32'sd-0.18645901254785308, 32'sd-0.04714663193999112, 32'sd-0.11356980619023553, 32'sd-0.07798925352056331, 32'sd0.005957191798366989, 32'sd-0.028658986715439667, 32'sd-0.20080820469228677, 32'sd-0.25596585430262003, 32'sd-0.2054500645816341, 32'sd-0.1572338805735524, 32'sd-0.24134230594501196, 32'sd-0.035917626087768696, 32'sd0.08283690086945347, 32'sd0.17254522012473308, 32'sd0.11706914276721962, 32'sd0.008547149206290785, 32'sd-0.004423033432010747, 32'sd0.034101962082155726, 32'sd0.060479706454724315, 32'sd0.0610848421457267, 32'sd0.07639656096540524, 32'sd-0.10903728437924098, 32'sd0.03998376188852352, 32'sd-0.032062012071035345, 32'sd-0.03357529413166268, 32'sd0.017358559459419227, 32'sd-0.01633733595213928, 32'sd0.00653852388652139, 32'sd-0.10408548671616577, 32'sd-0.14123543489342946, 32'sd-0.01869734307030415, 32'sd-0.03017069604160516, 32'sd0.02902644511469202, 32'sd-0.09124863509987044, 32'sd-0.055596768682003105, 32'sd0.03175979166279431, 32'sd-0.005749421341255418, 32'sd0.1392518668625025, 32'sd0.03572065165606963, 32'sd0.14240678179934416, 32'sd0.07548506342373155, 32'sd0.176224992899952, 32'sd0.19351264926119463, 32'sd0.15518553008325808, 32'sd-0.0492436549752466, 32'sd0.07635295369262991, 32'sd0.00813230262656249, 32'sd-0.05300638088352224, 32'sd0.12810931575192788, 32'sd0.04279800011664585, 32'sd0.008834943690651855, 32'sd0.04359457668352895, 32'sd-0.007419673684313446, 32'sd-0.07557309508963095, 32'sd-0.1399994991760412, 32'sd-0.12338294742207519, 32'sd0.014238371590294584, 32'sd-0.13737974467763564, 32'sd-0.14462048809116473, 32'sd-0.02011139237336105, 32'sd-0.012916597669750477, 32'sd0.0542403576436268, 32'sd0.09523194333897055, 32'sd0.14884874572583134, 32'sd0.2212334925571347, 32'sd0.17248294480562593, 32'sd0.23036649166010922, 32'sd0.12728098096272514, 32'sd0.18385408569143308, 32'sd0.17477908568933087, 32'sd0.16938833831577016, 32'sd0.11657109073804237, 32'sd0.10048337214084074, 32'sd-0.014071020970651322, 32'sd0.026092711645590447, 32'sd-0.0033762516308020597, 32'sd-0.003510817949161476, 32'sd-0.053173053903269464, 32'sd0.007261054979109062, 32'sd-0.06371302588608456, 32'sd-0.06387387605913648, 32'sd0.003941931897419328, 32'sd-0.020879022410522342, 32'sd-0.06595064865457714, 32'sd-0.07403519222618267, 32'sd-0.03595028652360169, 32'sd-0.07450937044280792, 32'sd-0.08484907425152972, 32'sd0.05312508566548204, 32'sd0.09289853039822919, 32'sd0.20016401942511425, 32'sd0.27989346196511455, 32'sd0.1831916043322045, 32'sd0.12977528132952007, 32'sd0.16775179634292509, 32'sd0.038418173028564456, 32'sd0.19530867725726966, 32'sd0.24624123015029312, 32'sd0.0005693735631476593, 32'sd0.018108360588345477, 32'sd0.07604717407592697, 32'sd-0.047904199474131784, 32'sd0.12699576942479157, 32'sd0.03988274571140344, 32'sd-0.009210335534622676, 32'sd0.049924770990866674, 32'sd0.07766810192364475, 32'sd-0.03387457534774433, 32'sd-0.012283827646908104, 32'sd-0.028099354250202397, 32'sd-0.03294314517365172, 32'sd0.011245065696629536, 32'sd0.0505543476554223, 32'sd-0.0578909344414955, 32'sd-0.07005589603042589, 32'sd0.06000300370514291, 32'sd0.24152203240447803, 32'sd0.055630038875317527, 32'sd0.14029640107437785, 32'sd0.17611361671365902, 32'sd0.007860783507107389, 32'sd0.13859389504458278, 32'sd0.05926924577078475, 32'sd-0.02927850724386927, 32'sd0.007899932933391144, 32'sd-0.01166931092065662, 32'sd-0.07759937069711069, 32'sd-0.03465297281175916, 32'sd-0.0238938332382102, 32'sd-0.13857708050655776, 32'sd0.056561184187062366, 32'sd0.0930286272627042, 32'sd0.07569826522692616, 32'sd0.01608290283530089, 32'sd-0.020737965200894545, 32'sd0.005978210628160927, 32'sd-0.015172234744865225, 32'sd-0.13258436705655668, 32'sd0.11878310162904372, 32'sd0.08126614830519242, 32'sd-0.01173990045631789, 32'sd-0.06551521975088855, 32'sd-0.07115151514311088, 32'sd0.12751534117967167, 32'sd-0.05523887349084103, 32'sd0.1155540034477712, 32'sd0.07981695336458007, 32'sd0.09721245361029494, 32'sd0.011642877147611747, 32'sd0.06678800281772553, 32'sd-0.05384593017682763, 32'sd-0.1082351332011997, 32'sd-0.05906355562447039, 32'sd-0.13347289523667652, 32'sd-0.10733906490310688, 32'sd-0.19077132022820084, 32'sd-0.07297082178203443, 32'sd-0.0987842435019752, 32'sd-0.08841207873192418, 32'sd0.037007738169945764, 32'sd0.005820540817033481, 32'sd0.12056774441905348, 32'sd0.013903537459775737, 32'sd0.010845372961810382, 32'sd0.01878831056641224, 32'sd0.029174582143170532, 32'sd0.033329588667144895, 32'sd0.063577128380327, 32'sd-0.032268220140684145, 32'sd-0.09381710975550517, 32'sd0.036847860767181446, 32'sd0.019270247399255525, 32'sd-0.052444933848449095, 32'sd-0.045772994275614064, 32'sd-0.027641868031100896, 32'sd0.0658602401628911, 32'sd-0.014791168731536361, 32'sd-0.03548104299150111, 32'sd-0.0823298722904528, 32'sd-0.16229324002233528, 32'sd0.04733314178574783, 32'sd-0.08678098717939296, 32'sd-0.05213508421232943, 32'sd-0.0369354632453668, 32'sd-0.03991661378660415, 32'sd-0.032981199837427526, 32'sd-0.011204575051429707, 32'sd-0.1406995152665423, 32'sd-0.014812209651185647, 32'sd-0.06111322873972515, 32'sd0.02495951888940355, 32'sd0.012829851813120508, 32'sd0.013638031798818485, 32'sd0.042938621644720155, 32'sd0.005520561035082236, 32'sd-0.04293353659246869, 32'sd-0.03392893066325124, 32'sd-0.059418652660849, 32'sd-0.028797793489877186, 32'sd-0.1554661941869421, 32'sd-0.0558757177783043, 32'sd-0.02508094298750629, 32'sd-0.0652863002673582, 32'sd0.061661306219240396, 32'sd-0.03893837526615953, 32'sd0.001561186952805569, 32'sd-0.16071782255267755, 32'sd-0.16788404747244423, 32'sd-0.08441906194788473, 32'sd-0.0006882575216848, 32'sd-0.06883995278624448, 32'sd-0.11435451878252503, 32'sd-0.054958936175439815, 32'sd-0.07620927109655166, 32'sd-0.13211295289652228, 32'sd-0.1900941908467865, 32'sd-0.034614060334895724, 32'sd0.017914096501371737, 32'sd0.06701176028563335, 32'sd0.0029207859659597154, 32'sd0.043697102185575584, 32'sd-0.045676598547395024, 32'sd0.1448692945246807, 32'sd-0.07526559585171726, 32'sd0.05170088679997658, 32'sd-0.01849131991203076, 32'sd-0.06760612953604517, 32'sd0.012546451229969004, 32'sd-0.0894829944398961, 32'sd-0.012486012142285762, 32'sd-0.0337850406350452, 32'sd0.038870849393279144, 32'sd0.05768891630016023, 32'sd0.06148055293124081, 32'sd-0.0003094835192113443, 32'sd-0.13942514237541856, 32'sd0.009051430852619766, 32'sd-0.1854045243310062, 32'sd0.06464287924040418, 32'sd-0.08008450774313598, 32'sd-0.0811930460507051, 32'sd-0.030310312352590022, 32'sd0.12779035382320317, 32'sd-0.025082791663584857, 32'sd-0.06963260966812782, 32'sd-0.00022223444537955507, 32'sd0.05803430113836818, 32'sd-0.004934839048267891, 32'sd-0.08160383835862524, 32'sd0.00022749303595336133, 32'sd0.2021546744754711, 32'sd0.19364878698896426, 32'sd0.03843810792411728, 32'sd-0.05200613164193777, 32'sd-0.04293487274891968, 32'sd-0.07207328118033608, 32'sd0.09207158933649734, 32'sd-0.01822661574247617, 32'sd0.11446757723030815, 32'sd0.03173874132878525, 32'sd0.04463856952608443, 32'sd-0.12134872184146171, 32'sd-0.0876913192239938, 32'sd-0.033499091744992555, 32'sd-0.07447791495554625, 32'sd-0.028130995948955257, 32'sd0.019425722357596827, 32'sd0.052194900703406426, 32'sd-0.050004886600396, 32'sd-0.06314579946390549, 32'sd-0.010934675951763702, 32'sd0.05762536130653367, 32'sd0.0925001258861553, 32'sd0.025671689608327525, 32'sd0.007994203634531093, 32'sd0.030381281347660657, 32'sd-0.013066508737215177, 32'sd0.0003489647367228179, 32'sd0.0027687717724909204, 32'sd0.07103413498901182, 32'sd0.08301244900635678, 32'sd0.04200127207847072, 32'sd0.05848563966520648, 32'sd-0.07509261140352358, 32'sd-0.0793717313501973, 32'sd0.01159512859471804, 32'sd0.03517749777574776, 32'sd-0.030154087896998284, 32'sd-0.12012386078667464, 32'sd-0.13498285944475158, 32'sd-0.08105092959275063, 32'sd-0.013001763517002154, 32'sd-0.05848329886594281, 32'sd-0.039199996182713207, 32'sd-0.07576249371199051, 32'sd-0.011807329794687332, 32'sd0.013578111489861905, 32'sd-0.06291688815230861, 32'sd-0.01908948134019761, 32'sd0.08956990044025834, 32'sd0.027907206232809886, 32'sd0.031893068046368496, 32'sd2.728402479084134e-116, 32'sd0.023231949932184144, 32'sd-0.04444218351264332, 32'sd0.10496873151397695, 32'sd-0.1160403505863221, 32'sd0.09981602549657263, 32'sd0.19226653992334378, 32'sd0.10399912110380588, 32'sd0.07150202619966788, 32'sd0.08100830354745209, 32'sd0.06976669848081651, 32'sd-0.027555934458934537, 32'sd-0.07682377134372816, 32'sd-0.07530924676092157, 32'sd-0.023956325762718663, 32'sd0.012074151823853295, 32'sd-0.14203308229550815, 32'sd-0.11702552563948192, 32'sd0.047403518567619006, 32'sd2.952976802484423e-05, 32'sd-0.010200023444062973, 32'sd-0.05261746768394823, 32'sd0.023424759028613112, 32'sd0.0017750504718628706, 32'sd-0.17022670687680652, 32'sd-0.061562419320834984, 32'sd-0.01026673713985159, 32'sd0.006858778016132888, 32'sd0.030845250698555836, 32'sd0.04633442240913198, 32'sd-0.039142516245669515, 32'sd0.0665132763875265, 32'sd-0.02742482117409372, 32'sd0.04933877359947496, 32'sd0.07614366173522562, 32'sd0.18171008654604306, 32'sd0.10718281784223593, 32'sd-0.007138458821520725, 32'sd-0.0382438343425838, 32'sd0.02334633259476731, 32'sd0.0394308669921858, 32'sd-0.08405940831065695, 32'sd0.10407633630581405, 32'sd-0.01399899142086869, 32'sd0.044962465322891325, 32'sd0.012188792894843094, 32'sd-0.09910323739650356, 32'sd0.04026947556449388, 32'sd0.03804849477027475, 32'sd-0.11845834281475895, 32'sd-0.06417835241077188, 32'sd0.051215252584192204, 32'sd-0.04002481312994027, 32'sd-0.019748328656130174, 32'sd0.10061462726839966, 32'sd-0.07470512377734087, 32'sd0.02203813975682383, 32'sd-0.00903625543929317, 32'sd-0.09649364894304335, 32'sd0.011830673520782448, 32'sd0.049491347085446113, 32'sd-0.02161757107937246, 32'sd0.07257270631511034, 32'sd0.08155745851448455, 32'sd0.016152458787323614, 32'sd-0.008044755992266226, 32'sd0.03948765110131742, 32'sd-0.05270130484256702, 32'sd-0.012845709842132515, 32'sd-0.136266107239329, 32'sd0.07830748679081345, 32'sd-0.011900853588363226, 32'sd-0.055694915430815985, 32'sd-0.008303969663609884, 32'sd0.03247807040648958, 32'sd0.12469188202645314, 32'sd0.0398001762605715, 32'sd-0.055658674886860944, 32'sd0.05662608217540551, 32'sd0.181347169519419, 32'sd-0.0996312482126098, 32'sd0.02686832569429161, 32'sd0.10069151495080281, 32'sd-0.05800299169213112, 32'sd1.4460420364999323e-115, 32'sd0.01602857522725158, 32'sd0.025758180301946834, 32'sd0.016453821249580163, 32'sd0.0036479055053174197, 32'sd0.1509745547947051, 32'sd0.03618062186594855, 32'sd0.022991279373470924, 32'sd-0.06923791671034422, 32'sd-0.07108287483811541, 32'sd-0.05560950030062223, 32'sd-0.11042266878492518, 32'sd-0.15359154109209314, 32'sd-0.10748286868221095, 32'sd-0.01420413574554573, 32'sd0.0199947360898339, 32'sd0.020025614064095792, 32'sd0.10369725641118048, 32'sd0.02051387532679761, 32'sd0.06618997011741067, 32'sd0.09870905949105258, 32'sd-0.06261004756809482, 32'sd0.01129000063929495, 32'sd0.10319389416856191, 32'sd-0.10832547223867213, 32'sd0.08896122213777935, 32'sd0.0891861993168463, 32'sd0.05047649919608674, 32'sd0.03113006097014289, 32'sd-0.05417837967381112, 32'sd-0.12220585673309749, 32'sd0.03184619132423062, 32'sd-0.04079118526071326, 32'sd0.01820525596612254, 32'sd0.011218716949357537, 32'sd-0.12042213212615219, 32'sd-0.1244257611333567, 32'sd-0.07397048977398449, 32'sd-0.15288240723125213, 32'sd-0.027087380112772296, 32'sd-0.04769419280752349, 32'sd-0.025946925673848313, 32'sd0.026633512663631963, 32'sd-0.011792771757149588, 32'sd0.07590383351295238, 32'sd0.04015385682393842, 32'sd-0.011009436954458704, 32'sd0.11257667823683237, 32'sd0.06900501961668559, 32'sd0.04502054817711838, 32'sd-0.031141647118419245, 32'sd0.0047377160702068415, 32'sd0.05341508827783035, 32'sd0.05182418145759246, 32'sd-0.014187698342544155, 32'sd0.01486360020619684, 32'sd-0.02946350766856984, 32'sd-0.07472715910020633, 32'sd0.06996283702830734, 32'sd-0.006936934171196554, 32'sd0.03490837082717029, 32'sd-0.062399555856027855, 32'sd-0.09996898053711123, 32'sd-0.05479047610659301, 32'sd-0.06106810431918946, 32'sd0.057086227527522924, 32'sd0.04691554647355217, 32'sd-0.036174812952956714, 32'sd0.008946687300795364, 32'sd0.05215331454104541, 32'sd0.07141162304704275, 32'sd0.08038921717607207, 32'sd-0.023219603758281082, 32'sd0.15338475513490335, 32'sd0.07015967996317787, 32'sd-0.0020517642601316746, 32'sd0.1454589604316528, 32'sd0.09641396406500415, 32'sd-0.09163729387387119, 32'sd0.009396773960750206, 32'sd0.03322896669196364, 32'sd0.08144186687315998, 32'sd-0.05999782143269565, 32'sd-0.01672364346220552, 32'sd6.0953047701049716e-120, 32'sd0.025859645069770867, 32'sd0.02213474439724474, 32'sd0.03756526887400529, 32'sd-0.009611437443622986, 32'sd0.0417327287306676, 32'sd-0.027947733697720856, 32'sd0.05211519824027466, 32'sd-0.06360167600981202, 32'sd-0.04124779202545609, 32'sd-0.025910278321417863, 32'sd0.1657754492093696, 32'sd0.10792751235124821, 32'sd0.0219989301454848, 32'sd-0.00987975049715303, 32'sd-0.015067921771203146, 32'sd-0.030437096029132134, 32'sd0.08422969552348675, 32'sd-0.052204814079794895, 32'sd0.03309875170252998, 32'sd0.14767384209779388, 32'sd0.02151547501738871, 32'sd-0.03271145698240925, 32'sd-0.03673163461607611, 32'sd-0.07955110505097292, 32'sd-0.03347093517937728, 32'sd-0.006093366019148513, 32'sd3.606239658538682e-114, 32'sd7.255167094228249e-121, 32'sd1.664020690577963e-116, 32'sd0.013245991238566594, 32'sd-0.0593721575886466, 32'sd-0.008686253764440537, 32'sd-0.03182550934956571, 32'sd-0.011203193854285724, 32'sd-0.019820122552987745, 32'sd0.03543795918854373, 32'sd0.009356079055276707, 32'sd0.07407245035299685, 32'sd0.05218172402553369, 32'sd0.16080931869829193, 32'sd0.024754895625046316, 32'sd-0.001385977090719054, 32'sd0.05280615891139124, 32'sd0.003241482676317336, 32'sd0.06419020127185508, 32'sd-0.00957021883477293, 32'sd0.05031464277264339, 32'sd-0.1280582723528466, 32'sd-0.09548691150736711, 32'sd-0.0426085056470341, 32'sd-0.027638287074306506, 32'sd-0.048603747825875884, 32'sd0.001635746608955883, 32'sd0.051471341397543, 32'sd9.848917435089896e-126, 32'sd9.800467360702545e-117, 32'sd-5.727547114980149e-123, 32'sd0.004010700332439143, 32'sd-0.025382860296860692, 32'sd-0.09743829070234875, 32'sd-0.07871605977822793, 32'sd0.12971821102751646, 32'sd0.03136691001634402, 32'sd0.033330349031984105, 32'sd-0.02436313190137236, 32'sd0.024005744698858, 32'sd0.1002495138470066, 32'sd0.10068001399050712, 32'sd0.007241628018816604, 32'sd-0.07333367274301023, 32'sd0.04301102705551453, 32'sd0.08911415740873765, 32'sd0.10033697727774381, 32'sd-0.10252058911386157, 32'sd0.002358612618946273, 32'sd0.0013816566521575701, 32'sd0.04849234254507806, 32'sd-0.0034504549896320668, 32'sd-0.03245867548944135, 32'sd-0.08396823968542133, 32'sd0.004231840975315308, 32'sd-0.057205276757823366, 32'sd1.3959490039169888e-127, 32'sd-8.812057563127323e-125, 32'sd5.700060345231977e-123, 32'sd-3.4690130981797965e-116, 32'sd0.08717910433673678, 32'sd-0.11829588587188854, 32'sd0.013295425796608296, 32'sd0.08290931352971882, 32'sd0.0063983882876759825, 32'sd0.17568344705331862, 32'sd0.027208627569769526, 32'sd0.0005649045082652028, 32'sd0.07826528383221465, 32'sd0.07630422013186032, 32'sd0.12319569466748123, 32'sd0.043044661042671746, 32'sd0.21305202958114222, 32'sd0.017213495637253037, 32'sd0.07457025544307577, 32'sd0.08881240821017206, 32'sd0.08620935847384827, 32'sd0.028097501944095004, 32'sd-0.06992256231205549, 32'sd-0.1077424535004501, 32'sd-0.008182977137086307, 32'sd0.07588380707016165, 32'sd0.04491692705724429, 32'sd-4.187162402574463e-122, 32'sd-1.4905480617431254e-127, 32'sd6.0346211423226426e-120, 32'sd-1.7925905829758595e-118, 32'sd1.66729830243286e-124, 32'sd2.3354550385918979e-119, 32'sd0.09526541492954232, 32'sd0.006391077225831558, 32'sd0.0621423653675027, 32'sd0.08441272833075192, 32'sd0.11114079670616359, 32'sd0.056006344935978496, 32'sd0.13419739616718732, 32'sd0.023774367925965774, 32'sd0.04012072217218672, 32'sd0.08583198402799298, 32'sd0.01804517983929397, 32'sd0.06597832537432616, 32'sd0.0961917807016357, 32'sd0.014371100337503452, 32'sd-0.06877451386445463, 32'sd0.007723741463050341, 32'sd0.05438982336168008, 32'sd0.04529801838268916, 32'sd0.06912774064438727, 32'sd0.06608812195262835, 32'sd-5.192907781482702e-118, 32'sd8.88233949236996e-127, 32'sd-1.4383183677171495e-125, 32'sd-1.3478816409004365e-128},
        '{32'sd2.9533738175535224e-118, 32'sd-3.8566306990495066e-122, 32'sd-7.674361951270156e-127, 32'sd-6.121170527521603e-127, 32'sd-6.439788848191075e-128, 32'sd2.539779586501511e-123, 32'sd-1.3892463160581542e-118, 32'sd-8.835218142375711e-122, 32'sd-2.5759143224367645e-120, 32'sd1.285989334465638e-124, 32'sd5.026900060812104e-117, 32'sd1.8803618380245911e-121, 32'sd-0.07794241910739698, 32'sd-0.03015081182062807, 32'sd-0.005357363683594889, 32'sd-0.0015384978843547758, 32'sd1.0916321997922024e-123, 32'sd-2.715539234423651e-115, 32'sd-8.52652895070583e-117, 32'sd4.4248919279649235e-125, 32'sd-1.160541371277695e-122, 32'sd-4.462107233567505e-126, 32'sd-7.106479736180278e-120, 32'sd2.5692549884443056e-126, 32'sd3.393282511948431e-121, 32'sd2.436239346041197e-124, 32'sd6.967645156621258e-120, 32'sd-6.436632559687403e-124, 32'sd-5.0886321988489885e-118, 32'sd1.088288422638703e-127, 32'sd3.167244384682591e-121, 32'sd-2.868729274020956e-119, 32'sd0.008204893792301566, 32'sd-0.08036634106510356, 32'sd0.007151822692411485, 32'sd-0.01637146742634566, 32'sd-0.06279908890696122, 32'sd-0.022819553119058762, 32'sd-0.09328740699207276, 32'sd0.026700238238151434, 32'sd-0.03245530133803505, 32'sd0.03605152548495178, 32'sd-0.005719622874388484, 32'sd-0.025710859306022966, 32'sd0.0972312277711968, 32'sd0.08155606550610525, 32'sd-0.07681236239467343, 32'sd0.005244474568066567, 32'sd0.031656360520227696, 32'sd0.057628120539081014, 32'sd0.07101385193368571, 32'sd0.030979708226746883, 32'sd1.564811099668948e-114, 32'sd2.333656107166592e-117, 32'sd-6.950033615674302e-124, 32'sd-2.1725765370045153e-122, 32'sd7.193354534300797e-115, 32'sd-1.737793451344267e-125, 32'sd0.019975889328321804, 32'sd0.014925791102188482, 32'sd0.08307393777383963, 32'sd-0.006543316827115643, 32'sd0.04529373558877048, 32'sd0.046562050667646765, 32'sd-0.06054010923157889, 32'sd-0.03843276712774827, 32'sd0.04339323135381648, 32'sd-0.045585987834897056, 32'sd-0.08347942646348816, 32'sd0.1311883345492077, 32'sd0.0431613729628274, 32'sd0.050871300460724085, 32'sd0.0772812333128413, 32'sd-0.06220866388397358, 32'sd-0.003487183117343305, 32'sd0.026564399067511287, 32'sd0.0994300966777601, 32'sd0.12754586409151433, 32'sd0.03925696483292211, 32'sd-0.04793997332526285, 32'sd0.07291828894368274, 32'sd0.0067114238983339135, 32'sd-4.67939066655055e-123, 32'sd7.399776979648051e-122, 32'sd-1.2237918221398358e-124, 32'sd-1.0093809142028222e-117, 32'sd0.018558652479891767, 32'sd-0.021301242516058597, 32'sd-0.07220494440439011, 32'sd-0.0038381619983484877, 32'sd0.04133429770647603, 32'sd-0.06215013712916081, 32'sd-0.045042050168403854, 32'sd0.0886812747452297, 32'sd0.057361465747666165, 32'sd0.015664378794144583, 32'sd0.13980301903601014, 32'sd0.27970328341977313, 32'sd0.11330036497034214, 32'sd0.10937339347523721, 32'sd0.042693784169400416, 32'sd0.024649298028392445, 32'sd-0.011098256257890574, 32'sd-0.018976085108868366, 32'sd0.030490694843874722, 32'sd-0.001607463695239752, 32'sd-0.009723442490460421, 32'sd-0.029295264693469054, 32'sd0.01864407295593407, 32'sd-0.05753229879476058, 32'sd-0.020667356413703267, 32'sd-1.0688357581049005e-124, 32'sd1.5675025230486738e-124, 32'sd0.00855874047022101, 32'sd0.02291365227813399, 32'sd-0.06455145704737536, 32'sd0.060784294448302, 32'sd0.013046100586614654, 32'sd-0.030333396844567158, 32'sd-0.1439446939741144, 32'sd-0.11565279211417656, 32'sd0.01264248002781408, 32'sd0.13624322648056914, 32'sd0.05565979127468688, 32'sd0.07831874236397748, 32'sd0.07321928056753704, 32'sd0.03448116641459238, 32'sd-0.07205745615125157, 32'sd-0.016163888051483048, 32'sd0.032698217944860775, 32'sd0.031381326510684364, 32'sd0.09654750022380587, 32'sd0.059377173298337804, 32'sd-0.07245400222530696, 32'sd0.008399113770635519, 32'sd0.10041574263412986, 32'sd-0.006832175918044147, 32'sd0.029926070733143968, 32'sd0.010086383499241207, 32'sd-0.010896785035616375, 32'sd1.7754970916278474e-115, 32'sd0.015471411857716357, 32'sd-0.04957294992169235, 32'sd-0.02937372406201477, 32'sd0.01706529568973769, 32'sd-0.11667636795444565, 32'sd0.005268709897162422, 32'sd-0.05225021416819271, 32'sd0.014970926739712417, 32'sd0.09562932943977716, 32'sd0.12374754299945862, 32'sd0.04790710576709186, 32'sd0.11798947539330909, 32'sd0.09161132843395292, 32'sd0.20473468830487593, 32'sd0.01553769386182791, 32'sd0.18775089686212199, 32'sd0.11352952763460242, 32'sd0.16132375105763636, 32'sd0.0934368247168982, 32'sd-0.018534283443774467, 32'sd-0.05045776293317494, 32'sd0.01209737440515512, 32'sd-0.014430880644487597, 32'sd0.013665525254424151, 32'sd0.09580378800591849, 32'sd0.02584853897202604, 32'sd0.0017831669932662252, 32'sd1.1690366327149184e-123, 32'sd0.032082653156824625, 32'sd-0.01911697904774699, 32'sd-0.0002623553194948652, 32'sd-0.0025492473935363707, 32'sd-0.12265655037827602, 32'sd-0.11478389745493041, 32'sd0.01975327307995164, 32'sd-0.051801397472694174, 32'sd0.02503045275092342, 32'sd-0.07756514890703343, 32'sd0.10366753772008981, 32'sd0.028388324451619363, 32'sd0.10308985670999316, 32'sd0.12447280179866085, 32'sd-0.009389664707498684, 32'sd0.08295148705987672, 32'sd0.01040139904789796, 32'sd0.03572679078988156, 32'sd-0.030741126940501608, 32'sd-0.012709087379952893, 32'sd-0.11040352837548384, 32'sd0.01628715990878055, 32'sd-0.06596410738904321, 32'sd-0.09649755240989837, 32'sd-0.045875358167571295, 32'sd0.05152517854213922, 32'sd0.05130965044549123, 32'sd0.019320254808799203, 32'sd0.07676151495538103, 32'sd-0.05384077726725081, 32'sd-0.037481540442270894, 32'sd-0.023959034713367574, 32'sd-0.06537194378620265, 32'sd-0.08544319747535302, 32'sd-0.07685028277504036, 32'sd0.049709633486931484, 32'sd-0.0006728912735152621, 32'sd0.07522835975449507, 32'sd0.058121287867528286, 32'sd0.04302862928768408, 32'sd0.047064448191794665, 32'sd0.013890657545307649, 32'sd-0.011891527272766156, 32'sd-0.0579002762621367, 32'sd-0.08694306412708282, 32'sd-0.1137308433101974, 32'sd-0.07122514961402107, 32'sd-0.08639006398229168, 32'sd-0.10376099821709399, 32'sd-0.16342393021204096, 32'sd-0.09012516903229417, 32'sd-0.11791538090515696, 32'sd-0.04189739573119676, 32'sd-0.0012623197579178793, 32'sd-0.05608251558652229, 32'sd0.05225885954806033, 32'sd-0.007815211346954103, 32'sd0.04397582491258995, 32'sd-0.01668414470733484, 32'sd-0.10217607408557748, 32'sd-0.030686832072716757, 32'sd0.0217069852533767, 32'sd-0.003818115045826096, 32'sd0.11229373699281918, 32'sd0.11435286799122743, 32'sd0.09641746963455239, 32'sd0.11740211146226086, 32'sd0.08282156115473475, 32'sd0.0017018983149424307, 32'sd-0.015515090207198204, 32'sd-0.17349782803424052, 32'sd-0.15705386747617583, 32'sd-0.026934998286648776, 32'sd-0.13016937503689202, 32'sd-0.1781322738985728, 32'sd-0.07416458622177997, 32'sd-0.09441915565852131, 32'sd-0.10669356987800106, 32'sd-0.07343055848589812, 32'sd-0.08130764919741372, 32'sd-0.06974998718103173, 32'sd-0.0043827645250951045, 32'sd0.06983880612538142, 32'sd0.036081132329388046, 32'sd0.07541738727418894, 32'sd0.004206132632871969, 32'sd-0.06312395123401801, 32'sd-0.07161951179796157, 32'sd-0.020509463313204163, 32'sd0.11081029418571384, 32'sd0.12301697959245127, 32'sd0.12293017575220715, 32'sd0.07423846836221518, 32'sd0.03589390437819953, 32'sd0.054945913752661946, 32'sd-0.04096193906632886, 32'sd-0.04510148896487856, 32'sd-0.11037833456405716, 32'sd-0.08997278145026072, 32'sd-0.2477741302025897, 32'sd-0.13386792743816706, 32'sd-0.007658903134397621, 32'sd-0.08112250886073336, 32'sd-0.16431240280749326, 32'sd-0.0262824700885305, 32'sd-0.09464795426116539, 32'sd-0.10595000766210884, 32'sd0.08987764453850472, 32'sd-0.04976543367069724, 32'sd0.06427916029604752, 32'sd0.07703828970803554, 32'sd0.00859188390023449, 32'sd0.07220720765694423, 32'sd0.08597614643710183, 32'sd-0.11786633099802732, 32'sd-0.17211830766533462, 32'sd-0.018604443214245214, 32'sd-0.016679533146713357, 32'sd-0.036777989054366335, 32'sd0.0802673244036422, 32'sd0.011889985268743441, 32'sd0.00047458983514779926, 32'sd-0.00044659016822419794, 32'sd-0.08418973990017117, 32'sd-0.026010002194737248, 32'sd-0.04680865719832838, 32'sd-0.10893366595835542, 32'sd-0.15296984643435937, 32'sd-0.02344450555440832, 32'sd-0.0509830878162863, 32'sd0.0434952539580213, 32'sd0.022988338533452373, 32'sd0.022203955106076156, 32'sd0.04920589095058779, 32'sd0.058194553379900094, 32'sd0.09944703679536639, 32'sd-0.03439030677849634, 32'sd0.030083745638773477, 32'sd-0.02932305491355376, 32'sd-0.026685164900378824, 32'sd0.003394910290584911, 32'sd0.010881099792428415, 32'sd0.021626928900114764, 32'sd-0.08626143570655066, 32'sd-0.09304616840083946, 32'sd-0.04670461959458634, 32'sd-0.04335424068556237, 32'sd-0.1023230742911636, 32'sd-0.11921300586489657, 32'sd-0.07642966342570136, 32'sd-0.1383675498191478, 32'sd-0.20520668931016273, 32'sd-0.010159190849347077, 32'sd0.06584516948234345, 32'sd0.08600797405863203, 32'sd0.05249376728803677, 32'sd-0.037974252064477944, 32'sd0.09248081645582301, 32'sd0.112155363861861, 32'sd0.013079986926104998, 32'sd0.08350767324775467, 32'sd0.061744323271475124, 32'sd0.2516686252827062, 32'sd0.0956798745404152, 32'sd0.04704502406678147, 32'sd0.07421730500871349, 32'sd0.09523802966047162, 32'sd0.022654668602199408, 32'sd-0.05949942047946985, 32'sd-0.012794435148211861, 32'sd0.05955014817861784, 32'sd-0.009238024469241296, 32'sd-0.008335578631007914, 32'sd-0.06232208066035201, 32'sd-0.03262496214600414, 32'sd-0.07053553464029919, 32'sd-0.09956820135197568, 32'sd-0.08935729522784058, 32'sd-0.06486226294914257, 32'sd-0.11083138159239178, 32'sd-0.03981803734545173, 32'sd0.006928765901770189, 32'sd0.13762160194972206, 32'sd0.033008654242409556, 32'sd-0.09270572141975847, 32'sd-0.06072078217601771, 32'sd0.06821368596106922, 32'sd-0.06832349429299585, 32'sd0.01650074466910924, 32'sd-0.04167394870158497, 32'sd0.1312503031432787, 32'sd0.12270795951608436, 32'sd0.04683579223832583, 32'sd-0.04385081419720166, 32'sd-0.0006935805669818659, 32'sd0.01716426230414684, 32'sd0.013752496884011324, 32'sd0.030945379042386215, 32'sd-0.05645839582394019, 32'sd-0.13091443968988833, 32'sd0.038225704083912314, 32'sd-0.03490125280683452, 32'sd0.046642463347356694, 32'sd-0.13428680491693026, 32'sd0.04427986873559337, 32'sd0.04765830756239304, 32'sd-0.03870357957609465, 32'sd-0.12427984202801633, 32'sd-0.07088319342685374, 32'sd0.16708232343253906, 32'sd-0.001425472837941155, 32'sd-0.13975801327005694, 32'sd-0.12388797053919036, 32'sd-0.15185081535559897, 32'sd0.01602568317613826, 32'sd0.01810574680981159, 32'sd0.007574994901834061, 32'sd0.013353293973062669, 32'sd-0.008299441064602819, 32'sd0.0605592136737731, 32'sd0.014826728391586039, 32'sd-0.00011716908270768594, 32'sd0.07285405443351428, 32'sd0.04634137226491836, 32'sd-0.04026211079448035, 32'sd0.04243880930277351, 32'sd0.05680253005107063, 32'sd0.06590566020432073, 32'sd0.14321244515605916, 32'sd0.008825216585859852, 32'sd0.010635635137061355, 32'sd0.016229941655657467, 32'sd0.009209968948532805, 32'sd0.1118250174639791, 32'sd-0.05963723070242757, 32'sd0.020070262835717417, 32'sd-0.09123082022211271, 32'sd0.013358832563581087, 32'sd-0.12486943796176209, 32'sd-0.14470791504703917, 32'sd-0.1531041980126751, 32'sd-0.07717137318369494, 32'sd-0.06222653886607931, 32'sd-0.034250512273645096, 32'sd0.0013091421554907892, 32'sd0.08707369204973739, 32'sd0.07571872998801013, 32'sd0.0861937851364097, 32'sd0.013015208776947519, 32'sd-0.07108145972188659, 32'sd0.05683570594466269, 32'sd0.07209400566071622, 32'sd-0.0692875195513121, 32'sd0.034467804001933285, 32'sd-0.11090570360148722, 32'sd0.005716206276391571, 32'sd0.05043929042477383, 32'sd0.0284470615656904, 32'sd-0.03598304577307567, 32'sd-0.0047654062143183285, 32'sd0.06079107777257569, 32'sd-0.019851186381016447, 32'sd-0.05772842079946775, 32'sd-0.06422411812876504, 32'sd0.08246886989387911, 32'sd0.02195297416671902, 32'sd-0.15108545575933227, 32'sd-0.20426167846199156, 32'sd-0.08550901845588127, 32'sd-0.016448538908295493, 32'sd0.10050970240022078, 32'sd-0.05053096351860765, 32'sd-0.03545997670277687, 32'sd-0.013792294519679631, 32'sd-0.028759359200122396, 32'sd-0.07806183126510872, 32'sd-0.08375860885997993, 32'sd-0.019865881703128, 32'sd0.04022039451949784, 32'sd0.03025969908897544, 32'sd0.057245956130178105, 32'sd-0.06452240467726049, 32'sd-0.10883543012398264, 32'sd-0.039722983310934434, 32'sd0.08216915545392448, 32'sd0.028037399735507867, 32'sd-0.0773712498869289, 32'sd-0.13437716797042465, 32'sd-0.07726346368867526, 32'sd-0.05057728925056443, 32'sd-0.18688200741655134, 32'sd-0.06146056774430665, 32'sd0.06385883566206318, 32'sd0.11814049112832516, 32'sd-0.09361202664578838, 32'sd-0.22535381521069653, 32'sd-0.08843741950682464, 32'sd0.0011553953868401127, 32'sd0.012523788958222122, 32'sd-0.04872375714380406, 32'sd0.002241690309088715, 32'sd-0.020456739589340987, 32'sd-0.011205164810546868, 32'sd-0.08528226570689898, 32'sd0.015060618376467074, 32'sd0.04085952295485229, 32'sd-0.019244559917043033, 32'sd6.762994907278849e-116, 32'sd-0.0015199918102724468, 32'sd0.0033109140511149225, 32'sd-0.14380216632889256, 32'sd0.06136876958722622, 32'sd-0.0020349250777306066, 32'sd0.03672512079036577, 32'sd-0.08657863890425327, 32'sd-0.026015792338491883, 32'sd-0.0711368603049913, 32'sd-0.11576407271509145, 32'sd-0.06371272587080011, 32'sd-0.0788324594516189, 32'sd-0.05417475088083694, 32'sd0.1580061470921332, 32'sd0.055421214383528386, 32'sd-0.01208219152440933, 32'sd0.026043885428399787, 32'sd-0.035640393202864266, 32'sd0.021908894982760576, 32'sd0.036149516180929445, 32'sd-0.02018579753180296, 32'sd0.01076670681180184, 32'sd-0.005321700488285469, 32'sd-0.06771041818828316, 32'sd-0.02575179067781273, 32'sd-0.04507006766491042, 32'sd0.023245156706180093, 32'sd0.036074703139200845, 32'sd0.05009590427854066, 32'sd0.03916161652077676, 32'sd-0.08179157372408251, 32'sd-0.04112128832545355, 32'sd0.07192782318336699, 32'sd0.07579027697961338, 32'sd-0.08607009883701046, 32'sd-0.05579140792707119, 32'sd0.016799691474542307, 32'sd0.010828533275839606, 32'sd-0.18389546415735736, 32'sd-0.052471878155586335, 32'sd0.028218443811661234, 32'sd0.19509674571232308, 32'sd0.005017736417485962, 32'sd0.04159708680782173, 32'sd-0.01670252987910795, 32'sd0.03758332402846048, 32'sd-0.092601408757397, 32'sd-0.025362205507933236, 32'sd-0.03157178573409213, 32'sd0.04551714369051748, 32'sd-0.0059008430840047634, 32'sd0.13883408020260757, 32'sd-0.03121675598513552, 32'sd-0.07258103343333028, 32'sd-0.01598397350843732, 32'sd0.03150867678025974, 32'sd0.07054888536384951, 32'sd-0.11838286101492944, 32'sd-0.06988525718705413, 32'sd-0.11566675578097613, 32'sd0.0837532699111663, 32'sd0.08863647406371838, 32'sd0.058751599112235105, 32'sd0.024474523060338923, 32'sd-0.011508194581250027, 32'sd-0.017933538516737096, 32'sd0.043499023255527756, 32'sd0.04433667212968601, 32'sd0.2099834303885589, 32'sd0.20723542500487513, 32'sd0.04622421997615392, 32'sd-0.042719513831985245, 32'sd-0.03885294228509601, 32'sd-0.09205897342918433, 32'sd-0.06957769462296665, 32'sd0.03845019497891892, 32'sd-0.06569561899263965, 32'sd0.020755998308603654, 32'sd-0.015073453349059185, 32'sd-0.02193659469271894, 32'sd0.023176397969652773, 32'sd-0.11866536873834999, 32'sd-0.006895039456235233, 32'sd-5.136923237408402e-117, 32'sd0.010135062132307535, 32'sd-0.02272162428038178, 32'sd-0.05529198436230017, 32'sd-0.0025935828873172454, 32'sd0.1256403845773489, 32'sd0.04043051965633881, 32'sd-0.07473653339213437, 32'sd-0.1523420810465341, 32'sd-0.04557311899401764, 32'sd-0.08377727365595608, 32'sd0.10795128355081841, 32'sd0.16408422234219114, 32'sd0.18903942607002105, 32'sd0.05518771997030872, 32'sd0.1665895598124557, 32'sd0.04268089742804406, 32'sd-0.10144809089760644, 32'sd0.017234285845719323, 32'sd-0.0003187027753932638, 32'sd-0.07648597077448319, 32'sd-0.11404565324967354, 32'sd-0.004777661937663869, 32'sd-0.02887610527847701, 32'sd0.008010562126571875, 32'sd-0.09509527835007181, 32'sd-0.09141951076538582, 32'sd0.007710214088095978, 32'sd-0.003513785063998238, 32'sd-0.07220323396887587, 32'sd0.05364421238517928, 32'sd0.045873010059216686, 32'sd0.025112402924226937, 32'sd0.0468026072633016, 32'sd0.11680147804472306, 32'sd-0.06566884915555624, 32'sd-0.11520799244127508, 32'sd-0.15097016859260692, 32'sd-0.0024656316263851285, 32'sd0.050075959909789636, 32'sd0.12890759439859426, 32'sd0.11260071043101542, 32'sd0.08965336737266681, 32'sd0.15100617920305737, 32'sd-0.01659753657817513, 32'sd-0.0034808095885398255, 32'sd0.012361181540288976, 32'sd-0.028144568058301848, 32'sd0.030920486057246937, 32'sd0.03043328755702814, 32'sd0.003141648739090746, 32'sd-0.026308930576320673, 32'sd0.060360279354158865, 32'sd-0.10534955633905811, 32'sd0.042829973050616865, 32'sd0.02722265398505814, 32'sd0.11077815587499994, 32'sd0.07145406246114867, 32'sd-0.1284841695272892, 32'sd-0.043427145573171844, 32'sd0.007907507309916169, 32'sd-0.08624949429838932, 32'sd0.0537732863742098, 32'sd0.06412215277494557, 32'sd0.03154475937581273, 32'sd0.027470093943927656, 32'sd0.04739799170921205, 32'sd0.009492677992495532, 32'sd-0.06328786063054453, 32'sd-0.007846598681703846, 32'sd0.09126500819256443, 32'sd0.11163691608897926, 32'sd0.12305443848579332, 32'sd0.01939813118103971, 32'sd0.06786697756623332, 32'sd-0.07535680860284222, 32'sd0.03773660835723556, 32'sd-0.01091876456650612, 32'sd0.06855914663130827, 32'sd-0.013849951626897816, 32'sd0.11713196875024381, 32'sd-0.10638315310917826, 32'sd-0.017898187990778865, 32'sd0.025668504608582512, 32'sd-4.632299452766162e-126, 32'sd0.00037520051095766877, 32'sd0.03487493686927073, 32'sd-0.034474171552035755, 32'sd-0.047002026583620016, 32'sd0.061088691839936995, 32'sd0.06075118866900445, 32'sd-0.009833681504068974, 32'sd0.015281124439664763, 32'sd0.04088542439408856, 32'sd0.028194428744226462, 32'sd-0.027454109833909897, 32'sd-0.04830960138536162, 32'sd-0.045548229729805226, 32'sd0.06231793802341421, 32'sd0.09155078495111857, 32'sd0.10902295462644537, 32'sd0.10026260792758654, 32'sd-0.14593648032745912, 32'sd-0.07568450832915746, 32'sd0.10061849912377366, 32'sd-0.02469983981354213, 32'sd0.07021197683084938, 32'sd-0.04358298188997183, 32'sd0.029897700810334542, 32'sd-0.060902664966082674, 32'sd-0.023883554627883608, 32'sd-1.4299434697933812e-118, 32'sd-9.537954082633708e-120, 32'sd3.856051168264958e-119, 32'sd-0.006685114680582315, 32'sd-0.021301147633536674, 32'sd-0.1053799482138367, 32'sd-0.026243058417426114, 32'sd-0.00017870012218987205, 32'sd-0.041175724612910566, 32'sd0.035012701339591557, 32'sd-0.026278680444321852, 32'sd-0.07741153266920461, 32'sd0.09151492803836234, 32'sd-0.01655709926336672, 32'sd0.019963911889734693, 32'sd-0.08690342649402263, 32'sd-0.04585490065267741, 32'sd0.05993336513994919, 32'sd0.10511434924647878, 32'sd0.10845569541847404, 32'sd0.04731896710798976, 32'sd0.08709854196046173, 32'sd-0.05104701626884038, 32'sd-0.010739838282689117, 32'sd0.035441465700594706, 32'sd0.06915729282876434, 32'sd0.016262040747687046, 32'sd-0.050313704013833595, 32'sd-3.504440916886034e-118, 32'sd-1.1275665463767658e-119, 32'sd1.8173208698329712e-123, 32'sd-0.050208482669456274, 32'sd0.10520558568447212, 32'sd0.006074943549940304, 32'sd0.014886926308425131, 32'sd0.05753413210854033, 32'sd0.10610805040486622, 32'sd-0.0998615458055132, 32'sd-0.10971482044613148, 32'sd-0.1512358502239909, 32'sd-0.007762629052997417, 32'sd-0.009823583579391023, 32'sd-0.010348420864192163, 32'sd-0.010313144364783512, 32'sd-0.056437561156745274, 32'sd0.021454939281549405, 32'sd0.09779648837304712, 32'sd0.10031288623265484, 32'sd-0.032471936998447574, 32'sd0.055473674354134514, 32'sd0.04713496442529571, 32'sd0.013277974854016395, 32'sd0.046904111585063704, 32'sd0.07612260495295826, 32'sd0.04833412803768767, 32'sd0.025934047139901918, 32'sd-7.831466259091532e-122, 32'sd2.4432196421724697e-120, 32'sd-8.514003871104247e-117, 32'sd-2.9629886698652646e-123, 32'sd0.05398620498455255, 32'sd0.02815485885155402, 32'sd0.018793717164746936, 32'sd0.01841983144892066, 32'sd0.0715865934567064, 32'sd0.12367198230817258, 32'sd0.013759584559931197, 32'sd0.02867139711387309, 32'sd0.054366223833412906, 32'sd-0.10598682756300674, 32'sd-0.07024045249522261, 32'sd0.04738804087256013, 32'sd0.10471345017752931, 32'sd0.007920074754715779, 32'sd-0.1358132412524612, 32'sd-0.0034580811308491575, 32'sd-0.05889257871616996, 32'sd0.03699462348280159, 32'sd-0.12583538779787007, 32'sd-0.07345292705899287, 32'sd0.01707314431122076, 32'sd0.07653517622684329, 32'sd0.00422440856088464, 32'sd-6.878233147311448e-124, 32'sd1.4262392706475576e-122, 32'sd-9.857992123709217e-121, 32'sd2.5132428685688463e-116, 32'sd2.6600567342375505e-124, 32'sd4.311209763372958e-122, 32'sd0.013109433212931601, 32'sd0.041596584072382044, 32'sd0.0857728076435945, 32'sd-0.06254896612946398, 32'sd0.049598551416426856, 32'sd-0.01642165230021805, 32'sd0.04551135593814263, 32'sd0.061666570404211384, 32'sd0.042932251289854305, 32'sd0.0519887888940412, 32'sd-0.03975157767604816, 32'sd0.045855600328566684, 32'sd0.036587011597508094, 32'sd0.052035225046313555, 32'sd-0.03778322876428211, 32'sd0.014225701025670511, 32'sd-0.027292682055229566, 32'sd-0.06258683788424593, 32'sd-0.059450616641794296, 32'sd0.047675705319445975, 32'sd3.517566431363039e-119, 32'sd9.878795128523307e-125, 32'sd3.393564779451949e-120, 32'sd-1.4386226843646451e-123},
        '{32'sd-7.382731741296083e-115, 32'sd-3.08654917348385e-116, 32'sd6.274868762279328e-124, 32'sd-2.3852152784808256e-120, 32'sd4.0740931366548166e-120, 32'sd3.0664801851244664e-114, 32'sd-1.3114945064478622e-122, 32'sd-1.0749444178224322e-122, 32'sd-2.9004115930175244e-118, 32'sd-1.558362876582376e-115, 32'sd5.6019823624733426e-121, 32'sd1.7413093981659968e-124, 32'sd0.03593551953457973, 32'sd-0.06455326571341057, 32'sd0.02528551400409072, 32'sd-0.06281194862183231, 32'sd3.1895546559889024e-122, 32'sd-1.1933586041551465e-118, 32'sd2.9752305664727153e-120, 32'sd3.36863443574848e-120, 32'sd-8.632504874673312e-119, 32'sd-4.620250740231205e-118, 32'sd1.572326716590439e-123, 32'sd1.0163771384538593e-115, 32'sd-9.884079306387111e-116, 32'sd2.5059142039871994e-124, 32'sd-4.6967184667091724e-117, 32'sd-1.2114641846318098e-118, 32'sd-9.499738383547784e-120, 32'sd1.0437778798145477e-117, 32'sd-2.5503754171643342e-121, 32'sd-4.844911217634635e-118, 32'sd0.06897157710808947, 32'sd0.028987196242506508, 32'sd-0.030160707949772533, 32'sd-0.04091987381120009, 32'sd-0.03736120821088807, 32'sd0.014120736790867658, 32'sd0.050942165640312884, 32'sd-0.019738205791299673, 32'sd-0.002039257336495711, 32'sd0.016393198447518843, 32'sd0.06611488950804315, 32'sd-0.04132245530751839, 32'sd-0.08211880129639089, 32'sd0.028814222398680745, 32'sd-0.07167390437604719, 32'sd0.032644773284774345, 32'sd-0.02316099282458919, 32'sd0.00298002813718725, 32'sd-0.06761193373307153, 32'sd0.014837908472059921, 32'sd-5.009576354684116e-127, 32'sd-2.1365883776612814e-127, 32'sd-1.688898522346423e-125, 32'sd7.673411656982317e-119, 32'sd-4.9023444640673674e-116, 32'sd1.053312617646864e-119, 32'sd0.0020469605585092527, 32'sd-0.020920576717813968, 32'sd0.1138225988734886, 32'sd-0.0016130147273712195, 32'sd-0.02382845042651285, 32'sd-0.06593086009994847, 32'sd0.052758176031962756, 32'sd0.08860624539512768, 32'sd0.04710180011709409, 32'sd0.025621121428216487, 32'sd-0.01536030736191907, 32'sd-0.02497363721291632, 32'sd-0.06074428051952563, 32'sd-0.06387217505270035, 32'sd-0.08990193608671265, 32'sd-0.05917485146463331, 32'sd0.004935193135861935, 32'sd-0.027344854734991927, 32'sd0.03401452314869646, 32'sd-0.028389196660651282, 32'sd-0.010389074898362554, 32'sd0.039197915714517854, 32'sd-0.0462131609472287, 32'sd0.02897596239017973, 32'sd-3.968914732210722e-119, 32'sd-8.630696121479122e-122, 32'sd-7.56717367973444e-115, 32'sd5.930146850589243e-126, 32'sd-0.020685380454963456, 32'sd-0.010485824228043807, 32'sd-0.027534458243497654, 32'sd-0.06122499741851199, 32'sd-0.07318900201008699, 32'sd0.04025060897762235, 32'sd-0.013600227556845465, 32'sd-0.044309358372617166, 32'sd-0.10520515671857904, 32'sd0.010579564287974604, 32'sd-0.03340575322126175, 32'sd-0.0041842877738369425, 32'sd0.1477372239765039, 32'sd-0.015840333845709174, 32'sd-0.16725271497886154, 32'sd-0.049993191557557895, 32'sd-0.11223186676373541, 32'sd-0.07702137038535709, 32'sd-0.07394739745183926, 32'sd0.060941726232771117, 32'sd-0.02283073783495317, 32'sd0.01902895489176401, 32'sd-0.0002532265754825538, 32'sd-0.04838974205879872, 32'sd0.06311127299391849, 32'sd1.3924879638243813e-120, 32'sd4.7850984324764805e-123, 32'sd-0.006648635583214185, 32'sd-0.023294853258100198, 32'sd0.013597073115283796, 32'sd-0.17318999325814685, 32'sd0.020484359301900172, 32'sd0.00499077285378198, 32'sd-0.03025756161850701, 32'sd-0.014158621013231499, 32'sd-0.149685105220724, 32'sd-0.08391543472646272, 32'sd0.002810686264983526, 32'sd-0.0010749060358938578, 32'sd-0.059964279508735056, 32'sd-0.11134834209793436, 32'sd-0.1470360704905551, 32'sd-0.02254955371092002, 32'sd-0.060899979319636886, 32'sd0.0523858066809587, 32'sd-0.05414079352149052, 32'sd-0.014785543942708078, 32'sd0.1234443120278814, 32'sd0.13626120334028455, 32'sd0.02964676394518779, 32'sd-0.04150125291097394, 32'sd0.008332535075822947, 32'sd0.03564954600790963, 32'sd0.0534292039323166, 32'sd4.877888425008389e-119, 32'sd0.02466581016868004, 32'sd-0.04690009066732317, 32'sd0.03755980395492952, 32'sd0.07621425254087168, 32'sd0.012687414321159246, 32'sd0.05831920649653111, 32'sd0.09869028992724459, 32'sd0.08962886802934332, 32'sd-0.03222871344628275, 32'sd0.03967252325054412, 32'sd0.0432696379971518, 32'sd0.06728084909169227, 32'sd0.025470115649257483, 32'sd-0.03638793693488843, 32'sd-0.10879905864366346, 32'sd-0.09109437703004383, 32'sd-0.027783896780351494, 32'sd-0.046118997005539085, 32'sd-0.07242297682351298, 32'sd-0.09593659326465888, 32'sd0.011455334511302729, 32'sd0.06261040722300566, 32'sd0.025933693852599752, 32'sd-0.06751089906474657, 32'sd0.10002536696330408, 32'sd-0.04138626830525991, 32'sd-0.07443450994383166, 32'sd-2.901095957486821e-122, 32'sd-0.0026970564151274673, 32'sd-0.11760900976810908, 32'sd0.047031063090101036, 32'sd0.09438247663645757, 32'sd0.0351461608548458, 32'sd-0.018032437420351047, 32'sd0.0633864020860423, 32'sd0.045825778927505195, 32'sd-0.14110753293429384, 32'sd-0.04359299989701485, 32'sd0.019684927667203856, 32'sd-0.03729882403231426, 32'sd-0.03448159351554842, 32'sd-0.04803799594126019, 32'sd0.032181386239138084, 32'sd0.06938561083994876, 32'sd0.05008830162584427, 32'sd-0.027990329667391036, 32'sd0.04649759988582163, 32'sd0.0637110240468514, 32'sd-0.0025763282846603423, 32'sd-0.006699200439089504, 32'sd0.15246018087354532, 32'sd0.05283966584300511, 32'sd-0.011036550427211063, 32'sd0.09236490113163527, 32'sd-0.002311036246757043, 32'sd0.0255007322221554, 32'sd-0.02638670929062993, 32'sd-0.058004340246290885, 32'sd0.015482409063521184, 32'sd-0.029265000659055206, 32'sd0.003582748345043262, 32'sd-0.08584675628393086, 32'sd-0.11357205571294118, 32'sd-0.09897317707601491, 32'sd-0.1987052376239931, 32'sd0.008148519093536326, 32'sd-0.03045980837614183, 32'sd-0.05891617378877435, 32'sd-0.043613243642113, 32'sd0.07769933007279708, 32'sd0.06124517701397387, 32'sd0.09747381120257591, 32'sd0.05439203619131474, 32'sd-0.06525350018757464, 32'sd0.1568423541864238, 32'sd0.008566338323776823, 32'sd0.048067018249837126, 32'sd0.03535271211747309, 32'sd0.146777909509921, 32'sd0.05909653822649878, 32'sd0.0600042889728155, 32'sd-0.04894569680278559, 32'sd-0.01590797698093643, 32'sd0.06107562604258422, 32'sd0.011024523954049167, 32'sd0.004807611367533129, 32'sd0.09895166545668539, 32'sd-0.13954654990626128, 32'sd-0.03726647875235696, 32'sd-0.07529370742861823, 32'sd-0.061940325259342836, 32'sd-0.10828802417401627, 32'sd0.03476116116380941, 32'sd0.05150868616935957, 32'sd8.347222762764529e-05, 32'sd0.13036650804498068, 32'sd0.10266309531710002, 32'sd-0.020316630085111594, 32'sd-0.019775149819708737, 32'sd-0.15685586224165304, 32'sd-0.11083815198309263, 32'sd0.014908513909943572, 32'sd-0.05254204772379813, 32'sd0.051566749807088245, 32'sd0.007815867091872281, 32'sd0.039465809875253104, 32'sd-0.05122555693623719, 32'sd0.12911001859852542, 32'sd0.09384122034517663, 32'sd0.012703241745962985, 32'sd0.07316453805203305, 32'sd0.040656404552659633, 32'sd0.006967441004482398, 32'sd0.0003965275692576292, 32'sd-0.07987953078553814, 32'sd-0.1668057679232553, 32'sd-0.026543235489147804, 32'sd-0.008756116823786023, 32'sd-0.1391668538550512, 32'sd-0.12017823658536339, 32'sd-0.05367480632887936, 32'sd0.03621831820099179, 32'sd0.05875006230663387, 32'sd0.1815317229705537, 32'sd0.03444939856424875, 32'sd-0.09664145302334529, 32'sd-0.054021634594958595, 32'sd-0.07097851612011283, 32'sd-0.04365011869468381, 32'sd-0.08898172178786716, 32'sd0.0826771221572574, 32'sd0.061456615228653456, 32'sd0.018046734277800777, 32'sd0.012862372302608258, 32'sd-0.05286744324116216, 32'sd0.05661326289870969, 32'sd0.03161239631823375, 32'sd-0.0008839643941701591, 32'sd-0.028968788816699103, 32'sd-0.015676604038244585, 32'sd-0.012022650576266362, 32'sd-0.06370979680966005, 32'sd0.054326724936984136, 32'sd-0.1379671305270435, 32'sd0.0539407311410985, 32'sd-0.05517011726186381, 32'sd-0.11342034122544244, 32'sd-0.14459491511525385, 32'sd-0.034413497150219505, 32'sd0.02655973369178021, 32'sd0.13337783211155815, 32'sd0.0627554665679371, 32'sd-0.16946496415317983, 32'sd-0.19444932871660855, 32'sd-0.19874179030248712, 32'sd-0.1549495954277017, 32'sd-0.10382281634646826, 32'sd-0.10911335413727018, 32'sd0.0838879472306094, 32'sd0.06572162455768879, 32'sd0.0056231148086551995, 32'sd0.11898698493090039, 32'sd0.11514333079149942, 32'sd-0.02723308288992203, 32'sd0.07703839075330578, 32'sd-0.06943453469604643, 32'sd0.024437398814745905, 32'sd-0.0352181399725937, 32'sd-0.06261129329108386, 32'sd0.10803020931191624, 32'sd0.012671283092369727, 32'sd-0.06454717838915357, 32'sd-0.009328143797135069, 32'sd-0.11987574709940876, 32'sd-0.08912932140219078, 32'sd-7.223188893736687e-05, 32'sd0.1467832878073831, 32'sd0.15647778388611325, 32'sd-0.01882409433980064, 32'sd-0.06212501624657856, 32'sd-0.25392725611588934, 32'sd-0.14905419476770282, 32'sd-0.13626720797172384, 32'sd-0.013022429058375808, 32'sd0.030577862271304355, 32'sd-0.0657926374488037, 32'sd0.02172554145935023, 32'sd0.11659657543601809, 32'sd0.12129924409188228, 32'sd0.07123621380733826, 32'sd0.13664201669538395, 32'sd0.04873493949140366, 32'sd0.0321422488015943, 32'sd-0.09863722103283482, 32'sd-0.12408330925271836, 32'sd0.03902771044498512, 32'sd-0.06974003838765558, 32'sd0.06774074296316449, 32'sd0.057305385689078045, 32'sd0.032261952631342565, 32'sd-0.016604695147626053, 32'sd-0.0983487081076525, 32'sd-0.09483336314893939, 32'sd0.09414205147770031, 32'sd0.06477419459495386, 32'sd0.13778300996043114, 32'sd-0.12139419782758358, 32'sd-0.1334805836182858, 32'sd-0.08653819212014435, 32'sd-0.11888544459626917, 32'sd-0.02000319635000072, 32'sd0.1943405506377534, 32'sd0.012770203093594166, 32'sd0.04072882495775687, 32'sd0.1437924679338185, 32'sd0.20489585370368357, 32'sd0.1937129612651938, 32'sd0.09807287016437048, 32'sd0.09205013317817538, 32'sd0.09074586403143421, 32'sd-0.11305513690737047, 32'sd-0.06887734397090418, 32'sd0.007521019964717577, 32'sd-0.0013942599426303296, 32'sd-0.007271678083599267, 32'sd-0.032545660247128703, 32'sd-0.08277596443063236, 32'sd-0.048246838530149785, 32'sd-0.14316543825535713, 32'sd-0.040263908541850586, 32'sd0.06369687186132907, 32'sd0.06488110634715515, 32'sd0.09954990963936151, 32'sd-0.07613871461984636, 32'sd-0.02333908944509296, 32'sd0.045374055702092325, 32'sd0.00389786629545069, 32'sd0.1305618017870471, 32'sd0.29368138729264853, 32'sd0.07122380959593608, 32'sd0.0496148095636474, 32'sd0.008688217264625455, 32'sd0.04966334595009615, 32'sd0.1029092084364947, 32'sd0.12650936282873848, 32'sd0.042701517913906153, 32'sd0.0725158241353346, 32'sd-0.027536688789447684, 32'sd-0.10690829613611491, 32'sd-0.11628926368204805, 32'sd0.03381248470001651, 32'sd0.04443151510581478, 32'sd0.037161376971175115, 32'sd-0.007373036128931075, 32'sd-0.0474322771109221, 32'sd-0.012005698581212398, 32'sd-0.0464014223613209, 32'sd-0.1846653601495665, 32'sd0.053969439338939766, 32'sd-0.039258947843534515, 32'sd-0.021902673592846228, 32'sd-0.07599087512321955, 32'sd-0.032016069826702444, 32'sd0.032282477704712105, 32'sd0.2757205095248918, 32'sd0.1964486640920359, 32'sd0.18654885691235304, 32'sd0.1596100357598424, 32'sd0.06792032954763823, 32'sd-0.022355983773863913, 32'sd0.014014447517807883, 32'sd0.07782202887597672, 32'sd0.02238501464495827, 32'sd-0.06307609294328598, 32'sd-0.03626110331074568, 32'sd-0.12364543041902626, 32'sd0.04032514568679231, 32'sd-0.03839890688351406, 32'sd-0.026242817455029068, 32'sd0.02787389329937602, 32'sd0.06070707762253129, 32'sd-0.04896159634612808, 32'sd0.02187978671289167, 32'sd-0.08028744995604524, 32'sd-0.0769038698074719, 32'sd-0.050123094378283155, 32'sd0.008322893748960461, 32'sd0.04238622149241624, 32'sd-0.07897712929226519, 32'sd-0.017377587225107082, 32'sd0.08300375728588182, 32'sd0.09093183022211779, 32'sd0.12474546900964502, 32'sd0.2875480033178878, 32'sd0.1783738773672373, 32'sd0.15191981471603574, 32'sd0.03127422063150046, 32'sd0.03900803468472279, 32'sd-0.1447450998538807, 32'sd-0.14253025244172216, 32'sd-0.021777993679851917, 32'sd0.031310024476536885, 32'sd0.04161383276673798, 32'sd-0.041553637084474085, 32'sd-0.07264628500077124, 32'sd0.06308133422944238, 32'sd0.05573042449129611, 32'sd0.0004820832763690228, 32'sd0.06570608694937541, 32'sd-0.03052714799415066, 32'sd0.02868219528574874, 32'sd0.07176988239096367, 32'sd-0.033010069728658144, 32'sd-0.0638141940840452, 32'sd0.03211112431045028, 32'sd0.03881486791225786, 32'sd-0.01802815994125822, 32'sd0.05718243605366281, 32'sd0.0341141989976846, 32'sd0.20143048709949915, 32'sd0.21985739838401136, 32'sd0.10953667952251567, 32'sd0.018471393984759735, 32'sd-0.010334195803432205, 32'sd-0.057356998460802326, 32'sd-0.10751949326769791, 32'sd-0.12328544102469519, 32'sd-0.004278415472813309, 32'sd0.020635271248957174, 32'sd-0.058147403872697775, 32'sd0.07553387765768606, 32'sd0.07628383354906074, 32'sd-0.07899308854532468, 32'sd0.017180328990572136, 32'sd0.08153459427735517, 32'sd3.0022361489924304e-123, 32'sd-0.023823966363826655, 32'sd-0.09712063053097605, 32'sd-0.00874353795896392, 32'sd0.029444167472209695, 32'sd-0.16773232026113286, 32'sd-0.13826288275639964, 32'sd0.020685067767373725, 32'sd0.02026367913338615, 32'sd-0.18569586058774554, 32'sd-0.025598359738003035, 32'sd0.07415357448654655, 32'sd0.09295518281774957, 32'sd0.16037860255963157, 32'sd0.045674198914857765, 32'sd-0.016568069465795275, 32'sd-0.05707952858120656, 32'sd-0.131686842484223, 32'sd-0.14114066349200113, 32'sd-0.0357945461818087, 32'sd-0.11890223376272081, 32'sd-0.01639104249181645, 32'sd0.003593159483360799, 32'sd-0.06282922189790184, 32'sd-0.14696420728124443, 32'sd-0.005764497185882569, 32'sd-0.07042208051109448, 32'sd-0.10357057487291677, 32'sd0.0026504891877725052, 32'sd0.050056730978095536, 32'sd-0.06848818890605847, 32'sd-0.13151927712063174, 32'sd-0.07377420707622095, 32'sd-0.1187397430251029, 32'sd-0.10806810482393277, 32'sd-0.008261700958726113, 32'sd-0.08589090478496124, 32'sd0.013584358121439094, 32'sd-0.015704633988030476, 32'sd0.09806552846293994, 32'sd-0.035968929612210876, 32'sd0.024424943353279008, 32'sd0.09709390286754106, 32'sd0.06570270446708508, 32'sd-0.12413325135224428, 32'sd-0.18681850252956708, 32'sd-0.1066573600855481, 32'sd-0.04305083117651977, 32'sd-0.10132955953882905, 32'sd-0.09654817189952726, 32'sd-0.09925404073445146, 32'sd-0.04975693477790993, 32'sd-0.06619675724292044, 32'sd0.0039359903868922685, 32'sd0.03572961088283031, 32'sd0.06672463807490786, 32'sd0.011766814198002873, 32'sd-0.04658985746812418, 32'sd0.08721786721732369, 32'sd-0.02211948503693079, 32'sd0.003828889556446194, 32'sd-0.06585769175811053, 32'sd-0.05712980297626594, 32'sd-0.021265271147321952, 32'sd-0.0873913157099935, 32'sd0.022654779182943684, 32'sd0.015931158747184194, 32'sd-0.07991526513580358, 32'sd-0.04902590751957333, 32'sd0.05781747545960411, 32'sd0.23631975033716474, 32'sd-0.026089419934080472, 32'sd-0.10069361531114851, 32'sd-0.018804932743221908, 32'sd0.008511741306729825, 32'sd0.055764415053473786, 32'sd-0.06844517624715812, 32'sd0.04394461824096313, 32'sd-0.027279699034990237, 32'sd-0.1498958838985914, 32'sd-0.022428719333916478, 32'sd-0.03385381574612902, 32'sd0.07912869708661001, 32'sd0.008745276387480648, 32'sd-8.08824320495131e-123, 32'sd0.046875485505713375, 32'sd0.10408347453588714, 32'sd-0.05642326507184003, 32'sd0.019538057930147772, 32'sd0.005129920733295539, 32'sd-0.026431892972542458, 32'sd0.03971910036894139, 32'sd-0.04940066170873357, 32'sd-0.11302396246490164, 32'sd-0.03103955919038215, 32'sd-0.1434782903952584, 32'sd0.00976295193079742, 32'sd0.12630796914216694, 32'sd0.20159427462097634, 32'sd0.07941112157716497, 32'sd-0.06574252415164167, 32'sd0.004083852054597783, 32'sd-0.005217612193553367, 32'sd-0.05034099765462764, 32'sd-0.030649215332224804, 32'sd0.004300239616013014, 32'sd-0.04878804547300405, 32'sd-0.008400487218540536, 32'sd-0.03649884962228944, 32'sd0.06990722662453268, 32'sd0.08182118823728794, 32'sd-0.04076200127558456, 32'sd0.0009771072238521936, 32'sd0.001964467355553217, 32'sd-0.008116562973213717, 32'sd0.07190346841330202, 32'sd-0.014380969284673337, 32'sd-0.058778322324168276, 32'sd0.06136291924830777, 32'sd0.001034684796329164, 32'sd-0.11317333504695838, 32'sd0.01579019119051412, 32'sd-0.01563592269059748, 32'sd-0.018686891307651016, 32'sd0.04044797298134506, 32'sd0.03705947899938416, 32'sd0.014218556605071738, 32'sd-0.022339402910550914, 32'sd-0.12975586169425027, 32'sd-0.237559230708794, 32'sd-0.03180312249043321, 32'sd-0.11290888044676539, 32'sd-0.0370945725858769, 32'sd-0.0631174170554903, 32'sd-0.05259030768957825, 32'sd0.053559284485290654, 32'sd-0.10529794169781796, 32'sd-0.05282304639010733, 32'sd0.004265789608217207, 32'sd0.013294976011580872, 32'sd0.08670812057563472, 32'sd0.00488004963776967, 32'sd-0.032537409613397864, 32'sd-0.10772626889943149, 32'sd0.00018308171290159093, 32'sd-0.03451413792268433, 32'sd0.1680589834699379, 32'sd0.09578013774705377, 32'sd-0.02990022265425742, 32'sd-0.06845318649255215, 32'sd0.030706579522830974, 32'sd0.005314048365014071, 32'sd-0.00973007607524094, 32'sd-0.04775699750235062, 32'sd0.09217790541623055, 32'sd-0.18329499484478678, 32'sd-0.3015898471317711, 32'sd-0.36177770220827854, 32'sd-0.10376288098101476, 32'sd-0.006516174332592304, 32'sd-0.058811914933533514, 32'sd-0.027578920144548685, 32'sd-0.04613542772281426, 32'sd-0.03367450066857431, 32'sd-0.006245185278597423, 32'sd-0.0017919345880029786, 32'sd-0.035873183291771873, 32'sd0.020798663903236543, 32'sd3.976528296517856e-117, 32'sd0.00347914758263012, 32'sd-0.021595879173111385, 32'sd0.03866330573332653, 32'sd-0.1200040219865396, 32'sd0.08542096898905237, 32'sd0.021500602391007883, 32'sd0.04681288769997221, 32'sd0.1664237282811724, 32'sd-0.032546038434303655, 32'sd0.07017445638297237, 32'sd0.07565660409486102, 32'sd-0.08344034701348275, 32'sd-0.08908253006878915, 32'sd0.008890674346782399, 32'sd-0.24818378427023743, 32'sd-0.22312089722581546, 32'sd-0.2400116054140103, 32'sd-0.011772564431894415, 32'sd-0.1672549025518825, 32'sd-0.08385922141971208, 32'sd-0.0450819491457144, 32'sd-0.08344783361671052, 32'sd0.017962340824783415, 32'sd0.03256767753948059, 32'sd0.01811548769700683, 32'sd0.005997851033402956, 32'sd6.2361512858829464e-117, 32'sd3.5359786329305106e-114, 32'sd-1.9903706257005845e-129, 32'sd0.08464329735479204, 32'sd-0.1432197251496791, 32'sd-0.05598118365267417, 32'sd0.0346512642829816, 32'sd-0.0073554896539753094, 32'sd-0.055440790124634626, 32'sd0.07390991796397745, 32'sd0.03777112191594569, 32'sd0.056702061331194244, 32'sd-0.03060486157468723, 32'sd0.010716546634477549, 32'sd0.023981537682064, 32'sd0.1672892715350891, 32'sd0.054143619219053585, 32'sd-0.07614569115843899, 32'sd-0.23250103004329759, 32'sd0.014600806507219954, 32'sd-0.045906142503648814, 32'sd-0.0325754173882102, 32'sd0.054480785073269304, 32'sd0.07077788705712876, 32'sd0.09274241053645194, 32'sd0.04964630244067555, 32'sd0.0017618105038847288, 32'sd0.048393246059976594, 32'sd3.1754097985556417e-116, 32'sd-4.406753652507551e-123, 32'sd-5.383791013204291e-118, 32'sd0.055132688482175125, 32'sd-0.10922718493431968, 32'sd-0.019498925627942018, 32'sd0.0306309170143, 32'sd-0.011027735527976517, 32'sd0.05621386655695153, 32'sd0.021357127471231804, 32'sd-0.020777056771007836, 32'sd-0.020660951214666764, 32'sd0.045592122651083214, 32'sd-0.06037807784114766, 32'sd0.023911189841137114, 32'sd0.010577344418423076, 32'sd-0.023072993162168594, 32'sd-0.03475765100327499, 32'sd-0.11448980192880948, 32'sd0.08927280998828944, 32'sd0.028108943296619216, 32'sd-0.0639269991108289, 32'sd-0.13470181043152507, 32'sd0.028067192624434988, 32'sd0.03049579574746439, 32'sd-0.0644722635922239, 32'sd0.03918073144938076, 32'sd-0.0013043904955503769, 32'sd-1.3798392654271456e-115, 32'sd-2.3951611796857957e-124, 32'sd3.6668125748179616e-119, 32'sd3.547898531652776e-123, 32'sd0.037571860328596496, 32'sd0.028545891854245994, 32'sd0.06083143054669173, 32'sd-0.02619858504631945, 32'sd-0.004209599171631595, 32'sd0.027304738833037297, 32'sd0.022846910617036052, 32'sd0.06977307753876975, 32'sd0.12323899471533387, 32'sd0.10695474348231207, 32'sd0.11954313066100603, 32'sd0.06392919036651228, 32'sd-0.017613021804233076, 32'sd0.020551996019726078, 32'sd0.054372772597615526, 32'sd0.14388782680798853, 32'sd0.0025656587461353455, 32'sd0.04283938371685788, 32'sd-0.04170453738791843, 32'sd0.03774202775365244, 32'sd0.005188483795323415, 32'sd0.055075800173527915, 32'sd0.05170709376317549, 32'sd-2.7258549031171525e-120, 32'sd-3.097019404832373e-119, 32'sd2.8820245614068053e-115, 32'sd1.772965128498441e-116, 32'sd-2.0632811661105602e-126, 32'sd-6.575002108709592e-124, 32'sd0.03049697323977652, 32'sd0.05461822398484115, 32'sd0.010760349314220206, 32'sd0.003534777577786361, 32'sd0.024821122510995983, 32'sd-0.002613266856018199, 32'sd0.0232241376019245, 32'sd0.009577595709191112, 32'sd0.059611339773706334, 32'sd0.010895763345229428, 32'sd0.06093373509631367, 32'sd0.06101602039582476, 32'sd0.13716846734901542, 32'sd0.00918335033365622, 32'sd0.13573535935229697, 32'sd-0.0021069219371206275, 32'sd-0.027819775905217278, 32'sd0.014578032347374826, 32'sd0.011587452027999436, 32'sd0.005656383256070148, 32'sd-1.5596117760744503e-115, 32'sd-4.67325051207548e-117, 32'sd1.1526519373800116e-125, 32'sd-7.871217440455424e-116},
        '{32'sd-6.567396500981041e-124, 32'sd-1.8381107648602545e-124, 32'sd-6.97702759622446e-121, 32'sd-4.051284432712837e-125, 32'sd1.2250487652424049e-115, 32'sd6.90603866550868e-121, 32'sd5.7474385799412385e-123, 32'sd-8.951463925882333e-121, 32'sd2.1242172049319907e-127, 32'sd3.054612874515979e-126, 32'sd-4.001607669812232e-130, 32'sd5.451639810406055e-117, 32'sd0.07991779365792082, 32'sd0.059227243173999224, 32'sd0.08056688567183043, 32'sd-0.027908032451118177, 32'sd4.243024659487106e-123, 32'sd9.730403265775987e-123, 32'sd2.4280066472255936e-123, 32'sd1.6784328341826533e-125, 32'sd1.9095515904393722e-118, 32'sd6.945871207340902e-127, 32'sd2.48669200010424e-125, 32'sd-3.8778145371754586e-119, 32'sd6.42701459481325e-126, 32'sd-3.343753204121962e-123, 32'sd-1.5147417047311836e-126, 32'sd-1.5629888054117688e-115, 32'sd-1.9938480212994436e-124, 32'sd-6.886931607588972e-124, 32'sd7.015157748327062e-120, 32'sd-9.717439412497161e-118, 32'sd0.007873646538059439, 32'sd0.05371085184671167, 32'sd-0.031656418042275015, 32'sd0.033429117942991714, 32'sd0.00022693836737977492, 32'sd0.08460472110276408, 32'sd-0.050989640457284914, 32'sd-0.048069442528498506, 32'sd-0.016751299620183582, 32'sd0.008860493073569618, 32'sd-0.018844528351777527, 32'sd-0.008894178361805817, 32'sd0.09998362994272973, 32'sd0.10069743143581873, 32'sd0.09245904371857255, 32'sd0.014946962765189835, 32'sd0.0975086226147354, 32'sd0.13166938714141938, 32'sd0.06915191285793557, 32'sd0.04290138153289246, 32'sd1.4311928534510202e-118, 32'sd-3.888476998813347e-119, 32'sd3.2020084864435285e-124, 32'sd2.1177662374351284e-117, 32'sd-8.630992547063356e-117, 32'sd-1.1791808557329178e-115, 32'sd0.07949325330537844, 32'sd0.04913059105131639, 32'sd-0.09595600718624944, 32'sd0.01370793042187003, 32'sd0.03796027295069339, 32'sd0.07562334806612594, 32'sd0.027680130913198507, 32'sd-0.04789627877110561, 32'sd0.025299477678144815, 32'sd-0.01029419311805109, 32'sd-0.04413186261869604, 32'sd-0.07477266268913316, 32'sd0.10347572854969125, 32'sd0.07606667349028205, 32'sd0.045386582834703995, 32'sd0.06526324999924912, 32'sd-0.02534215951761483, 32'sd-0.060550225796012755, 32'sd0.025812923341679277, 32'sd0.14984519804521879, 32'sd0.0867815331140866, 32'sd0.08682241467056771, 32'sd0.13223622462255508, 32'sd0.07088721209730711, 32'sd1.133417021179394e-118, 32'sd3.01446633113289e-125, 32'sd2.6035861133751515e-115, 32'sd1.7022317066268751e-127, 32'sd0.019228005926091793, 32'sd0.08092017980433451, 32'sd0.06469522318712473, 32'sd0.032347280966643584, 32'sd-0.050290345867143, 32'sd-0.0004379797407354909, 32'sd0.09486003887024157, 32'sd0.10557035530692226, 32'sd0.01988957440926107, 32'sd0.11412714822945971, 32'sd0.05147011827085626, 32'sd0.028159686407267417, 32'sd0.014568572795423415, 32'sd0.03532057210172966, 32'sd0.03214040629332733, 32'sd-0.004474005276388976, 32'sd0.027353849501786986, 32'sd-0.07080003387100509, 32'sd-0.09637347538564399, 32'sd-0.013275591910446152, 32'sd-0.004828452752046354, 32'sd0.0020751072617973118, 32'sd0.11620915221125994, 32'sd0.02102272707924667, 32'sd0.0020284325757819062, 32'sd1.0984606025489672e-117, 32'sd1.5300476160022303e-123, 32'sd0.0491077615899661, 32'sd-0.016734045895772206, 32'sd0.02540263141011368, 32'sd0.07028850746212159, 32'sd0.024516492512010223, 32'sd0.02266846085286791, 32'sd-0.017991291734210848, 32'sd0.07992783522313343, 32'sd-0.052730044467321206, 32'sd-0.03711759416681431, 32'sd0.10125616241498778, 32'sd0.08306152502031997, 32'sd0.005224290490554454, 32'sd0.017089765827408662, 32'sd0.0030426484734969476, 32'sd0.004064450862474785, 32'sd-0.039230450758650046, 32'sd-0.00581920067716424, 32'sd0.07362851747532866, 32'sd-0.00225226944186217, 32'sd-0.03574699322658745, 32'sd-0.06516900108822657, 32'sd-0.08205473980064774, 32'sd-0.03965256422576516, 32'sd0.0016255786212540362, 32'sd0.04380105054884713, 32'sd0.07451992376799041, 32'sd-2.3259589284588818e-127, 32'sd0.07535955583998706, 32'sd-0.01736198570645516, 32'sd-0.05256018593557932, 32'sd0.02003615692213382, 32'sd-0.062488654295696805, 32'sd0.12744679832532316, 32'sd0.10278312973963234, 32'sd0.11278199729736586, 32'sd0.017863121101317683, 32'sd0.19622062938756246, 32'sd0.21017404731412623, 32'sd0.1264756383167639, 32'sd0.060400486456301944, 32'sd-0.05639163775349521, 32'sd-0.12764287315823353, 32'sd0.005476089402930895, 32'sd-0.07489159650825968, 32'sd-0.017813847590434643, 32'sd0.047988262817437434, 32'sd0.07293399611641661, 32'sd0.020929371668791365, 32'sd-0.07342404871640364, 32'sd-0.03905055842641002, 32'sd-0.16959704814044127, 32'sd-0.10186126901102557, 32'sd-0.021123936595043486, 32'sd-0.0033296099002960143, 32'sd1.5832032329317917e-127, 32'sd0.05633540449208943, 32'sd-0.01369575563229655, 32'sd-0.01349560723798649, 32'sd-0.07721154963701307, 32'sd0.03613143236087543, 32'sd0.022888333269768763, 32'sd-0.00337064973044598, 32'sd0.09937074879842776, 32'sd0.22146046935334646, 32'sd0.19029912861793952, 32'sd0.21102345141797418, 32'sd0.0635732311697294, 32'sd0.09844535332865745, 32'sd0.05309471879668871, 32'sd0.1334740527179649, 32'sd0.12319811071298878, 32'sd0.025473505316669403, 32'sd-0.04192878999030989, 32'sd0.05609220674877514, 32'sd-0.022601518309639, 32'sd0.023840237459163076, 32'sd0.03890238207310497, 32'sd-0.009388783579963459, 32'sd0.00998274451563969, 32'sd-0.003583877525423501, 32'sd0.044838261201050535, 32'sd-0.08567569950383513, 32'sd0.12915650622959854, 32'sd0.020284558050929515, 32'sd-0.02111576798357695, 32'sd0.06406791702433819, 32'sd-0.0009833964703730774, 32'sd-0.04751744952808008, 32'sd0.0661559261365421, 32'sd0.13703018966015476, 32'sd-0.056208727675881885, 32'sd0.06612647556304102, 32'sd0.11755511860174651, 32'sd0.15074401584823113, 32'sd0.16164005417866695, 32'sd0.14794620690983148, 32'sd0.16391654335969216, 32'sd0.03268740346924974, 32'sd0.09227138773183276, 32'sd0.07397938035581282, 32'sd0.029175932496276136, 32'sd0.16619261412204342, 32'sd0.10915810560917817, 32'sd0.03225674593677048, 32'sd-0.06454495710309821, 32'sd-0.01489119993464323, 32'sd0.12482323123428694, 32'sd0.09241608195651807, 32'sd0.1456026813013802, 32'sd-0.01863347760418871, 32'sd0.045865401060226546, 32'sd0.07127155457619926, 32'sd-0.1103797496030645, 32'sd0.08424766656407376, 32'sd-0.026472689136067873, 32'sd-0.018767219409833998, 32'sd-0.06964464751388781, 32'sd0.01973915686688684, 32'sd-0.03690791350854842, 32'sd-0.09616675013878502, 32'sd-0.06383585916583542, 32'sd0.049860691457493146, 32'sd-0.03788919735633797, 32'sd0.02462265512156192, 32'sd0.12474334070997446, 32'sd0.0669126712432863, 32'sd0.03694194153228147, 32'sd0.018461076508574033, 32'sd0.04308132061878264, 32'sd0.07779099972127179, 32'sd0.0027839092536644607, 32'sd0.03210034340039998, 32'sd0.008596414966562951, 32'sd0.047639106780977235, 32'sd0.028828146840776083, 32'sd-0.03255289103768322, 32'sd0.07497714955511853, 32'sd-0.05230065678898117, 32'sd0.03410994702882004, 32'sd-0.11468404113874973, 32'sd-0.07931914020466489, 32'sd0.011941297775858482, 32'sd0.02096884380896451, 32'sd-0.021331499291530744, 32'sd-0.11408280513859363, 32'sd0.0986933690721462, 32'sd-0.13366872721991255, 32'sd-0.17840398463972304, 32'sd-0.25157007831986605, 32'sd-0.11872146521659621, 32'sd-0.176568651218239, 32'sd-0.19818092126378614, 32'sd-0.19960039090317466, 32'sd-0.06388123352575122, 32'sd-0.018946112116252904, 32'sd0.011703057539308764, 32'sd0.06669815036525888, 32'sd0.09605898685680574, 32'sd0.05265878651162231, 32'sd-0.01715836350043218, 32'sd0.11479991492887891, 32'sd0.06679229063014144, 32'sd-0.11937428683629227, 32'sd0.020789439112658355, 32'sd0.031191992133071996, 32'sd0.057355527245785146, 32'sd-0.031775841558852436, 32'sd0.018780200166168028, 32'sd-0.023498351756079897, 32'sd-0.0485781776925862, 32'sd0.05030030280734116, 32'sd-0.08454258917377497, 32'sd-0.052663489188347325, 32'sd-0.0833027627703676, 32'sd-0.13881572695195807, 32'sd-0.18451741439445465, 32'sd-0.31929269832194496, 32'sd-0.33028488067011924, 32'sd-0.19759254751930477, 32'sd-0.33673779404762466, 32'sd-0.2345066584667496, 32'sd-0.19448762529227853, 32'sd-0.021199312061458284, 32'sd0.07326944310347543, 32'sd0.06737805340541847, 32'sd0.07957111909633426, 32'sd0.031592860226283825, 32'sd-0.018681853835869178, 32'sd0.005385681419649193, 32'sd-0.06059448729354259, 32'sd0.05006939120110089, 32'sd-0.0191827207125258, 32'sd0.12930914881473818, 32'sd0.02054532492769744, 32'sd-0.026686096548765113, 32'sd-0.007572238353177308, 32'sd-0.02007835536462794, 32'sd-0.04866907125524147, 32'sd-0.03610146294220614, 32'sd-0.0951457741714398, 32'sd-0.14200663844559125, 32'sd-0.2237216930576775, 32'sd-0.31790340884295737, 32'sd-0.2602372089566173, 32'sd-0.3317184190934062, 32'sd-0.3618165591321085, 32'sd-0.4197199862334572, 32'sd-0.2817214526982706, 32'sd-0.18829937999346363, 32'sd-0.1583494539541713, 32'sd-0.042560236245581404, 32'sd-0.009115839744162663, 32'sd0.049206198475493505, 32'sd-0.056012015898144155, 32'sd-0.027024245430624576, 32'sd0.004150247716368077, 32'sd-0.03484887118421751, 32'sd-0.028234281624993616, 32'sd0.02756698014331892, 32'sd-0.014338550006521249, 32'sd-0.047103431171766706, 32'sd-0.05263979212169409, 32'sd0.04441601430352822, 32'sd-0.02612537055526742, 32'sd-0.10552062115020178, 32'sd-0.05446659673472694, 32'sd-0.1659006486100565, 32'sd-0.28457546282907953, 32'sd-0.21802816996314162, 32'sd-0.2578923725392069, 32'sd-0.26387508821205935, 32'sd-0.23736146739263445, 32'sd-0.15407406801048307, 32'sd-0.22632679300473255, 32'sd-0.13389793285552387, 32'sd-0.017195458774167057, 32'sd-0.07613113217085202, 32'sd0.05820936703982045, 32'sd-0.0865364642181756, 32'sd-0.0771316491741439, 32'sd-0.026607030902258785, 32'sd-0.05002451011037829, 32'sd0.00920839168284246, 32'sd0.021964422471937497, 32'sd-0.20342287266597622, 32'sd0.08302394664126411, 32'sd0.018127016510943467, 32'sd-0.009638161656638626, 32'sd-0.10564696391606797, 32'sd0.039311886515472565, 32'sd0.08313191828897623, 32'sd0.006008935594779465, 32'sd-0.007834755011440264, 32'sd-0.1255232518001431, 32'sd-0.11116922040859835, 32'sd-0.16824536287736294, 32'sd-0.29153268017090755, 32'sd-0.26328508260406497, 32'sd-0.1710215339010284, 32'sd-0.04738761043778143, 32'sd-0.11982706266314122, 32'sd-0.11411937257757354, 32'sd-0.03907868560393981, 32'sd0.20662801861347693, 32'sd0.047174131288593844, 32'sd0.01461756294092578, 32'sd-0.11615356796435951, 32'sd-0.16499444486207565, 32'sd-0.0074988601467626415, 32'sd-0.0025657627565203087, 32'sd-0.01984036835135488, 32'sd-0.05453278110871674, 32'sd-0.12678900291172485, 32'sd-0.04294953381432259, 32'sd0.005669579591503649, 32'sd-0.01813802687914171, 32'sd0.02738706670293283, 32'sd0.006079740860202347, 32'sd0.022673552465014346, 32'sd-0.006636465372434989, 32'sd-0.009821670999082618, 32'sd-0.08496141219524732, 32'sd-0.05021416816239332, 32'sd-0.0348617382511571, 32'sd0.07231013433967805, 32'sd-0.04565677388256194, 32'sd0.10750587851459363, 32'sd0.17927833766069246, 32'sd0.1426116312389201, 32'sd0.03513012495022495, 32'sd0.17371894776882962, 32'sd0.21707393405796266, 32'sd0.0193267660598604, 32'sd-0.0033187988465441056, 32'sd-0.11195609888837521, 32'sd-0.08241958704473351, 32'sd0.03271832508392695, 32'sd0.012199494579509676, 32'sd0.015461726550838115, 32'sd-0.015563820876020847, 32'sd0.04219094678183595, 32'sd-0.04430040670850827, 32'sd0.08786868221467642, 32'sd0.02462632862276575, 32'sd0.031576377947922896, 32'sd-0.0699479967375946, 32'sd-0.016047407717274906, 32'sd-0.09115607358503935, 32'sd-0.00784242989446106, 32'sd0.00031427636707235276, 32'sd-0.05501253844217224, 32'sd0.10386604663404742, 32'sd0.15769009953284538, 32'sd0.1869202362197939, 32'sd0.17223467865358122, 32'sd0.12140685325099654, 32'sd0.08128234036858553, 32'sd0.05402378440855882, 32'sd0.03010210803337153, 32'sd0.10001203704472353, 32'sd-0.031725448460489684, 32'sd-0.014971211908230652, 32'sd-0.040733381967378766, 32'sd0.06770130073861025, 32'sd0.02811289389481596, 32'sd-0.06793506815045232, 32'sd-0.015241400843118353, 32'sd-0.024610646866164054, 32'sd-0.06444799597114072, 32'sd0.11223670252673408, 32'sd0.042116738635469296, 32'sd-0.02885694441790689, 32'sd-0.04336114800222996, 32'sd0.10368885607140406, 32'sd0.056884045266837824, 32'sd-0.0188124039866827, 32'sd0.05703246794365584, 32'sd-0.03460853031281239, 32'sd0.07292678524324887, 32'sd0.14289191142073968, 32'sd0.1772179228375605, 32'sd0.187856666424142, 32'sd0.1697496349945929, 32'sd0.19051149213981033, 32'sd0.029328505006781854, 32'sd0.11156780336191752, 32'sd0.012969676362241094, 32'sd-0.014267206521700685, 32'sd-0.013416729458763483, 32'sd-0.03257212547795579, 32'sd0.01869940736964712, 32'sd-0.04001530631922758, 32'sd0.00427852665876092, 32'sd0.05316448216478306, 32'sd-0.03292720657760348, 32'sd-0.0427658108269174, 32'sd-0.03222585952773431, 32'sd-0.009594596616876564, 32'sd-0.05197860945228047, 32'sd-0.035325088637424756, 32'sd-0.04815518677241716, 32'sd0.16780784650694716, 32'sd-2.535940336800084e-119, 32'sd0.008373277156734981, 32'sd-0.01940991648197783, 32'sd-0.0014095552824313138, 32'sd0.013455793228592007, 32'sd0.14125897141954355, 32'sd0.20283747613704164, 32'sd0.09958561034406935, 32'sd0.043167091425173915, 32'sd-0.018799550605914483, 32'sd-0.1039523164771545, 32'sd-0.06134117883550855, 32'sd0.1460425067338198, 32'sd0.08928918726388406, 32'sd0.05508979876282236, 32'sd-0.002415509557292137, 32'sd-0.04839237195586229, 32'sd-0.04002748576538745, 32'sd-0.15178266414192398, 32'sd0.057839967023799954, 32'sd0.0070455239299542045, 32'sd-0.08262132534732086, 32'sd-0.07989635355549936, 32'sd0.04096443525491526, 32'sd0.09928518898464428, 32'sd-0.025409612847847124, 32'sd-0.011244158985014858, 32'sd-0.024944225678512198, 32'sd0.03208095385328928, 32'sd0.09901406381765537, 32'sd-0.005911173572392059, 32'sd0.12654741649444023, 32'sd0.03037625807207156, 32'sd0.1463819424838353, 32'sd0.07474551141825192, 32'sd0.011569440269470679, 32'sd-0.0964880093173456, 32'sd-0.09820345668645344, 32'sd-0.12866372790886452, 32'sd-0.056514127063504185, 32'sd0.10756606658379719, 32'sd0.13700042053757963, 32'sd-0.08649456956493962, 32'sd0.06863630413736535, 32'sd-0.06262806951304913, 32'sd0.0698739242524242, 32'sd-0.03674245962149959, 32'sd0.0685425034929752, 32'sd0.06125136767574741, 32'sd0.038187846961482634, 32'sd-0.05327381552862408, 32'sd0.12705611059793578, 32'sd0.0017971915661116878, 32'sd-0.11893973623593561, 32'sd0.01585716552100947, 32'sd-0.035132652483743046, 32'sd0.07712269010483469, 32'sd0.07612704723227598, 32'sd0.035385958893269835, 32'sd0.056660206171035676, 32'sd-0.05350789944813124, 32'sd0.06461288895081857, 32'sd-0.10984433713108695, 32'sd-0.0902360429795341, 32'sd-0.08709832412127312, 32'sd-0.07556358549759314, 32'sd-0.08304120799241889, 32'sd0.05800736257304952, 32'sd-0.007557355770110445, 32'sd0.12083148444894255, 32'sd-0.051898667839434184, 32'sd-0.08959477190452124, 32'sd0.07003546149133798, 32'sd0.04526053550481312, 32'sd0.018983997038019774, 32'sd0.08417875867015272, 32'sd0.10317916157131728, 32'sd-0.029911986268976867, 32'sd0.06432886189184117, 32'sd0.015082517889713803, 32'sd-0.05855733388200904, 32'sd0.13574425446156532, 32'sd0.09881161559336848, 32'sd0.04298323207647282, 32'sd-3.0839324418170685e-116, 32'sd0.005007701683355641, 32'sd0.07420766216643793, 32'sd-0.009720856854140765, 32'sd-0.059551110656386165, 32'sd0.001996159569371725, 32'sd0.05853510448069133, 32'sd0.006238671042400501, 32'sd0.007062186297173896, 32'sd-0.12079032189331172, 32'sd0.08796147936234096, 32'sd-0.019933487610125766, 32'sd0.022625046600819546, 32'sd-0.07036569631655497, 32'sd-0.010051063879981992, 32'sd0.056673285827631543, 32'sd-0.02402620417864574, 32'sd0.019242081181906175, 32'sd0.08024601779081628, 32'sd-0.0430003403712295, 32'sd0.04316681080104417, 32'sd-0.02060770396039285, 32'sd0.03053968905206323, 32'sd0.045180580101917944, 32'sd0.034970308427406595, 32'sd0.05473787224980777, 32'sd0.09141427619514197, 32'sd0.014123206249356675, 32'sd0.0022843055850172377, 32'sd0.02095998867073778, 32'sd0.09699008301982345, 32'sd0.019474952628298424, 32'sd0.010285772127669821, 32'sd-0.01928290787482762, 32'sd0.006355831794556273, 32'sd-0.01751610200177405, 32'sd0.01333816702576153, 32'sd-0.08254769195112267, 32'sd0.007129948301823307, 32'sd-0.10206730937920382, 32'sd0.07274956936395312, 32'sd0.06390847641626281, 32'sd0.10534380648373005, 32'sd0.029509461738898655, 32'sd-0.05405195062402922, 32'sd-0.03634257909965154, 32'sd0.008897849879799101, 32'sd0.15639930976956073, 32'sd-0.01931765023789609, 32'sd0.09952146847309752, 32'sd0.006021938303235742, 32'sd0.005869986967869506, 32'sd0.05452463520702028, 32'sd0.12983877141712297, 32'sd0.006674392496652649, 32'sd0.0019570496613516477, 32'sd-0.05147036380906223, 32'sd0.034159218822862415, 32'sd0.12023199754807944, 32'sd0.0703857910307328, 32'sd0.027638828261134916, 32'sd0.09506263828286758, 32'sd0.048689915687000505, 32'sd0.0007648503128768191, 32'sd0.061090529416343235, 32'sd-0.012545096488165772, 32'sd-0.029387133784178877, 32'sd0.0019650160674263683, 32'sd-0.032308832532667836, 32'sd0.016827350467313717, 32'sd-0.11469922007648584, 32'sd-0.08206137232875678, 32'sd-0.011727100704455902, 32'sd0.06659406447147656, 32'sd0.023700673959757307, 32'sd-0.04351992854342005, 32'sd0.06426820327401082, 32'sd0.007479813358552741, 32'sd-0.1463024456811188, 32'sd-0.06970051475364752, 32'sd0.010843676309867996, 32'sd0.01982775101319239, 32'sd0.07658117358311484, 32'sd0.09442290008833301, 32'sd-6.811644853493241e-126, 32'sd0.06286272895869661, 32'sd-0.014280863764077983, 32'sd0.029729725893687962, 32'sd0.0063281601329632795, 32'sd0.03279095466285376, 32'sd-0.059717453170152736, 32'sd0.09325241892906924, 32'sd0.036177679520745076, 32'sd-0.0006226622539417404, 32'sd-0.039631050697493564, 32'sd-4.7789191066189264e-05, 32'sd-0.06924498581809481, 32'sd-0.012209342607210452, 32'sd-0.02989268466045924, 32'sd-0.07133486890858574, 32'sd-0.11561421466468753, 32'sd-0.18336756208785854, 32'sd-0.1252245772066194, 32'sd-0.07883711726724478, 32'sd-0.037498417161087726, 32'sd0.018615869480767593, 32'sd-0.05414591578082389, 32'sd-0.0397173251748005, 32'sd0.031160522973326183, 32'sd0.07912206368310568, 32'sd-0.023217062520545437, 32'sd-2.3446924399362935e-116, 32'sd-9.133818785196426e-124, 32'sd-1.0533090823230917e-124, 32'sd-0.0891830843406005, 32'sd0.020173296683659116, 32'sd0.04138274473537182, 32'sd0.018226733460349167, 32'sd-0.061459323354191416, 32'sd0.022867397575554234, 32'sd0.15343814703187192, 32'sd0.06125996295524795, 32'sd0.055259232680010414, 32'sd0.12074553738176355, 32'sd0.04641815505605698, 32'sd-0.025039125736139024, 32'sd0.1525628594325409, 32'sd-0.05677539160165878, 32'sd-0.12087973404796329, 32'sd-0.047933701876013535, 32'sd-0.024431307421440382, 32'sd0.03498858186897032, 32'sd-0.021536972994224232, 32'sd0.0036312551558599013, 32'sd0.10241245630801071, 32'sd-0.03671142648329521, 32'sd0.08048283216294541, 32'sd0.015009998270185714, 32'sd-0.00492996036448244, 32'sd-1.5010659162555626e-125, 32'sd1.0468217864848844e-124, 32'sd-4.699507417086011e-124, 32'sd0.02531048276308599, 32'sd0.06781067989984421, 32'sd0.012679955991806543, 32'sd-0.04300396620528817, 32'sd0.058617902117449286, 32'sd0.030061939368013504, 32'sd-0.014969267434207602, 32'sd-0.02249736963066504, 32'sd0.05670713117875818, 32'sd-0.008400393246124061, 32'sd0.12693259420856642, 32'sd-0.09754978828855214, 32'sd0.030667754383559998, 32'sd0.10539545074254841, 32'sd-0.10709740809693122, 32'sd0.04871965899322492, 32'sd-0.18151921075809324, 32'sd-0.06994070308615356, 32'sd-0.0736453479003233, 32'sd0.014610182844981492, 32'sd0.04070129119806146, 32'sd0.0021410531524356817, 32'sd-0.08672466552452177, 32'sd0.04827361977521473, 32'sd0.0372669118821532, 32'sd-1.7379657260496208e-125, 32'sd-2.149138119575137e-116, 32'sd1.2145745112176135e-120, 32'sd-1.7117373312281265e-127, 32'sd0.06620637119408297, 32'sd0.0013269569258849386, 32'sd0.03759655055595706, 32'sd-0.013927241353864877, 32'sd-0.06557394043118404, 32'sd-0.06122207718163858, 32'sd0.028770180111301256, 32'sd0.08518873204505752, 32'sd0.1147152542679812, 32'sd0.02526579954382609, 32'sd0.06347581944825159, 32'sd0.055610715312037665, 32'sd-0.047581329873774614, 32'sd0.04609152599032645, 32'sd-0.0065330198196078, 32'sd0.11329454623569817, 32'sd-0.009923598746820188, 32'sd-0.009589207304428013, 32'sd-0.08034881745792682, 32'sd-0.03390838999675115, 32'sd0.10664922537780155, 32'sd-0.011245762328317074, 32'sd0.1229214353343739, 32'sd6.180570941167006e-122, 32'sd1.1515291174337733e-122, 32'sd-5.674095168741158e-124, 32'sd-6.167538619296633e-126, 32'sd-3.180040260692619e-120, 32'sd6.741345811916526e-120, 32'sd0.1452569453292282, 32'sd0.03904145903773453, 32'sd0.10941596910341786, 32'sd0.09288038115472325, 32'sd0.14828372040204307, 32'sd0.06122411593884774, 32'sd0.03253241645327648, 32'sd0.10761027745466298, 32'sd0.1772461889052077, 32'sd0.10918510903974872, 32'sd0.08093677225847956, 32'sd0.1233176214527298, 32'sd0.0632848486168273, 32'sd0.05855702826792357, 32'sd0.029247094936431874, 32'sd-0.026697261201339594, 32'sd0.04586763528685485, 32'sd0.0313181873941732, 32'sd-0.05630902848002758, 32'sd0.16531895576741257, 32'sd3.4224007640726203e-124, 32'sd-2.084476039565583e-117, 32'sd-1.2338057876477506e-118, 32'sd1.6778065951300006e-124},
        '{32'sd2.7203193200622043e-121, 32'sd1.7760670830993558e-124, 32'sd1.7031752603658355e-125, 32'sd-4.20215268266087e-118, 32'sd1.6724865010893093e-123, 32'sd2.1164762427753106e-117, 32'sd-4.871879862691078e-123, 32'sd-5.670040465329354e-115, 32'sd4.23562926311185e-125, 32'sd2.8337708273048686e-120, 32'sd-2.0456273902435625e-117, 32'sd-1.9392043932926444e-127, 32'sd0.03725511070992748, 32'sd-0.041224758803930214, 32'sd0.01655726032070195, 32'sd-0.036559052236487005, 32'sd1.6148290542086118e-125, 32'sd2.5359114400859135e-114, 32'sd1.0766972941290774e-115, 32'sd2.499414134541422e-126, 32'sd5.231682548484362e-123, 32'sd-2.116518305524964e-117, 32'sd-6.922155259480574e-124, 32'sd-4.288969309460744e-121, 32'sd-4.869890398357605e-123, 32'sd-2.5201645529588797e-117, 32'sd1.2144522957399582e-122, 32'sd1.9956005945663752e-120, 32'sd-9.049868619082261e-121, 32'sd-3.7022892340518877e-122, 32'sd-3.189400130730237e-120, 32'sd-1.0692610698939833e-121, 32'sd-0.018119680093324216, 32'sd0.04730723720452995, 32'sd0.002196557683993877, 32'sd0.0008127789885522116, 32'sd0.055988180492472665, 32'sd0.09734431300743504, 32'sd0.0434915027013099, 32'sd0.09900214808092882, 32'sd0.06787711194483335, 32'sd-0.05292222493499177, 32'sd-0.012613063233608151, 32'sd0.024553977356923787, 32'sd0.07781132656920121, 32'sd-0.03453625200534552, 32'sd0.04645119348129703, 32'sd0.04788831237994902, 32'sd0.028395895315710115, 32'sd-0.006576486639799591, 32'sd0.03812398786058374, 32'sd-0.0073262570646366685, 32'sd4.898907803765875e-124, 32'sd-2.486356724507068e-123, 32'sd2.0447695981561277e-127, 32'sd-1.6249930438384443e-115, 32'sd2.8678029318681185e-128, 32'sd-2.1518954145872025e-126, 32'sd0.056778928310836314, 32'sd-0.04221950979357201, 32'sd-0.07917897991858484, 32'sd-0.044510951630107466, 32'sd0.09000279487711561, 32'sd0.024965062979986984, 32'sd0.011156556780273833, 32'sd-0.02009733647181441, 32'sd-0.007267103576670621, 32'sd0.010605543725451878, 32'sd0.11823713186697533, 32'sd0.09153810601962692, 32'sd0.08391300502465929, 32'sd0.07472760633852726, 32'sd0.06750093832781606, 32'sd-0.04211165521456264, 32'sd-0.03006216631929911, 32'sd0.021229521004006324, 32'sd0.04879696756712068, 32'sd-0.03477254399153985, 32'sd-0.07074241071736528, 32'sd0.08489955331388363, 32'sd-0.027121546707612236, 32'sd0.0216898075516093, 32'sd1.6504089604961308e-123, 32'sd-1.875381381846591e-129, 32'sd-7.740772079428661e-125, 32'sd1.461367862471763e-126, 32'sd-0.04227647355461197, 32'sd0.02131740751397237, 32'sd0.014477523904915031, 32'sd0.039397949706378374, 32'sd-0.006067871844444399, 32'sd-0.09680632424020577, 32'sd-0.13290918154031472, 32'sd0.08498321834417115, 32'sd0.0292573509441313, 32'sd-0.023886821474641003, 32'sd0.08977228928699033, 32'sd0.018740531371270932, 32'sd0.0034776413460569874, 32'sd0.0450424743566902, 32'sd0.20689344340222693, 32'sd0.06211934870564649, 32'sd0.0697212895599276, 32'sd0.015121003619761708, 32'sd-0.012983390228831368, 32'sd-0.015494206717699034, 32'sd-0.012598839826582966, 32'sd-0.08526623232024147, 32'sd-0.05543409230003524, 32'sd0.06727294050809982, 32'sd0.11867438457437054, 32'sd3.338349125847422e-121, 32'sd-2.1309858102532348e-126, 32'sd-0.004938154281902406, 32'sd0.037698954677085, 32'sd-0.0677289615773344, 32'sd0.03704423855485997, 32'sd-0.023448410541060824, 32'sd-0.12040583830338658, 32'sd-0.05647727981534438, 32'sd-0.08811294089804803, 32'sd-0.08435278228940629, 32'sd-0.19998524557953262, 32'sd-0.16520029962392002, 32'sd-0.029048504001818142, 32'sd-0.06910562713726182, 32'sd-0.006228888238791824, 32'sd0.07084250328822721, 32'sd0.07490201693910678, 32'sd-0.06813463240703085, 32'sd0.044640149336087794, 32'sd0.046243869845171856, 32'sd-0.06419664815830621, 32'sd-0.07605515095801549, 32'sd-0.07626554776536514, 32'sd-0.042355698034323847, 32'sd-0.014500627662243807, 32'sd-0.007685252440764933, 32'sd-0.056731580770855876, 32'sd0.004981597133476551, 32'sd1.294003762198183e-125, 32'sd0.03144443423762249, 32'sd-0.023293344753905657, 32'sd-0.04749897902853855, 32'sd0.03874948594649611, 32'sd-0.1481221599964417, 32'sd-0.08650018819357305, 32'sd-0.158040172372474, 32'sd-0.07070120870612219, 32'sd-0.0021852026232921976, 32'sd-0.07593595149124797, 32'sd-0.0621491463643934, 32'sd-0.15633652857801342, 32'sd0.06785716457086426, 32'sd0.10024505678232364, 32'sd-0.015916628373165556, 32'sd0.0008798567432108834, 32'sd-0.03762199997046848, 32'sd0.04393449626670541, 32'sd0.001297547608017481, 32'sd-0.15067679464317377, 32'sd-0.004003464617726642, 32'sd0.007652893831374029, 32'sd-0.04297565059701648, 32'sd0.0011210335524740932, 32'sd-0.004451724302179653, 32'sd0.03946495604790299, 32'sd0.03737941392123711, 32'sd7.065499236138096e-115, 32'sd0.02709667070684926, 32'sd0.046864679980703955, 32'sd-0.09270232584110119, 32'sd-0.013267021889612436, 32'sd0.06489776608624255, 32'sd0.04382099797685055, 32'sd-0.08455462080379315, 32'sd-0.16738092501460383, 32'sd-0.056945677285203035, 32'sd0.013324063252420639, 32'sd-0.16303735437130076, 32'sd-0.1704391440734967, 32'sd-0.02486349612289675, 32'sd-0.09953943248921572, 32'sd-0.07427421107896873, 32'sd-0.044724120378457834, 32'sd0.10878410006908358, 32'sd0.008208867521331962, 32'sd0.08350977859810552, 32'sd0.05601484194146503, 32'sd0.04353683997297933, 32'sd0.07043000342867752, 32'sd-0.012686139387785626, 32'sd0.05066134619341376, 32'sd-0.11315867976357645, 32'sd0.014357386366088475, 32'sd0.03036378121969056, 32'sd0.06971884932240897, 32'sd-0.013648812084398337, 32'sd-0.02436434218038157, 32'sd-0.0644620022990403, 32'sd-0.06110073720263891, 32'sd0.06308306502391559, 32'sd0.06295618059116778, 32'sd-0.010148207970682534, 32'sd-0.13099002861259648, 32'sd-0.05851124768194239, 32'sd-0.07519544260339946, 32'sd-0.11409730174212893, 32'sd-0.061071199624309395, 32'sd-0.004142708906534414, 32'sd0.02046816681201026, 32'sd0.03900947306019873, 32'sd0.06692608131494847, 32'sd0.04100667660417718, 32'sd0.15338080877086563, 32'sd0.022543032479906043, 32'sd0.1358752341398199, 32'sd-0.0395603917158174, 32'sd0.017520532507805206, 32'sd0.059396088770220686, 32'sd0.005763350461701616, 32'sd-0.12810644423515682, 32'sd0.08201453091492747, 32'sd-0.06623854821054943, 32'sd0.04608239845529834, 32'sd0.06946605889586109, 32'sd0.013082845377145194, 32'sd0.019778389873643172, 32'sd0.012251978215465649, 32'sd0.0337739538240603, 32'sd0.026873850615893383, 32'sd-0.0514735675782691, 32'sd-0.16951322197297444, 32'sd-0.11752375372468309, 32'sd-0.0919585055233746, 32'sd0.047580257368703215, 32'sd0.021209299695861716, 32'sd-0.059224418318936135, 32'sd0.10441268206947021, 32'sd0.054114172956552666, 32'sd0.1309271208292541, 32'sd0.11696081749964297, 32'sd0.14322318019228722, 32'sd0.18484624567640406, 32'sd0.2032572733897184, 32'sd0.11403142681616608, 32'sd0.1822469231334259, 32'sd0.14457137295517727, 32'sd-0.10519773010799917, 32'sd0.001715724799823218, 32'sd0.022370767730213088, 32'sd0.0843202119772354, 32'sd-0.01465222795681911, 32'sd-0.09306202086119608, 32'sd0.026386633256185236, 32'sd0.01790142764250628, 32'sd-0.05595394741519874, 32'sd-0.05274202358433773, 32'sd0.012400351895118905, 32'sd0.021600615617400724, 32'sd-0.04333004305351249, 32'sd-0.007849951852210978, 32'sd-0.0775330159948153, 32'sd-0.03663352291847478, 32'sd0.20148406439533698, 32'sd0.015080946144854123, 32'sd0.04754508712033846, 32'sd0.12752934434362367, 32'sd0.037898124313879435, 32'sd0.09589695982205346, 32'sd0.131646543297877, 32'sd0.028726651461063256, 32'sd0.16059221916756786, 32'sd0.1639609938874005, 32'sd0.07381628508030193, 32'sd0.1041052575737486, 32'sd0.006882543655712343, 32'sd0.044503411639865306, 32'sd-0.052305351506414285, 32'sd-0.006752896536972345, 32'sd0.018499986741162558, 32'sd-0.07883377844066534, 32'sd-0.007689474651119074, 32'sd-0.12802846717117183, 32'sd0.014437727253494266, 32'sd-0.06614708910788089, 32'sd-0.08335050429990114, 32'sd-0.07665929365205064, 32'sd-0.020924729699430104, 32'sd-0.029920730841760466, 32'sd0.06762342674722607, 32'sd-0.03001267012943784, 32'sd0.04402582155970883, 32'sd0.08596950462494202, 32'sd0.12671177312320225, 32'sd0.037588660422115755, 32'sd0.14806084418854523, 32'sd0.003239987313777795, 32'sd0.07859322352915547, 32'sd-0.03090880670950759, 32'sd0.04358583146890677, 32'sd0.09077232056155525, 32'sd0.07990710807540555, 32'sd0.036962272430654274, 32'sd0.05141664603368261, 32'sd0.02454402583089781, 32'sd0.08975886304326224, 32'sd0.04970134888619216, 32'sd0.062259201628825686, 32'sd0.11644334441529838, 32'sd-0.028227370931893273, 32'sd-0.06791137848770573, 32'sd-0.09081083620057911, 32'sd-0.12194966371059039, 32'sd-0.00032677155042984304, 32'sd0.007913939845518593, 32'sd-0.031110454976556637, 32'sd0.020420047503790114, 32'sd0.026449102425049168, 32'sd0.04703127513496473, 32'sd-0.11650185027141279, 32'sd-0.004962616133548869, 32'sd0.027660400669204287, 32'sd0.09991187018846522, 32'sd-0.02579207039222797, 32'sd-0.08780889527693543, 32'sd-0.057469291759107, 32'sd0.06320275227417008, 32'sd0.07723107324358389, 32'sd-0.06228574711196731, 32'sd-0.051074906238649236, 32'sd0.0018118205916746748, 32'sd0.13144816785735994, 32'sd-0.013539696948244771, 32'sd-0.012854953243206117, 32'sd0.058327004990408896, 32'sd0.07665295621788752, 32'sd-0.03133334414309997, 32'sd0.018210567630163054, 32'sd0.0758537491490093, 32'sd-0.13954647344193225, 32'sd-0.11720629072665639, 32'sd0.007813897130656926, 32'sd-0.06569804867929564, 32'sd-0.1052253135988808, 32'sd-0.014911083305951802, 32'sd0.014465499045697269, 32'sd-0.026486582160198207, 32'sd-0.10673403056804863, 32'sd0.020930282550515565, 32'sd0.06664504086963263, 32'sd0.014764790006906926, 32'sd0.05226254984063395, 32'sd-0.033012649391104806, 32'sd0.12046610882665815, 32'sd-0.010218827236616816, 32'sd-0.07689494908916496, 32'sd0.01958611804358384, 32'sd0.10616500461579481, 32'sd0.08631764226674317, 32'sd-0.0023958410387738085, 32'sd0.029631360061472132, 32'sd-0.05445770579481221, 32'sd0.0850776008614873, 32'sd0.0238178104862602, 32'sd0.09169899494629068, 32'sd0.04453142349985219, 32'sd0.07527273274298853, 32'sd-0.06520456516782457, 32'sd-0.09276993348873515, 32'sd0.0669149032782853, 32'sd0.018175764840312632, 32'sd-0.0058487748996740455, 32'sd-0.013629008719168311, 32'sd0.095404954805602, 32'sd0.026115971453250904, 32'sd0.05952173200558897, 32'sd0.09030484996348678, 32'sd0.08304786542333757, 32'sd-0.022771524832564508, 32'sd-0.07874207867315428, 32'sd-0.018068314724127076, 32'sd-0.10867626179885946, 32'sd-0.10001167567488374, 32'sd-0.04438119953993422, 32'sd0.03539848876009003, 32'sd0.07455156701621714, 32'sd0.03960793687874029, 32'sd9.103859995578254e-06, 32'sd-0.028693213940025216, 32'sd-0.06316264273521727, 32'sd0.09754772402211163, 32'sd0.028425979567537615, 32'sd0.04502038249172956, 32'sd-0.005406639887784578, 32'sd0.03604495363519927, 32'sd-0.04383234804013815, 32'sd0.1741693854312536, 32'sd0.024637738770045218, 32'sd-0.0862837694775237, 32'sd-0.04592071759315774, 32'sd0.05594094497469166, 32'sd0.08360107752866854, 32'sd0.14449624883427298, 32'sd0.021834589596655306, 32'sd0.06253440389323599, 32'sd-0.057578412686843806, 32'sd-0.05843744096540922, 32'sd-0.15680541915886695, 32'sd0.03189409379750299, 32'sd-0.06555365199056726, 32'sd-0.07186979311193718, 32'sd0.004237013640981143, 32'sd0.042759637685628266, 32'sd-0.05970177827314678, 32'sd0.05742611938978986, 32'sd0.07193807024022815, 32'sd-0.09670217876337017, 32'sd-0.07349368599329378, 32'sd-0.013283892314720908, 32'sd-0.01723709214262414, 32'sd0.011021195102601076, 32'sd-0.10576053027137913, 32'sd-0.1461493969187878, 32'sd0.03753739250247953, 32'sd0.2126170704231297, 32'sd0.10621632632152951, 32'sd-0.0202428735814925, 32'sd0.006194867218677349, 32'sd-0.020507758839563784, 32'sd0.1027488919664642, 32'sd0.09965911738844356, 32'sd0.010302523201047431, 32'sd-0.1419229056937219, 32'sd-0.2320486785357557, 32'sd-0.007652221273752737, 32'sd-0.08843122803060575, 32'sd-0.03148961031350175, 32'sd0.08685933147316316, 32'sd-0.009942425242203587, 32'sd-0.037976018771292454, 32'sd-0.035046304867795586, 32'sd0.04310496047676538, 32'sd-0.00048460858069884636, 32'sd0.17533044808256174, 32'sd0.013153198773310275, 32'sd-0.026703695170484713, 32'sd-0.017955670349369346, 32'sd0.023973155478543604, 32'sd0.04372511492344673, 32'sd0.004944826948499794, 32'sd-0.09158416967297345, 32'sd-0.005662014717492641, 32'sd0.10052734355406812, 32'sd0.028576991174832013, 32'sd-0.08181661567517755, 32'sd-0.02976176703141577, 32'sd-0.03207844853853933, 32'sd0.05336394719083076, 32'sd0.08924989088595679, 32'sd-0.050790522233231404, 32'sd-0.27795917331409514, 32'sd-0.1534493121106674, 32'sd-0.022642929353793508, 32'sd0.022095323276258603, 32'sd-0.008997168281057571, 32'sd0.018370933437936113, 32'sd-0.05399205490885282, 32'sd0.02780819735747473, 32'sd-0.03232005804077436, 32'sd0.049226838415821234, 32'sd-0.0807283067135108, 32'sd-0.022385739480568188, 32'sd0.10340712739663374, 32'sd0.09420359408993266, 32'sd0.04865931962949981, 32'sd-1.6802230184272158e-124, 32'sd-0.03645771026893751, 32'sd-0.03418008519602534, 32'sd-0.00026345172165363436, 32'sd-0.0006074325318233826, 32'sd-0.005789700596893442, 32'sd0.07718960232074147, 32'sd0.10626657014329706, 32'sd-0.007296557473414641, 32'sd0.10026193188413897, 32'sd0.04907275915925615, 32'sd-0.07558068957614605, 32'sd-0.05034144307253937, 32'sd-0.1189402995164515, 32'sd-0.09046556744801573, 32'sd-0.05935337286761663, 32'sd0.10028748321121764, 32'sd-0.001720668426929609, 32'sd-0.017403524518678225, 32'sd0.030959175507129007, 32'sd0.007243625111332168, 32'sd-0.0762920861763547, 32'sd-0.12315263486191141, 32'sd0.03331601149330116, 32'sd0.026829066978719743, 32'sd0.007041331230672923, 32'sd-0.009176004785560665, 32'sd0.047929827309090636, 32'sd-0.04582944511918873, 32'sd0.03524033231863689, 32'sd-0.03003052826135033, 32'sd-0.13628137221429762, 32'sd0.04610391060625424, 32'sd0.029287046862328168, 32'sd0.03692736710679844, 32'sd-0.03944151719103321, 32'sd0.10004446670561258, 32'sd0.14378208157614492, 32'sd0.07611175705808178, 32'sd-0.1094497100431037, 32'sd-0.18651313743104986, 32'sd-0.18623617128260037, 32'sd-0.027490368080945488, 32'sd0.10493528806456529, 32'sd-0.018856277617113403, 32'sd0.003047997199044535, 32'sd-0.12066270676783969, 32'sd-0.11780441703601724, 32'sd0.03116659362275707, 32'sd-0.0919804573399642, 32'sd-0.014374701799871019, 32'sd-0.08120377646770818, 32'sd0.06258350238803187, 32'sd-0.03535854306216218, 32'sd-0.04011144651157693, 32'sd0.047233396250050505, 32'sd0.09512829467247952, 32'sd0.05955369994571861, 32'sd0.014692798503782611, 32'sd-0.1456098781135377, 32'sd-0.0887552933340708, 32'sd0.06981298935971174, 32'sd0.013733370886308873, 32'sd0.09716230357961568, 32'sd0.1604164176668683, 32'sd0.015930655980064847, 32'sd0.1190154071984073, 32'sd-0.038986645920038476, 32'sd0.005380009985957397, 32'sd-0.08892986139673144, 32'sd-0.042123586085266944, 32'sd-0.04999616074987116, 32'sd-0.07539448589678621, 32'sd-0.05184985609915949, 32'sd-0.09040794461397005, 32'sd-0.11440613965208095, 32'sd0.01455232867182713, 32'sd0.030438446777233605, 32'sd0.0333285505241923, 32'sd0.029778427714662818, 32'sd0.02997335046701423, 32'sd0.06334215307171123, 32'sd0.03412700014789502, 32'sd-0.052842762464107525, 32'sd-8.003720578421207e-122, 32'sd0.07859530785598108, 32'sd-0.05732943367542639, 32'sd-0.043255744887655, 32'sd-0.04056904023505912, 32'sd0.051734708865567164, 32'sd-0.10684789272224728, 32'sd-0.08092244585935497, 32'sd0.00023047402985528785, 32'sd-0.005723601695202561, 32'sd0.0757751350825178, 32'sd0.006163219622214233, 32'sd0.04143485440131133, 32'sd-0.038507938204648345, 32'sd-0.10124044918925187, 32'sd-0.015249339431564144, 32'sd-0.06377148788938992, 32'sd0.040846862052900786, 32'sd-0.021461037112971922, 32'sd0.003948778766490037, 32'sd-0.009988472325820131, 32'sd0.09418583488471174, 32'sd-0.005256084931906864, 32'sd0.009568959402932328, 32'sd-0.06497692065645119, 32'sd-0.04441558441561691, 32'sd-0.05602133958569692, 32'sd0.11980991313278574, 32'sd0.030021978637911628, 32'sd-0.10505701308457237, 32'sd-0.01002808947974197, 32'sd-0.048766803325161735, 32'sd0.047009798030532894, 32'sd-0.01668038389250189, 32'sd0.023279327977699875, 32'sd-0.05212706505092888, 32'sd0.029902440427810904, 32'sd-0.007101520738313542, 32'sd0.07634576427831875, 32'sd0.051807565423754705, 32'sd-0.06134251980737829, 32'sd-0.0593879961799336, 32'sd0.0006143118519634644, 32'sd-0.005359908491401678, 32'sd-0.0019076022868135785, 32'sd-0.11702745398380171, 32'sd-0.03828177093592301, 32'sd-0.07577970613771563, 32'sd-0.09290802099300008, 32'sd-0.05324360065065261, 32'sd-0.02278822224640222, 32'sd0.038662078595041095, 32'sd-0.19019472061888604, 32'sd-0.17574838086539088, 32'sd-0.05463133019338848, 32'sd0.019105730261676706, 32'sd-0.03314500456472043, 32'sd-0.06010540396496553, 32'sd-0.0817147425750565, 32'sd0.0424457028186186, 32'sd-0.11728995850703905, 32'sd-0.07961566063488068, 32'sd0.16212340344553944, 32'sd0.060528649552451026, 32'sd0.05609259522032052, 32'sd-0.02209748087894162, 32'sd-0.025804558868044274, 32'sd-0.004622871980951635, 32'sd0.04484938213419195, 32'sd0.031133086609661256, 32'sd0.066750307199594, 32'sd0.06435758502589986, 32'sd-0.042561159475853164, 32'sd-0.07027729765597898, 32'sd0.07973168045535461, 32'sd0.0015006873220662956, 32'sd-0.03976195001050814, 32'sd-0.05357687705443592, 32'sd-0.12050789956954856, 32'sd-0.012126768016286555, 32'sd-0.07757012963848532, 32'sd-0.07583963291657697, 32'sd-0.04957248893735235, 32'sd0.0660514096040957, 32'sd-1.7582128553065455e-123, 32'sd-0.004049765813192201, 32'sd-0.058382201974428685, 32'sd-0.07048745724609802, 32'sd-0.04882508241626123, 32'sd-0.09935115222347835, 32'sd-0.027920857375229025, 32'sd0.06848132587188531, 32'sd-0.07734471500914755, 32'sd0.09114027692378716, 32'sd0.07530065222261864, 32'sd0.09615935903727513, 32'sd0.13864432990984918, 32'sd0.11196646128447896, 32'sd0.08545232474153713, 32'sd0.11846494780583225, 32'sd-0.043129402562885596, 32'sd0.10205178508003612, 32'sd-0.03443139604276427, 32'sd0.006268217392653861, 32'sd-0.0997718261803835, 32'sd-0.08642796147710471, 32'sd-0.06092081162177616, 32'sd0.030324284497895978, 32'sd0.08902584798290006, 32'sd-0.009054997649842259, 32'sd-0.03736736126977306, 32'sd-9.199749827859479e-125, 32'sd6.150219167775755e-116, 32'sd-5.219914907943343e-118, 32'sd0.006516909388524126, 32'sd0.011655425296761914, 32'sd-0.14756612650272688, 32'sd-0.10172651779235141, 32'sd0.051085059050875216, 32'sd-0.014329965853958085, 32'sd0.10441181653848891, 32'sd0.0029542260668428792, 32'sd0.07184455223059694, 32'sd0.14788061844842434, 32'sd0.33875822596746114, 32'sd0.07478100689895886, 32'sd0.10716166608203723, 32'sd0.07793425760322382, 32'sd-0.08375524710357644, 32'sd0.0936467940712974, 32'sd-0.06646384441291314, 32'sd0.03732088442492955, 32'sd0.08631311727887198, 32'sd0.023300482011156656, 32'sd-0.019676403492991174, 32'sd0.0247810810921679, 32'sd0.010888883364928072, 32'sd-0.06653989414626627, 32'sd0.05801883570634664, 32'sd4.2824377653246305e-120, 32'sd2.816940793173307e-116, 32'sd1.0499701742366077e-119, 32'sd0.04907612829090982, 32'sd0.060414054530950535, 32'sd0.045483190384252234, 32'sd-0.10053214242479154, 32'sd0.08188346263051843, 32'sd-0.07641115936904858, 32'sd-0.0890516510366693, 32'sd0.07377401954241683, 32'sd0.0234388319659917, 32'sd0.019720610250191863, 32'sd0.004814292372994208, 32'sd-0.07237902555037615, 32'sd-0.04730085626738428, 32'sd-0.06020207397954095, 32'sd-0.03978329672360896, 32'sd0.037993821720277696, 32'sd0.07300290648486941, 32'sd0.02658877558024434, 32'sd0.04500981897406448, 32'sd-0.043079674207401476, 32'sd-0.025876998678460772, 32'sd-0.06754438939584805, 32'sd0.010915505246354897, 32'sd0.004503326208192699, 32'sd0.024719304798574357, 32'sd1.3929778537020316e-117, 32'sd3.394176329760563e-120, 32'sd5.271946363735653e-118, 32'sd2.285954624035455e-120, 32'sd0.039419912380847834, 32'sd-0.10789785943982466, 32'sd0.048195602079328936, 32'sd-0.01954787895809854, 32'sd0.009181854851278634, 32'sd-0.07129164120798556, 32'sd-0.10934535746572571, 32'sd-0.009456929711943677, 32'sd-0.05731900263911434, 32'sd-0.02974832953202418, 32'sd-0.06976016009091758, 32'sd0.007967514879389601, 32'sd-0.030535991603098354, 32'sd-0.04440880161069435, 32'sd-0.00012415627755965725, 32'sd-0.03567410858821531, 32'sd0.026168748204246955, 32'sd0.020815948362238355, 32'sd0.06466719675565281, 32'sd0.08955749497728395, 32'sd0.07469464596358917, 32'sd-0.09425151997684678, 32'sd-0.015094416565581373, 32'sd-3.719527746710294e-122, 32'sd-1.3201969583150432e-122, 32'sd-3.5599854880396364e-126, 32'sd2.0527753587847513e-125, 32'sd2.863047691367077e-115, 32'sd2.9308786883976844e-127, 32'sd0.03649038044888768, 32'sd0.079713317353257, 32'sd0.006956477615783233, 32'sd0.014356885917220655, 32'sd-0.05388106982662673, 32'sd-0.020635165317889923, 32'sd0.07841077663849089, 32'sd0.017208956991423816, 32'sd0.016263625507577952, 32'sd0.12755043895924062, 32'sd0.09026348177817067, 32'sd0.025678338366781288, 32'sd-0.0795654560037978, 32'sd-0.016097988561790247, 32'sd-0.025562315861513172, 32'sd0.05623337994911092, 32'sd0.11555488960887482, 32'sd0.10739098679496913, 32'sd-0.01544094342030417, 32'sd0.030838854640660197, 32'sd5.5010860002712683e-129, 32'sd1.2050053356533887e-118, 32'sd-6.824812915190904e-124, 32'sd-1.0360087711170701e-120},
        '{32'sd-3.044857682492247e-122, 32'sd7.72196671716271e-121, 32'sd4.846856105075303e-123, 32'sd1.0212962333041857e-115, 32'sd-4.699111525204252e-123, 32'sd3.322031568747786e-121, 32'sd-8.489067386094868e-122, 32'sd-4.088067768056438e-125, 32'sd7.3256818177687845e-127, 32'sd-2.148576391500656e-126, 32'sd5.766861426192338e-125, 32'sd3.934745522776016e-119, 32'sd0.07199549339263406, 32'sd0.05870486424372548, 32'sd-0.041203608073295955, 32'sd-0.008423286921895791, 32'sd3.495202316132521e-125, 32'sd1.7767776660868935e-123, 32'sd1.3545419366652716e-126, 32'sd6.781931198545949e-124, 32'sd3.065485321059541e-122, 32'sd-6.329947278906752e-115, 32'sd3.3587282075674525e-121, 32'sd-4.993293381994596e-126, 32'sd-5.170219104514477e-115, 32'sd9.478613428617495e-121, 32'sd1.8800089509270512e-127, 32'sd1.3875706680587251e-123, 32'sd-3.126294392589585e-114, 32'sd-2.0984076333173834e-117, 32'sd1.3672195839943939e-120, 32'sd5.504226835785763e-117, 32'sd0.05100557757686656, 32'sd0.03364514357138432, 32'sd-0.016442701184569614, 32'sd0.024315809143171958, 32'sd0.079338056412569, 32'sd0.02398321362927545, 32'sd0.007912428106691018, 32'sd-0.06434229186467591, 32'sd0.02938306115452103, 32'sd0.08385888347295198, 32'sd0.034834710412038, 32'sd0.0008851614187212236, 32'sd-0.018489505707890784, 32'sd0.07113212355460194, 32'sd0.11294046768518388, 32'sd0.07279252269218019, 32'sd0.0568834841341314, 32'sd0.06452129563166682, 32'sd0.060178726385420905, 32'sd0.04521983075579121, 32'sd-2.457829053651765e-122, 32'sd9.240567174172725e-116, 32'sd9.922097885918091e-124, 32'sd1.034011712372873e-124, 32'sd6.555260287340994e-122, 32'sd9.845990739898308e-123, 32'sd0.11176209152376096, 32'sd0.07538377536780261, 32'sd0.08387423436323269, 32'sd-0.011304068155074998, 32'sd0.026980752682758097, 32'sd0.04165857515098606, 32'sd0.06996162997479738, 32'sd0.12100953967893635, 32'sd0.058495500581144826, 32'sd0.021101973862997073, 32'sd0.12996362956305302, 32'sd0.039025400465396834, 32'sd0.03222699138611335, 32'sd0.0036771168031013803, 32'sd-0.05852063864462186, 32'sd-0.02618385872697679, 32'sd-0.07731888151600047, 32'sd0.10573286511586003, 32'sd0.14458161316405216, 32'sd0.0047611049852894615, 32'sd0.0010258136003386416, 32'sd0.10260456418439504, 32'sd0.09467936247231841, 32'sd0.0902481239519427, 32'sd-6.892400620789928e-126, 32'sd3.3518549243025186e-115, 32'sd4.970197685997161e-129, 32'sd-1.8897522454263688e-116, 32'sd-0.03188565591525061, 32'sd-0.025211922445201113, 32'sd-0.016131775038318853, 32'sd0.10780221279261058, 32'sd0.05353551724775186, 32'sd0.052563342295744005, 32'sd0.043370286728418785, 32'sd-0.01244470146012528, 32'sd-0.041485021981995183, 32'sd-0.06733938227902318, 32'sd0.051698586097668565, 32'sd0.03303290028431229, 32'sd0.038865387183345895, 32'sd-0.07741985188183063, 32'sd0.011004920056775957, 32'sd-0.11368087529471198, 32'sd-0.14530671162483708, 32'sd-0.13836047845679753, 32'sd0.04255878507874945, 32'sd-0.01951648850937514, 32'sd-0.027019652770312652, 32'sd-0.0033067775982115284, 32'sd0.0951300566122217, 32'sd0.012230471655835892, 32'sd-0.049954594498696825, 32'sd9.112509057040917e-118, 32'sd-2.160203325484723e-126, 32'sd0.04178346250173083, 32'sd0.026821765472822164, 32'sd-0.005997364636513402, 32'sd-0.07760483526233031, 32'sd-0.05727389003096313, 32'sd0.01799814770956025, 32'sd0.026435181423814198, 32'sd-0.03698773875835965, 32'sd0.011587511460489775, 32'sd-0.045699342288926414, 32'sd0.07360405928173096, 32'sd0.03272220464913415, 32'sd-0.034239456320977045, 32'sd-0.05348918367694315, 32'sd-0.028234338116810902, 32'sd-0.1068963843386175, 32'sd-0.09194923481489728, 32'sd0.05301870820026093, 32'sd-0.002040475024987497, 32'sd0.06610699816317925, 32'sd0.11123658457759089, 32'sd-0.006656922062963065, 32'sd0.04282940114113818, 32'sd-0.0029221712237914297, 32'sd-0.10021647883721384, 32'sd-0.010366529345541645, 32'sd0.11098826973401991, 32'sd-4.141039878288517e-123, 32'sd0.057792176457267044, 32'sd-0.01442916240436051, 32'sd0.012920244066875941, 32'sd0.02207546230656465, 32'sd0.07417842266651217, 32'sd-0.03598512925766996, 32'sd-0.038092169365579735, 32'sd0.09024182822765289, 32'sd-0.07291573551108929, 32'sd-0.11496111887697076, 32'sd-0.1298983828055074, 32'sd-0.1267223396338283, 32'sd-0.17886811267309216, 32'sd-0.036028470996081655, 32'sd-0.1626841508135881, 32'sd-0.1450065971963636, 32'sd0.054018693764942755, 32'sd-0.06932554450112301, 32'sd0.09222798822753558, 32'sd0.060783605003165785, 32'sd0.06803111105948442, 32'sd-0.10465571250534875, 32'sd-0.04338290575527023, 32'sd-0.06411413074838712, 32'sd-0.014575813789307461, 32'sd-0.029022265678887816, 32'sd-0.017772453335221032, 32'sd6.954765076508898e-120, 32'sd0.05045862048914467, 32'sd0.05921450905621988, 32'sd-0.005132620974518225, 32'sd0.09916964933240834, 32'sd0.02425245163239404, 32'sd0.036612204294692786, 32'sd-0.02786531387138661, 32'sd0.055523758102861566, 32'sd-0.09217215761841077, 32'sd-0.041426756798379726, 32'sd-0.11189595673737113, 32'sd-0.035393574545273046, 32'sd-0.016242326586178357, 32'sd-0.02751583746343307, 32'sd-0.055147655488901465, 32'sd0.014805071580999361, 32'sd-0.05913893735685142, 32'sd0.019154508934682127, 32'sd-0.00239302011630668, 32'sd-0.020530734797828923, 32'sd0.08468689768276026, 32'sd0.07222935794897473, 32'sd-0.004912621267542846, 32'sd-0.067748773560143, 32'sd0.022464706429146736, 32'sd-0.020823274480009767, 32'sd0.09026988758288475, 32'sd0.11958036170444158, 32'sd0.02302856416294971, 32'sd0.05128714806207464, 32'sd0.04392351702328191, 32'sd0.00677895695292733, 32'sd-0.013973810190029043, 32'sd0.06298165708363979, 32'sd0.02489878006653785, 32'sd-0.05393309162639121, 32'sd-0.15297822268784012, 32'sd-0.11013397924852401, 32'sd-0.073121612181583, 32'sd0.0116958808133494, 32'sd0.06842259711009847, 32'sd-0.06028584670061334, 32'sd-0.11916034380460505, 32'sd0.07267655277319043, 32'sd0.07133620510905252, 32'sd0.09241716508375618, 32'sd0.05312103840482313, 32'sd-0.05818515420402045, 32'sd0.05893944186541664, 32'sd0.0033252361450497804, 32'sd-0.06420778734281472, 32'sd0.07481467886428894, 32'sd0.07002138640287968, 32'sd0.040586140226497744, 32'sd0.01903694253952747, 32'sd0.07142361878718242, 32'sd0.024651158911693387, 32'sd0.04359844615377067, 32'sd-0.009988441567936298, 32'sd0.007415111598749633, 32'sd-0.10595711548713083, 32'sd0.050329273965087566, 32'sd0.006791987924071187, 32'sd-0.030708769021774444, 32'sd-0.07508260651431194, 32'sd0.07516822308861486, 32'sd-0.030879480217344057, 32'sd0.028577526393874515, 32'sd-0.12346249880663511, 32'sd-0.031505313928099306, 32'sd0.01558916255780555, 32'sd0.0020944984654204446, 32'sd0.12550931899397064, 32'sd0.038256019359897586, 32'sd-0.07920462827547128, 32'sd0.10497879995033238, 32'sd-0.05986186733328558, 32'sd0.0038309246326627103, 32'sd-0.046716886054970146, 32'sd0.023650749135324542, 32'sd-0.012852450919876204, 32'sd-0.09183972930193998, 32'sd0.05235196397730456, 32'sd0.07566982364442949, 32'sd0.10700438180598833, 32'sd0.0653847269444049, 32'sd0.012017129599991848, 32'sd0.08055253883804209, 32'sd-0.08790471060624863, 32'sd0.0031997658832718916, 32'sd-0.07914652096740678, 32'sd-0.028599993155649085, 32'sd0.08147670725704677, 32'sd0.13689732367857682, 32'sd0.0802634268919766, 32'sd0.00858623919258787, 32'sd-0.007137977946936189, 32'sd-0.004599360599631151, 32'sd-0.03274741312919976, 32'sd0.008214231455202762, 32'sd0.021383479100179913, 32'sd0.012708472127287408, 32'sd0.11489487817323034, 32'sd0.018365229023072187, 32'sd0.08809593516983395, 32'sd0.041219498468621794, 32'sd0.020756500248453748, 32'sd0.008896846080577642, 32'sd0.028657460365648736, 32'sd-0.07584986124075983, 32'sd0.04012265701848432, 32'sd0.09204969667690047, 32'sd-0.01612945177980052, 32'sd0.17720122506435404, 32'sd0.0023405343432678733, 32'sd0.07443567017329866, 32'sd0.027100636753736224, 32'sd0.031482582174844266, 32'sd0.0849541905345107, 32'sd-0.0009838690496219685, 32'sd0.03557028799032434, 32'sd0.09783386033350587, 32'sd0.10273355626729966, 32'sd0.041166392500925984, 32'sd0.13448607638490664, 32'sd0.059457854893935444, 32'sd0.02927145081582741, 32'sd0.10927725358196211, 32'sd-0.027629428720387778, 32'sd0.13908419054482316, 32'sd0.012441042224565381, 32'sd0.06240129772435914, 32'sd0.14761676260908865, 32'sd0.10059317357816916, 32'sd-0.08275244417908259, 32'sd0.09566105352032164, 32'sd0.03952751495802709, 32'sd0.025296731547313652, 32'sd0.09466127021262233, 32'sd0.008425990753320718, 32'sd0.07301932573290401, 32'sd0.052029002124521335, 32'sd0.08273417966768701, 32'sd0.05536725718659854, 32'sd0.0459509748637448, 32'sd0.04608912097528694, 32'sd0.12468614277319083, 32'sd0.051429685764676915, 32'sd0.0251687461757689, 32'sd0.0029804663738250015, 32'sd0.22053753591459477, 32'sd0.02349541722435436, 32'sd0.14763795073696562, 32'sd0.23898482350714004, 32'sd0.198828216714653, 32'sd0.04992888721753743, 32'sd-0.027852879333132335, 32'sd0.05263472412036284, 32'sd0.1112704061029157, 32'sd0.1434627030437686, 32'sd0.11133471404858274, 32'sd0.16975368490312837, 32'sd0.07166639654886807, 32'sd0.08870531131552072, 32'sd-0.023190679428594457, 32'sd-0.034295551902727706, 32'sd0.01868410193134624, 32'sd0.044620132666231396, 32'sd0.04902494356416895, 32'sd-0.003991509793765213, 32'sd0.1005792777463313, 32'sd0.11872049048598231, 32'sd0.1829363479421653, 32'sd0.07379123529544976, 32'sd0.09223602304320565, 32'sd0.09352403959259258, 32'sd0.14469287822252916, 32'sd0.16030084374796127, 32'sd0.26782455909727765, 32'sd0.17426101921056278, 32'sd0.08473501921804089, 32'sd0.01579287751203345, 32'sd0.07406976126407261, 32'sd0.0004286414232881325, 32'sd-0.056744603941100015, 32'sd-0.0013305505102741534, 32'sd-0.01744965159431639, 32'sd0.11264190225180842, 32'sd0.17351483308873153, 32'sd0.08892550787695128, 32'sd0.09792024294773856, 32'sd0.029212034502986005, 32'sd-0.029486690991685622, 32'sd0.0039825971215062764, 32'sd-0.02366812282467752, 32'sd0.052707944567654666, 32'sd-0.06729992557196496, 32'sd0.05966671053551655, 32'sd-0.020681830297563496, 32'sd0.10372513845549781, 32'sd0.22714834742684123, 32'sd0.11051293628460108, 32'sd0.1081260661955682, 32'sd0.0413405713952153, 32'sd0.03010151507454832, 32'sd0.14384381845371616, 32'sd0.06297474302938416, 32'sd0.0007032853138905545, 32'sd-0.07372853053804966, 32'sd-0.15954694407914646, 32'sd-0.1773191554797642, 32'sd-0.1315703243104441, 32'sd-0.2569775385397254, 32'sd-0.06033798132636763, 32'sd-0.05745540721911201, 32'sd-0.035613837153613645, 32'sd0.10043944833387371, 32'sd0.15816147885706666, 32'sd0.15871673811902418, 32'sd-0.03243886787115613, 32'sd0.06032296912519923, 32'sd0.08024512436524275, 32'sd0.025152696256705916, 32'sd0.04525918111105514, 32'sd-0.054984711517018135, 32'sd-0.01948308748692174, 32'sd0.09631156019140352, 32'sd0.13354794356561778, 32'sd0.032650911411339315, 32'sd0.10585256720664783, 32'sd0.03689089054640336, 32'sd0.16455087228861487, 32'sd-0.0012168653644085555, 32'sd-0.02654572420094264, 32'sd-0.086845771502204, 32'sd-0.14584632341907233, 32'sd-0.1722044168998288, 32'sd-0.18198118864181587, 32'sd-0.020653185498936685, 32'sd-0.1936917031197815, 32'sd-0.19793466890539135, 32'sd-0.052698052781782856, 32'sd-0.10210309376686191, 32'sd0.07144794076784644, 32'sd0.12094803210860332, 32'sd0.16658106158656313, 32'sd0.0863865202727167, 32'sd-0.14846466432660813, 32'sd-0.16549871531111482, 32'sd-0.0095961515237127, 32'sd0.048437717284641524, 32'sd0.027093537809038448, 32'sd0.03662340127345632, 32'sd-0.01695422379481573, 32'sd0.04769345942286517, 32'sd0.049191841902408794, 32'sd-0.020355824093160273, 32'sd0.09903900391148969, 32'sd0.016014314914603207, 32'sd0.0341301977455, 32'sd-0.07813266394184135, 32'sd-0.0256878649580493, 32'sd-0.09582178892863542, 32'sd-0.13007359401415639, 32'sd-0.030450279973606307, 32'sd-0.008370600751544182, 32'sd-0.059880948405382224, 32'sd-0.1479955993037626, 32'sd-0.13644033837338773, 32'sd-0.12670197728010998, 32'sd-0.12449758649197182, 32'sd0.029234117423360344, 32'sd0.10085698538855126, 32'sd0.09052052730488093, 32'sd-0.037482786968822825, 32'sd-0.03581693845479823, 32'sd0.030430289119838128, 32'sd-0.05134183725307739, 32'sd0.05548524147303421, 32'sd0.045288506803331054, 32'sd-0.05496346947132533, 32'sd-0.023333070701790488, 32'sd-0.06324607721171098, 32'sd-0.02598066914171351, 32'sd0.08093693288792532, 32'sd-0.03264087967779405, 32'sd0.06170569613379094, 32'sd-0.003948767386165821, 32'sd-0.0796612958858213, 32'sd-0.04823347432671722, 32'sd-0.17964598918908578, 32'sd-0.194407364835282, 32'sd-0.1611961962601133, 32'sd-0.07588521528241393, 32'sd-0.0704361464863272, 32'sd-0.10250539910609208, 32'sd-0.10982388602527578, 32'sd-0.0663099882053598, 32'sd-0.06139711829007611, 32'sd0.049414573963342964, 32'sd0.027511875997838796, 32'sd0.07674968088532118, 32'sd0.09521595085234634, 32'sd-0.012964672662038726, 32'sd-0.07191081494589034, 32'sd-0.00922326452810284, 32'sd-0.01660995765731987, 32'sd1.4795182828980183e-124, 32'sd0.041467156812083336, 32'sd-0.022222821967529862, 32'sd0.007456448356551508, 32'sd0.05657998649860901, 32'sd0.06951095940401096, 32'sd0.0009733622616311724, 32'sd0.08776445788739501, 32'sd0.01275202821107763, 32'sd0.010204820534784534, 32'sd-0.13133326146929541, 32'sd-0.18297716055300048, 32'sd-0.0930647585072242, 32'sd0.008992393060968924, 32'sd-0.08622895286573631, 32'sd-0.07543998860991895, 32'sd-0.18761200636211353, 32'sd-0.0008617181458308508, 32'sd-0.04944849380089877, 32'sd0.07707492382905702, 32'sd0.004923071634915421, 32'sd0.03865770623447948, 32'sd0.12309952918846406, 32'sd0.01983910662829559, 32'sd-0.07733715793320717, 32'sd0.05469450711198294, 32'sd0.001157288512759669, 32'sd0.01866665671419643, 32'sd0.04008496448979363, 32'sd0.005586836358954364, 32'sd-0.08077720680495935, 32'sd-0.003589330665073963, 32'sd-0.04050706495367967, 32'sd-0.08666820732036706, 32'sd-0.03026636790807332, 32'sd0.06262917080931805, 32'sd0.12100277752976427, 32'sd0.06734459801657657, 32'sd-0.01063482025402754, 32'sd-0.09720222686680093, 32'sd-0.10472787166586554, 32'sd0.03097137572457415, 32'sd-0.02675899661798495, 32'sd-0.015695269341653193, 32'sd-0.09678893480287291, 32'sd0.08037391077978194, 32'sd0.07792453635323396, 32'sd-0.0483682231197653, 32'sd-0.01508289520108796, 32'sd0.03313791691340181, 32'sd0.08889350424228233, 32'sd-0.029377273708323014, 32'sd-0.028669029368251952, 32'sd-0.0065576589101554, 32'sd0.02420445128428834, 32'sd0.013397288795828995, 32'sd0.051726072286802434, 32'sd0.03733715906205591, 32'sd0.015396915778197124, 32'sd0.07819223261817138, 32'sd0.026563999323978592, 32'sd0.03303582195349318, 32'sd-0.0702656004275143, 32'sd0.08992891239593181, 32'sd0.06859119377547684, 32'sd0.0566468653241182, 32'sd0.08296689610756947, 32'sd-0.06079962345593922, 32'sd0.09573879750420991, 32'sd-0.0521035679234327, 32'sd-0.05044778049619646, 32'sd0.037935639516591145, 32'sd0.035855295601672464, 32'sd0.10297901786533517, 32'sd0.025709630704436333, 32'sd-0.08424262513706983, 32'sd0.05423688620316946, 32'sd-0.13826164464793733, 32'sd-0.041440455214155625, 32'sd-0.029329259425964534, 32'sd0.02264012985641329, 32'sd0.04527138976597495, 32'sd-0.10508700324389332, 32'sd0.031137537732398017, 32'sd-2.776563674199043e-120, 32'sd0.05750838414691167, 32'sd-0.09510277629507007, 32'sd-0.014347078475607653, 32'sd-0.009317319956281036, 32'sd-0.07261941315017742, 32'sd-0.035064088804320034, 32'sd0.09232428774373382, 32'sd0.16974929107636358, 32'sd0.09696991977322011, 32'sd0.13701639018913317, 32'sd-0.07030475063945761, 32'sd-0.01697202480260532, 32'sd0.08396325219256487, 32'sd0.006833221046144643, 32'sd-0.10268156262728237, 32'sd0.01688024184373108, 32'sd-0.021803036924287356, 32'sd0.009048704948289932, 32'sd-0.17994376660533526, 32'sd-0.1251920146064927, 32'sd0.001322723080512654, 32'sd0.012853111359020085, 32'sd-0.0802460081807184, 32'sd-0.044879725568596394, 32'sd0.12117562226259272, 32'sd-0.018402260329079427, 32'sd0.06453139993214217, 32'sd-0.0354358602295297, 32'sd0.003841201732699221, 32'sd0.02213248983915671, 32'sd0.08390895644431505, 32'sd-0.062031373321449, 32'sd-0.08878574577461887, 32'sd0.007335846525769317, 32'sd0.1709461823381369, 32'sd0.1183166159097463, 32'sd-0.006128855614955371, 32'sd-0.003841056915965637, 32'sd-0.022404800216109945, 32'sd0.06651212263316163, 32'sd-0.07982803226996284, 32'sd-0.119942817273966, 32'sd-0.036221187226773095, 32'sd0.029729706738292012, 32'sd-0.11285850535346025, 32'sd-0.0744932512942512, 32'sd-0.1565943194204281, 32'sd-0.12632401000635649, 32'sd0.008966321542826717, 32'sd-0.09289240671574142, 32'sd0.023231429685184962, 32'sd0.042831817154791896, 32'sd0.05175101062125955, 32'sd-0.049746862059440976, 32'sd-0.0030673669893830826, 32'sd0.03665501908178738, 32'sd-0.020621171269677253, 32'sd-0.12736720122903442, 32'sd0.09476315904521372, 32'sd0.04154020047759492, 32'sd0.07000055298073371, 32'sd0.02639238700869936, 32'sd0.08875815851957282, 32'sd0.13684282603777828, 32'sd0.09525345705034914, 32'sd0.07204935265694863, 32'sd0.01753522380039999, 32'sd0.008558859744872437, 32'sd0.04206241593813218, 32'sd-0.08908880806723356, 32'sd-0.028082706387654033, 32'sd-0.11894737202937893, 32'sd0.060220127055154754, 32'sd-0.051943042833175905, 32'sd-0.10085316241001115, 32'sd-0.13795728965231666, 32'sd-0.08328547320949897, 32'sd0.09487509758658978, 32'sd0.026012144880219062, 32'sd0.07045901046757724, 32'sd0.11498926064463233, 32'sd-0.05953139325700565, 32'sd0.07711511003329763, 32'sd-3.841703405565921e-116, 32'sd0.0480032727783811, 32'sd0.012931832429746194, 32'sd-0.10059947062922019, 32'sd-0.06501330552415514, 32'sd-0.03741290708151098, 32'sd-0.005374477211600229, 32'sd-0.03311310233263593, 32'sd0.04720824913008831, 32'sd-0.052901863303138855, 32'sd0.053289801319507286, 32'sd-0.001541495617980464, 32'sd-0.047138340170253645, 32'sd0.02712817996558022, 32'sd-0.0035696854685430338, 32'sd0.012450513629605154, 32'sd0.10202854465330259, 32'sd0.011829671810921176, 32'sd-0.006233379186354432, 32'sd-0.09021118992261015, 32'sd-0.05059139539560513, 32'sd-0.1074641813057895, 32'sd-0.04293344837836479, 32'sd0.04067233077473628, 32'sd-0.025766060672233818, 32'sd0.026445008026225503, 32'sd0.013793137508353797, 32'sd-3.470449428133299e-119, 32'sd-1.0961495478728664e-120, 32'sd-3.312110859663238e-120, 32'sd-0.07430505355142099, 32'sd0.0023464899601546756, 32'sd0.09120271501407427, 32'sd0.1118105489037684, 32'sd-0.007200072685206663, 32'sd0.004975875102025211, 32'sd0.04621980629013957, 32'sd-0.010085876708950886, 32'sd0.12483885869381837, 32'sd0.003016839822049621, 32'sd0.1297393868307442, 32'sd0.04814759667990818, 32'sd-0.005313835414661828, 32'sd0.013515629217595592, 32'sd0.08294788643852267, 32'sd0.13155793034752938, 32'sd-0.039591525351013325, 32'sd-0.03177306695901237, 32'sd-0.006673191380580031, 32'sd-0.05807373159874907, 32'sd-0.002966381124408978, 32'sd-0.0363140175490122, 32'sd-0.02648946699140619, 32'sd-0.06640460710558298, 32'sd0.09895569590465327, 32'sd7.647643164138783e-117, 32'sd-1.4237691738046051e-125, 32'sd-8.925532833832418e-120, 32'sd0.07840085264197409, 32'sd0.042884104500456634, 32'sd-0.04142101138787177, 32'sd-0.03744811132609253, 32'sd-0.022162208369248773, 32'sd0.004003061578177294, 32'sd-0.05907987653390276, 32'sd-0.024566115584233952, 32'sd0.031152047591266694, 32'sd-0.037822726798748436, 32'sd-0.17424330509693045, 32'sd-0.09763852651382382, 32'sd0.029606788239724638, 32'sd-0.02935800253501919, 32'sd0.19030407688575324, 32'sd-0.03893409525367066, 32'sd-0.1933969277838535, 32'sd-0.07535279504263111, 32'sd-0.004271778396533944, 32'sd-0.04451416722915039, 32'sd0.06845988163275679, 32'sd0.05106043528125976, 32'sd0.0042241941375116355, 32'sd0.09492362120039752, 32'sd0.0449500383613168, 32'sd1.79981556043014e-123, 32'sd-1.7046803543276936e-123, 32'sd-6.812704706133966e-118, 32'sd-5.023352158052482e-118, 32'sd0.051643909092740914, 32'sd0.052147592676870726, 32'sd-0.025471390369562585, 32'sd-0.010879149855996643, 32'sd-0.0872347661595003, 32'sd0.03498004350218339, 32'sd0.02303827635028754, 32'sd-0.03773344078020658, 32'sd0.007830584413388277, 32'sd-0.024508572458399686, 32'sd0.11446768106658624, 32'sd0.0601748637129722, 32'sd0.1296676953794195, 32'sd0.07984522114464991, 32'sd-0.002989972722012567, 32'sd-0.099505102866764, 32'sd0.051848359454452306, 32'sd-0.04491522387609021, 32'sd-0.025349340486536406, 32'sd0.09999566809186808, 32'sd-0.062076636079997916, 32'sd0.10830179932891269, 32'sd0.11792627927673267, 32'sd-7.70846582002139e-126, 32'sd-3.9909040861025966e-126, 32'sd-6.662437784327451e-126, 32'sd5.231566711261046e-125, 32'sd-1.0722643164802474e-124, 32'sd-1.0744517896088678e-123, 32'sd0.046182998035154375, 32'sd0.06571530172320707, 32'sd0.02735049684750867, 32'sd0.002003698257812914, 32'sd0.13837819728117787, 32'sd0.01591939300816211, 32'sd0.13571460621059914, 32'sd-0.018201037748641128, 32'sd0.06330073654668492, 32'sd0.023854249783257807, 32'sd0.11967480905515256, 32'sd-0.007220923370406583, 32'sd0.17053242715036326, 32'sd0.07413311851122215, 32'sd0.03967417882798246, 32'sd-0.05632234167470877, 32'sd-0.002591810703300406, 32'sd0.09661713954410453, 32'sd0.1500435488112679, 32'sd0.058527229609118187, 32'sd1.4355225513497718e-122, 32'sd7.021153516412456e-116, 32'sd1.2437591515404385e-116, 32'sd1.2195452513103073e-121},
        '{32'sd1.0483997105683838e-127, 32'sd-8.696075632603293e-122, 32'sd-8.604707383254111e-117, 32'sd5.722916791950364e-121, 32'sd2.0878125998074664e-126, 32'sd4.815586103246213e-118, 32'sd-3.387664601539319e-123, 32'sd1.016455490447119e-124, 32'sd1.4270752604844916e-125, 32'sd-7.527040486139849e-124, 32'sd-2.116232516902464e-127, 32'sd4.697389055463542e-115, 32'sd0.07967230360702317, 32'sd0.09569385598766222, 32'sd0.04777385331309479, 32'sd0.018837661613191538, 32'sd-2.4613095551139406e-122, 32'sd-3.1146441183828344e-118, 32'sd2.54990875818112e-126, 32'sd1.0754773904945274e-124, 32'sd-1.0192763766255604e-119, 32'sd1.3342729287264032e-122, 32'sd-5.709801631975198e-115, 32'sd2.4317346408862383e-119, 32'sd-5.561763523128446e-115, 32'sd2.892654205293785e-125, 32'sd7.314466560640699e-116, 32'sd3.734897944919391e-122, 32'sd1.1279184569518655e-119, 32'sd-2.9423168690754405e-128, 32'sd-1.4688609535426128e-119, 32'sd-2.4382630030436507e-121, 32'sd0.003779257795606728, 32'sd0.07796562675131519, 32'sd-0.10206906403029034, 32'sd-0.022552208108527205, 32'sd-0.03825686052940816, 32'sd-0.044855878833532266, 32'sd0.081518365391464, 32'sd0.06040584984426188, 32'sd0.05037548617406635, 32'sd0.11258326520766107, 32'sd0.012719429632765568, 32'sd-0.026694455893721526, 32'sd-0.05771083154031457, 32'sd0.04690153905427961, 32'sd-0.03825277911982984, 32'sd-0.05080085660675559, 32'sd0.05134183910631111, 32'sd0.0669726767016402, 32'sd-0.004487792367428299, 32'sd0.04749711107726116, 32'sd1.7330278386876074e-125, 32'sd1.4057391317951247e-115, 32'sd-1.1306017799115741e-116, 32'sd-3.521062324818266e-114, 32'sd4.263337178385112e-125, 32'sd2.6851155187667793e-116, 32'sd0.12444926978756844, 32'sd0.010431932937133504, 32'sd0.0283466450872653, 32'sd-0.07189229327084026, 32'sd0.0348439047517697, 32'sd0.06512829069379646, 32'sd-0.089543831292868, 32'sd-0.0884676770500879, 32'sd0.11778361335648127, 32'sd0.031031372769914693, 32'sd-0.029656740967108394, 32'sd0.0438029751570813, 32'sd0.03756273684991903, 32'sd-0.05810677215614269, 32'sd0.021934601081682797, 32'sd-0.06308339352628477, 32'sd-0.012295568709020896, 32'sd-0.03629627009139765, 32'sd0.04677748940874154, 32'sd0.14588281710285872, 32'sd0.009900941087622152, 32'sd0.07189825561129706, 32'sd0.05022831315659811, 32'sd0.07402213207779802, 32'sd-1.2258008450996585e-127, 32'sd-1.275818969435542e-116, 32'sd-1.075055973784076e-124, 32'sd5.723567837014276e-127, 32'sd0.03436584426357271, 32'sd-0.00551276871926278, 32'sd-0.012738907783194047, 32'sd0.06159483605252587, 32'sd0.03657185352329288, 32'sd0.05024393021971032, 32'sd-0.044002531393875534, 32'sd-0.1593639475643462, 32'sd-0.09584568754306254, 32'sd0.0022062753398327103, 32'sd-0.031199987927893573, 32'sd-0.06611140643686136, 32'sd-0.05432330135916442, 32'sd-0.10747735187790537, 32'sd-0.24008338578016303, 32'sd-0.1160717383810282, 32'sd-0.07702189430595233, 32'sd0.1153190949156361, 32'sd0.04008851770038705, 32'sd-0.027187771681662965, 32'sd0.025998727021168497, 32'sd-0.03325589484987753, 32'sd0.07667192858947587, 32'sd0.006857233924198563, 32'sd0.029652173198591217, 32'sd-4.1465684823190484e-123, 32'sd3.444674109411641e-129, 32'sd0.0747289189807931, 32'sd0.05416133017106962, 32'sd0.04917336796279522, 32'sd-0.018039175576674043, 32'sd-0.04202997231460979, 32'sd-0.029897984052803347, 32'sd-0.10042903684789228, 32'sd-0.0007563831122729952, 32'sd-0.022764453161086134, 32'sd-0.12767287544599465, 32'sd0.05898214950663449, 32'sd0.009414010620096162, 32'sd-0.036813197720639, 32'sd-0.018981048242040676, 32'sd-0.11388174544310255, 32'sd0.08079356717017508, 32'sd0.06636111060199741, 32'sd0.055162332507215535, 32'sd0.1313642314550666, 32'sd0.11785718155720697, 32'sd0.0657820778874038, 32'sd0.023192963832441182, 32'sd0.01402525125931951, 32'sd0.03537481266384685, 32'sd-0.07504834239502786, 32'sd0.1356236255176381, 32'sd0.02921943341222223, 32'sd2.132869274622323e-127, 32'sd0.08044676772613325, 32'sd-0.009447463147144754, 32'sd0.04722519314716216, 32'sd-0.060591608206783984, 32'sd0.05157103518849221, 32'sd0.04223109206060411, 32'sd-0.03909035599731223, 32'sd-0.012783568413732634, 32'sd0.09466455762541263, 32'sd-0.005096901538791547, 32'sd-0.12327252946442155, 32'sd-0.14244778225181612, 32'sd-0.09030438199830286, 32'sd-0.18739856616473685, 32'sd-0.14747402239454577, 32'sd0.0038431614955173245, 32'sd-0.03508133443122912, 32'sd0.15051225661418335, 32'sd0.11926825547749856, 32'sd0.1586263184933614, 32'sd0.05335866400971436, 32'sd0.035351495713675, 32'sd0.14588039169954886, 32'sd-0.05563281695238445, 32'sd-0.06898572020334494, 32'sd-0.01800072871477953, 32'sd0.005764024757799706, 32'sd6.4044597823446e-125, 32'sd0.019032484830865542, 32'sd-0.0006993166314517075, 32'sd-0.06360661926229585, 32'sd0.10895924863417793, 32'sd0.012435348993784253, 32'sd0.1603785446226451, 32'sd0.11720458585440757, 32'sd0.06829755646814305, 32'sd0.057070881752997966, 32'sd-0.02466084874849414, 32'sd0.0005076392497956956, 32'sd-0.019679941332207265, 32'sd-0.09657652383436031, 32'sd-0.20011131323562145, 32'sd-0.2649003236996921, 32'sd-0.07299918943317367, 32'sd0.09177877413467969, 32'sd0.10799568645427692, 32'sd0.14104900080572075, 32'sd0.07876854895735146, 32'sd0.15076901822411848, 32'sd-0.040078356611305654, 32'sd-0.038572524524876195, 32'sd-0.07431542301866642, 32'sd-0.11257966330053608, 32'sd0.0030466436130206563, 32'sd0.0412074026398377, 32'sd0.12657856115601618, 32'sd0.02693780434341926, 32'sd0.034521650685940077, 32'sd0.0260534161427137, 32'sd0.032726312032265635, 32'sd-0.03960829571644879, 32'sd0.05171034713016398, 32'sd0.08319301414509243, 32'sd-0.08121417919572439, 32'sd0.10966748793272997, 32'sd0.03064828164055637, 32'sd-0.09609929970560202, 32'sd-0.03617495197033646, 32'sd-0.09966823433733646, 32'sd-0.19732753215684717, 32'sd-0.19430233401002836, 32'sd0.06982751621657683, 32'sd0.2685606542560934, 32'sd0.2305845273653468, 32'sd0.20818083864116851, 32'sd0.052444693065204495, 32'sd0.1012615574554114, 32'sd0.1018068586655008, 32'sd0.057107146948561845, 32'sd-0.0026325038166674394, 32'sd-0.10792727234965163, 32'sd-0.052503360840928034, 32'sd0.012418863467499666, 32'sd0.05573513772334405, 32'sd0.0570387392429412, 32'sd-0.08390103848184095, 32'sd0.042215998582684204, 32'sd-0.09763051652213979, 32'sd-0.060113114413084666, 32'sd0.027391401357166167, 32'sd0.04398404543759151, 32'sd-0.08029908463170124, 32'sd0.034021846336395024, 32'sd0.014401922212042123, 32'sd-0.07225122703597718, 32'sd-0.06403779780308096, 32'sd-0.25028974041799545, 32'sd-0.30252622066635354, 32'sd-0.21282712453609656, 32'sd0.07914532798761446, 32'sd0.15995522751551766, 32'sd0.2399912152678947, 32'sd0.18650971469816535, 32'sd0.045549400645024454, 32'sd-0.048240084181975576, 32'sd0.052914514608499566, 32'sd0.06168495997065134, 32'sd-0.08554266867775732, 32'sd0.01584702376962175, 32'sd0.06985307390111385, 32'sd0.033385919072482076, 32'sd0.09234206480724237, 32'sd0.03597520549790236, 32'sd-0.030983458543797398, 32'sd0.03126104437422373, 32'sd-0.04267589045295936, 32'sd-0.14240694080100816, 32'sd-0.006687366587692158, 32'sd-0.039114725384743476, 32'sd-0.001472379006616676, 32'sd-0.046978042058414174, 32'sd-0.02087444766583551, 32'sd0.060339658931233664, 32'sd-0.011218522883491273, 32'sd-0.3320915426893499, 32'sd-0.30976753437100446, 32'sd0.04315706068093268, 32'sd0.16295878408904385, 32'sd0.26363571005736697, 32'sd0.13578706033871019, 32'sd0.08288477192757626, 32'sd-0.04946193950677275, 32'sd-0.02872347551757013, 32'sd0.0827530775844502, 32'sd-0.01403106261900398, 32'sd-0.009271348456302094, 32'sd0.003916799343535047, 32'sd-0.018259211501671084, 32'sd0.003642536996440166, 32'sd0.07940174764965442, 32'sd0.010192082030121273, 32'sd-0.010995370917502436, 32'sd-0.053368314566458755, 32'sd-0.0672999721490717, 32'sd0.03307971381283102, 32'sd0.05725361332771337, 32'sd-0.049316634731212186, 32'sd0.0059378174824368385, 32'sd0.09577277324706454, 32'sd0.015296071093251172, 32'sd-0.05535794225742517, 32'sd-0.14134712186696996, 32'sd-0.3010831044588365, 32'sd-0.1955967991211965, 32'sd0.18078909196189022, 32'sd0.20057060716967656, 32'sd0.2025915094485357, 32'sd0.05605090570539822, 32'sd-0.037463713695944874, 32'sd-0.09689637936400626, 32'sd-0.11509103578861248, 32'sd-0.018259061771623477, 32'sd-0.009550861449545756, 32'sd0.016680604521671017, 32'sd0.0892086754765955, 32'sd-0.09434494421549233, 32'sd-0.04088013165268004, 32'sd0.09742581692731421, 32'sd0.03914508840128782, 32'sd-0.04074317754616524, 32'sd-0.01822968121825108, 32'sd-0.05082772621340008, 32'sd-0.06612344625930099, 32'sd0.040378168299752965, 32'sd0.005368901959897814, 32'sd-0.07476390796386467, 32'sd0.013684516368511335, 32'sd0.05248603957456606, 32'sd-0.0840609709465614, 32'sd-0.15035381628218455, 32'sd-0.038826180748097336, 32'sd0.006944773995914433, 32'sd0.14570949591743748, 32'sd0.14715690480324498, 32'sd0.19564129058279048, 32'sd0.15106559169209896, 32'sd0.016124988989697654, 32'sd-0.015810387456084655, 32'sd-0.026742403737812576, 32'sd0.004019864248064625, 32'sd-0.09513637888634106, 32'sd-0.027007034498307513, 32'sd-0.03948536889296304, 32'sd0.0026316087773657166, 32'sd0.06066376588622913, 32'sd-0.020327358444932234, 32'sd0.004257788867177395, 32'sd0.025595583857822103, 32'sd-0.1228379812970499, 32'sd-0.02873649706906781, 32'sd0.0637280206903507, 32'sd-0.10371380075164133, 32'sd-0.07605406420533598, 32'sd0.03754087820288215, 32'sd0.13386581519210472, 32'sd-0.04248095365975773, 32'sd-0.17264011643005225, 32'sd-0.09767371014904976, 32'sd-0.07484125846530654, 32'sd0.004845885160047942, 32'sd0.10007179033210645, 32'sd0.05897973175045092, 32'sd0.04056511385928453, 32'sd0.07779142446934188, 32'sd-0.06199723341401341, 32'sd-0.15624091627536413, 32'sd-0.1299017680730304, 32'sd-0.05808941899401332, 32'sd0.012432996449105315, 32'sd0.08311693056215234, 32'sd0.07021709960180256, 32'sd0.013725875919508683, 32'sd0.057511851733102706, 32'sd0.03908388741721862, 32'sd0.023313273236817096, 32'sd0.010811843437946349, 32'sd-0.016748776192094497, 32'sd0.027068464760007106, 32'sd0.029168118176747988, 32'sd0.07297504873172984, 32'sd0.005647743160897759, 32'sd0.016229596526039208, 32'sd0.06432500957030043, 32'sd-0.08718865131130266, 32'sd-0.1207982809416074, 32'sd-0.09171825426248441, 32'sd-0.0912501769507241, 32'sd0.05054063578978186, 32'sd0.051231301178670245, 32'sd0.06215886480751288, 32'sd0.0845726710950121, 32'sd0.009262696201160263, 32'sd-0.001696328268467417, 32'sd0.007130136895715694, 32'sd0.026784327869543333, 32'sd0.051438143567354495, 32'sd-0.06281098551043132, 32'sd0.013391473759600907, 32'sd0.04885246826266015, 32'sd0.02612069924483748, 32'sd-0.07179130651893322, 32'sd0.06875377421992988, 32'sd0.003657386594562751, 32'sd0.014264741651832412, 32'sd0.000500589185780432, 32'sd0.03118075562001631, 32'sd0.06234692611403103, 32'sd0.02381051283079793, 32'sd0.026698695902249003, 32'sd-0.05840510712460787, 32'sd0.01636730009639353, 32'sd-0.025836782408988346, 32'sd0.056570828082122764, 32'sd-0.11296256859137324, 32'sd0.05758332873383537, 32'sd0.1469693518419558, 32'sd0.028470857846077762, 32'sd0.08633415648606399, 32'sd0.08881485508210761, 32'sd0.10001878839559267, 32'sd0.09114895986224349, 32'sd-0.014527956140787638, 32'sd0.0538266301225764, 32'sd-0.05385147073881696, 32'sd0.026606608799669328, 32'sd-0.03161514364548685, 32'sd0.04303261656374659, 32'sd-0.0026101808151899972, 32'sd0.01906420745289294, 32'sd-0.0888217146238085, 32'sd-0.03859209235361179, 32'sd0.01582642639568955, 32'sd0.043426114849711456, 32'sd-0.05440572243997343, 32'sd-0.04509635661259812, 32'sd-0.08520100862912881, 32'sd-0.023408174530729537, 32'sd-0.08753375179960902, 32'sd-0.10420127757516762, 32'sd-0.06715673974383338, 32'sd0.14412277050676134, 32'sd-0.09953393981001869, 32'sd0.07198360144486028, 32'sd0.05862109475479147, 32'sd0.013003517030932986, 32'sd0.015377166081454325, 32'sd0.012537151265745413, 32'sd-0.0058591168948771526, 32'sd0.0956839277043347, 32'sd-0.033680996821843584, 32'sd-0.051451571104175677, 32'sd-0.017120993559242268, 32'sd0.05452591065429634, 32'sd-0.06774294364478645, 32'sd0.021150958551783474, 32'sd0.04051474211001538, 32'sd0.0778224189780131, 32'sd0.03673894710806163, 32'sd0.0810684047130787, 32'sd-0.013158641223649783, 32'sd-0.007386499125188258, 32'sd0.03317465253349903, 32'sd-0.04731282435229839, 32'sd0.022793073467658697, 32'sd0.022452285487742422, 32'sd0.01904050979891791, 32'sd-0.05174414340021054, 32'sd0.07603644506700288, 32'sd-0.029836982768265127, 32'sd0.10718985320632149, 32'sd0.08661652146999015, 32'sd0.021955752581066405, 32'sd-0.003141437399136531, 32'sd0.03732084665857169, 32'sd0.050308674886706074, 32'sd0.052683484734359666, 32'sd0.02930504417888211, 32'sd0.052050967203646235, 32'sd0.00465099907490344, 32'sd-0.06564351383597086, 32'sd0.0122847700961957, 32'sd0.11002050136542772, 32'sd-0.0035130103713980755, 32'sd0.012187459204021216, 32'sd0.02298178614510382, 32'sd5.1800217252509615e-127, 32'sd0.0218655600626028, 32'sd-0.12959980496720278, 32'sd-0.061110441957601, 32'sd0.012638919272160584, 32'sd-0.03415872301603949, 32'sd-0.026901670968857254, 32'sd0.05935139228907866, 32'sd-0.02668930250250349, 32'sd-0.05007415519872584, 32'sd-0.06251437339743647, 32'sd0.052261064313105884, 32'sd0.03443152058697872, 32'sd0.16988306182258953, 32'sd0.1340034304711465, 32'sd-0.03832443906354983, 32'sd0.00013592459545899607, 32'sd0.04978393382147973, 32'sd0.10936118077350535, 32'sd0.15783052890952717, 32'sd0.10006194254576783, 32'sd0.08448930807519682, 32'sd0.030596412892719378, 32'sd-0.028366747584661373, 32'sd0.05056631865708143, 32'sd0.0166636829853156, 32'sd0.0027808985965912876, 32'sd0.006452426997065271, 32'sd-0.0038261154043797998, 32'sd0.048839664612355865, 32'sd0.023628245420077888, 32'sd-0.09248237910280761, 32'sd-0.0034098537752070683, 32'sd-0.060875855699247576, 32'sd-0.05250903706300925, 32'sd-0.06808082819472311, 32'sd0.008372668488046532, 32'sd0.07543869562705627, 32'sd-0.05798583883448711, 32'sd-0.020290282696816663, 32'sd-0.06987432423032239, 32'sd0.12882505993671073, 32'sd0.02558090524710208, 32'sd-0.0868901996155277, 32'sd-0.009575284309593781, 32'sd0.08144858590800674, 32'sd0.01146549903831838, 32'sd-0.0787693884426677, 32'sd0.003939675557086531, 32'sd-0.10637728037199809, 32'sd-0.016039329780309596, 32'sd-0.061057292459405416, 32'sd-0.15156764302230558, 32'sd-0.009646091810512524, 32'sd0.01861805718776038, 32'sd0.00826925640779237, 32'sd0.09089124671874231, 32'sd-0.07192721383133516, 32'sd0.08323566224750077, 32'sd0.04563867158124943, 32'sd-0.11051856431685986, 32'sd-0.10091482048660416, 32'sd-0.03412923660950113, 32'sd0.07419516476636531, 32'sd-0.10706594283416604, 32'sd0.08699216427429834, 32'sd-0.035453721236753444, 32'sd0.004408379504280439, 32'sd-0.013084872847142786, 32'sd-0.06718926600148725, 32'sd0.00624104290318342, 32'sd-0.03189843699495557, 32'sd-0.014845672816568638, 32'sd-0.052284563133284556, 32'sd-0.022886037389267165, 32'sd0.024895204381303312, 32'sd-0.034821341302206786, 32'sd-0.020619858838099275, 32'sd-0.05899908813164602, 32'sd-0.07417582996769294, 32'sd0.007814666793509438, 32'sd0.04264053985859428, 32'sd0.0026416215675955194, 32'sd0.033093045636362874, 32'sd-7.299843776248499e-115, 32'sd-0.010885508567628994, 32'sd-0.015249730981712699, 32'sd0.1760984495509815, 32'sd0.06965633576589104, 32'sd-0.06596211983824213, 32'sd-0.05077685457922076, 32'sd-0.03823929307267729, 32'sd0.016238587183586894, 32'sd-0.05674948113427634, 32'sd-0.09411444601568356, 32'sd-0.038283965269544806, 32'sd-0.026907572991139123, 32'sd-0.04793013818092821, 32'sd-0.04062352962890671, 32'sd-0.035056183310114536, 32'sd-0.06390668733535265, 32'sd-0.0036991576218406512, 32'sd0.034037296142085935, 32'sd-0.1259109212044086, 32'sd0.05175767141704469, 32'sd0.13083393105819774, 32'sd0.0039432086318529486, 32'sd0.1426643800181673, 32'sd-0.036474330210688057, 32'sd-0.055520751790138566, 32'sd-0.014418777557307883, 32'sd0.04987724473281934, 32'sd0.015906350309648373, 32'sd-0.0004109392701728821, 32'sd0.019413524059769937, 32'sd0.047288726139125443, 32'sd-0.016281399317782056, 32'sd-0.010569764155951587, 32'sd0.06388740593883398, 32'sd-0.08631564093020162, 32'sd0.01409196948656658, 32'sd-0.059830105549422904, 32'sd-0.009717821175781296, 32'sd0.027610948037065118, 32'sd0.0007149131329269524, 32'sd-0.010977665631842068, 32'sd-0.02589268500129731, 32'sd-0.12892064604593986, 32'sd0.034074037918917985, 32'sd0.038005756948869374, 32'sd-0.07557262012829545, 32'sd-0.08660973609410573, 32'sd0.04808431106940457, 32'sd0.08930407927492152, 32'sd0.07908680362017358, 32'sd0.0824392165877389, 32'sd0.021665001875642208, 32'sd-0.049714684593139304, 32'sd0.020192129146951843, 32'sd0.018606875885880305, 32'sd0.0625787173393062, 32'sd0.06466469281269625, 32'sd-0.006276977080014206, 32'sd0.0022794909719797427, 32'sd-0.058752224649782234, 32'sd0.1139919278773091, 32'sd0.0942084837593987, 32'sd-0.018174921954394286, 32'sd-0.04067003052611889, 32'sd-0.04303495718627691, 32'sd0.08372958694644073, 32'sd0.016881867489321457, 32'sd0.05453385725033473, 32'sd0.21870417491460825, 32'sd0.10281393520517272, 32'sd-0.05871079548679739, 32'sd0.004058788769361226, 32'sd0.0744108352994383, 32'sd0.0501162568264083, 32'sd-0.032587897404454606, 32'sd0.0005998648529439233, 32'sd0.0168858701603493, 32'sd-0.029682069120569015, 32'sd-0.11866205992459941, 32'sd0.03154986988365615, 32'sd-0.07027151678690316, 32'sd0.04431285598825586, 32'sd0.09057073304645874, 32'sd-6.401286454679294e-120, 32'sd0.10764269990233481, 32'sd-0.04239436074102311, 32'sd-0.0689019411111444, 32'sd0.009839425801091976, 32'sd0.018767758710940774, 32'sd0.004185062433867493, 32'sd0.1294621209300598, 32'sd-0.007812518349568568, 32'sd0.08849370358079628, 32'sd0.04165477436806581, 32'sd-0.007453224439243353, 32'sd0.08353897925092653, 32'sd0.14812079754494922, 32'sd0.03170166440918482, 32'sd0.012377309695089277, 32'sd0.0670439184586331, 32'sd0.03324482035986755, 32'sd-0.06416524228332629, 32'sd-0.07680062130790713, 32'sd-0.015519505530105903, 32'sd-0.034672382689083105, 32'sd0.016153257922046367, 32'sd0.05263738399383377, 32'sd0.014433228413601798, 32'sd0.053248075323772605, 32'sd0.06782493305525239, 32'sd-2.1388424277360033e-119, 32'sd-8.777105029807673e-116, 32'sd1.0714059344385894e-116, 32'sd0.05030194879376042, 32'sd0.08828044169404727, 32'sd-0.04521623529731823, 32'sd0.03481233562899411, 32'sd-0.01855058078241732, 32'sd0.028501836617312384, 32'sd-0.060422158718670196, 32'sd-0.01605044722381529, 32'sd0.03871997695739754, 32'sd-0.05944859929996758, 32'sd0.05813508610014859, 32'sd0.07348278563299127, 32'sd-0.0022494491706737613, 32'sd-0.07063390838074418, 32'sd-0.03591661551990255, 32'sd-0.04658117387813986, 32'sd-0.024045023559423805, 32'sd0.05193922829741625, 32'sd0.12645293876688268, 32'sd-0.03881193265408713, 32'sd0.05526153461914206, 32'sd0.044935982414533844, 32'sd-0.037601171036259234, 32'sd0.07908716316376972, 32'sd0.026399256584214218, 32'sd1.4931678104520767e-115, 32'sd1.2944360623435457e-121, 32'sd-3.5460757780178985e-116, 32'sd0.03285811023093558, 32'sd0.03570617030681058, 32'sd-0.04411203729544734, 32'sd0.07558613819100185, 32'sd-0.028125822782210416, 32'sd-0.05138671513740965, 32'sd0.00485319657948459, 32'sd-0.01443761906231282, 32'sd-0.07686786222374817, 32'sd-0.0474075199832657, 32'sd0.10987674227090856, 32'sd0.13741263898260736, 32'sd0.04993103715182283, 32'sd-0.15703577075043498, 32'sd-0.11462427741004158, 32'sd-0.1242458983375601, 32'sd0.018921692442791252, 32'sd-0.05307072739032775, 32'sd0.15134337337537818, 32'sd-0.03919768276011503, 32'sd0.0376974162946899, 32'sd-0.010931683334437394, 32'sd-0.03905248373964673, 32'sd-0.04791382820780753, 32'sd-0.05116166290690773, 32'sd1.8091266924760373e-122, 32'sd1.4965556343637332e-128, 32'sd5.408950810595762e-121, 32'sd-4.8062943656703075e-117, 32'sd0.09454454649826942, 32'sd0.04741100200065809, 32'sd-0.07770541427427376, 32'sd0.012928465427234574, 32'sd-0.00043696341911185987, 32'sd0.06586345931186327, 32'sd0.019223395785417652, 32'sd0.03597707689714144, 32'sd0.020934487318325652, 32'sd0.06676205696965173, 32'sd-0.011166739159964263, 32'sd-0.07974862720499505, 32'sd0.0007940665061374818, 32'sd-0.04683423915271496, 32'sd0.012075069051928122, 32'sd0.04943652820956019, 32'sd0.10716145032429165, 32'sd0.09698051557774671, 32'sd-0.050424296284579395, 32'sd0.15031359800010222, 32'sd0.044793908184646083, 32'sd-0.013235725717134652, 32'sd0.0745075352619378, 32'sd8.540033513095045e-122, 32'sd3.866110156091524e-128, 32'sd-1.682945855177561e-125, 32'sd2.1382809696222135e-127, 32'sd-1.399359108444809e-125, 32'sd5.598440224983468e-115, 32'sd0.0946836150263721, 32'sd0.14833336497700778, 32'sd0.055627867588408826, 32'sd0.17916997420484396, 32'sd0.043827268338930865, 32'sd-0.0471639393695123, 32'sd-0.028172414011151194, 32'sd-0.0545636168900115, 32'sd0.062395199943441254, 32'sd0.07879935573622429, 32'sd0.073792136695843, 32'sd0.03795681978042672, 32'sd0.059010699428170894, 32'sd-0.009294637591973059, 32'sd-0.08224830691652175, 32'sd0.005824800667849849, 32'sd-0.03486160949520586, 32'sd0.004590969633954171, 32'sd0.03181103274128673, 32'sd0.0864937608955418, 32'sd4.878727021962173e-115, 32'sd-7.392226239432882e-117, 32'sd7.572856696294681e-127, 32'sd2.893167748353696e-129},
        '{32'sd2.1222480992464883e-116, 32'sd-3.0286985873362334e-116, 32'sd-4.386870806976942e-117, 32'sd5.026588766969368e-118, 32'sd-8.157077939277735e-117, 32'sd-1.0452716671234247e-120, 32'sd-4.3195228792278606e-121, 32'sd-7.281478636953601e-125, 32'sd1.3656862859426167e-118, 32'sd-1.455365118023018e-114, 32'sd-2.1039298966916887e-124, 32'sd8.663088847632864e-115, 32'sd-0.002017727312279786, 32'sd-0.043849953048168896, 32'sd0.04412090253296877, 32'sd-0.017799524604578513, 32'sd1.4333539381377035e-118, 32'sd-2.599276426682807e-126, 32'sd-3.4342745749514395e-126, 32'sd-1.095351952947507e-119, 32'sd1.1172312573401862e-125, 32'sd7.564539961925873e-115, 32'sd5.399773492345636e-122, 32'sd8.550868845073863e-127, 32'sd2.2461121830467907e-123, 32'sd4.18240254824632e-125, 32'sd7.633223020250942e-117, 32'sd-1.5155345792025414e-117, 32'sd1.6303150294846782e-115, 32'sd-3.341891263739336e-125, 32'sd1.7363704011037977e-125, 32'sd-3.078945426143799e-122, 32'sd0.02665838097538289, 32'sd-0.07131848049212765, 32'sd0.0013731305060447003, 32'sd-0.11808366674048608, 32'sd0.026321091559412802, 32'sd-0.0024103052332647905, 32'sd0.008632547614146035, 32'sd-0.020646392076326778, 32'sd-0.008621175432136714, 32'sd-0.05206207909533145, 32'sd-0.031839655339443156, 32'sd-0.12038410990446236, 32'sd-0.020342536963684838, 32'sd0.0015103613690884215, 32'sd0.0477662239962685, 32'sd-0.07176131990769538, 32'sd0.01502693027150958, 32'sd0.055995648660521584, 32'sd0.04589945956260376, 32'sd-0.00872402294458992, 32'sd1.3278530648955313e-118, 32'sd-2.401156307012361e-127, 32'sd4.372743145129871e-126, 32'sd-1.0229939617307321e-120, 32'sd7.60031361914142e-122, 32'sd6.387781481969715e-124, 32'sd0.028284125359132408, 32'sd0.07371384987616889, 32'sd-1.8330416552335132e-05, 32'sd0.05661870845319388, 32'sd-0.05049207606889141, 32'sd0.039616073864469, 32'sd-0.029344923630161092, 32'sd-0.0891586266235708, 32'sd0.014448763732984798, 32'sd-0.09410493327787887, 32'sd-0.012976807083275053, 32'sd-0.06370071911235957, 32'sd-0.028490085762005915, 32'sd-0.18702586793332157, 32'sd-0.11726394859943741, 32'sd0.026853833200761464, 32'sd-0.147080644634931, 32'sd-0.04719592252161805, 32'sd-0.023087789606893575, 32'sd0.0097635500023474, 32'sd-0.06988490032536031, 32'sd-0.0543630659600163, 32'sd0.00637376518666011, 32'sd0.0955727499173786, 32'sd-8.853902697707031e-125, 32'sd1.0963733496763897e-121, 32'sd1.5357834286011238e-124, 32'sd-6.955577760191066e-124, 32'sd-0.014525999813638085, 32'sd0.013601355655815358, 32'sd0.002397163776766969, 32'sd-0.09677337997517939, 32'sd0.046468851508759006, 32'sd0.10802683190508237, 32'sd-0.0983295147846865, 32'sd-0.0946314872873314, 32'sd0.017136200382359443, 32'sd0.08446331121495373, 32'sd-0.12832297479898847, 32'sd-0.06764763317305923, 32'sd-0.013896748856778256, 32'sd-0.011056027569607593, 32'sd-0.1865822326876152, 32'sd-0.12427200647015235, 32'sd-0.007950188832348885, 32'sd-0.0019176167201327176, 32'sd-0.055617238801659696, 32'sd0.08609809099917502, 32'sd0.047105290722967715, 32'sd-0.032294774447789845, 32'sd-0.024318476064235227, 32'sd0.11421281726552272, 32'sd-0.04470599703029479, 32'sd-2.3654200926095348e-124, 32'sd1.1590205394401948e-115, 32'sd-0.0022965532081368465, 32'sd0.0377865776426531, 32'sd-0.05977833639839402, 32'sd-0.1418136381115877, 32'sd0.025107851273944333, 32'sd0.10691211872717153, 32'sd0.017760079456615653, 32'sd-0.01899681222773763, 32'sd-0.10992143821082363, 32'sd-0.18143085499211795, 32'sd-0.05856217516390404, 32'sd-0.10590278564476437, 32'sd-0.05510769935897141, 32'sd0.032951123197838814, 32'sd0.07069438179153982, 32'sd-0.06763843873333485, 32'sd-0.09181711107448319, 32'sd-0.13726129204888995, 32'sd-0.17918889245782535, 32'sd0.046777560064098445, 32'sd-0.04849525152212349, 32'sd0.0903901013068905, 32'sd0.017297862211576857, 32'sd-0.06201522781087083, 32'sd0.07719709448066302, 32'sd0.06531194365431679, 32'sd-0.03470608728975428, 32'sd7.522873838407047e-119, 32'sd0.02581082404917076, 32'sd0.0049856735014313725, 32'sd0.033917228242176634, 32'sd-0.20260093809785368, 32'sd-0.18994349476022915, 32'sd-0.008151226675631926, 32'sd0.061184653308684556, 32'sd0.05015884064446716, 32'sd0.050936629960701016, 32'sd-0.022681055329874786, 32'sd0.04720320781818478, 32'sd-0.01959583518633825, 32'sd-0.10231047849112818, 32'sd-0.12606221957990216, 32'sd-0.0032123413367918887, 32'sd-0.11582169412661424, 32'sd-0.0700853462788916, 32'sd-0.11230548251416983, 32'sd-0.136914793686649, 32'sd-0.01941822356541525, 32'sd-0.051593167441208995, 32'sd-0.025139681202937542, 32'sd0.07683504527536655, 32'sd0.0429951349897359, 32'sd-0.07722616222012853, 32'sd-0.025944154821917066, 32'sd0.02219475851461254, 32'sd-1.0228286040360778e-124, 32'sd0.014937745674448048, 32'sd-0.08820320653655113, 32'sd0.06432530616449417, 32'sd-0.07487862290781787, 32'sd-0.024538744206325656, 32'sd0.03724547353457361, 32'sd0.06684311563719356, 32'sd-0.05009436998679706, 32'sd0.14916269267607674, 32'sd0.0832663552837179, 32'sd0.02640899107202257, 32'sd-0.0802520994735238, 32'sd0.06360414384947864, 32'sd0.09603685814375987, 32'sd-0.05020493349919738, 32'sd-0.022606371733374625, 32'sd-0.017433134678917207, 32'sd0.006961082949189715, 32'sd-0.009932787125714623, 32'sd0.07984083123010886, 32'sd0.099595790585725, 32'sd0.00857765681571649, 32'sd0.03365676722591979, 32'sd0.0763050836207052, 32'sd-0.06676427583826186, 32'sd0.025094623460320042, 32'sd-0.044381522076909666, 32'sd0.010434435674049976, 32'sd0.06429495386075333, 32'sd-0.036815402904380366, 32'sd0.11248581845197411, 32'sd-0.03717027002581815, 32'sd-0.00020171180128280734, 32'sd-0.052054211625308225, 32'sd-0.03689524228751652, 32'sd-0.014672565366552755, 32'sd0.03412440186552579, 32'sd-0.10181780516201107, 32'sd-0.08019016632216375, 32'sd0.025418028327697316, 32'sd0.07627296710456091, 32'sd-0.0336742439080492, 32'sd-0.008225394146137098, 32'sd-0.04435734667043363, 32'sd-0.0983943865926415, 32'sd-0.022133318337752395, 32'sd0.002694441010720527, 32'sd-0.007235126970578988, 32'sd0.07307638775124427, 32'sd-0.03400482889591495, 32'sd-0.019190308785972554, 32'sd-0.10590405516089076, 32'sd-0.02734410839677667, 32'sd-0.04579594693676795, 32'sd-0.011377083753718325, 32'sd-0.031673140063217045, 32'sd-0.009868392263842658, 32'sd-0.03219900359307295, 32'sd0.0007469769073621388, 32'sd-0.07044029382696884, 32'sd-0.07353702106495577, 32'sd0.03863079107056611, 32'sd-0.06155484167582351, 32'sd0.023922744616737546, 32'sd-0.04588570543070318, 32'sd-0.05841119568989012, 32'sd0.004052512632877024, 32'sd-0.028687366863648082, 32'sd0.02770393385307379, 32'sd0.002315199149746981, 32'sd-0.04371205540628919, 32'sd-0.21321984002736588, 32'sd-0.14758522055437603, 32'sd-0.104421107683462, 32'sd-0.010755860563607021, 32'sd-0.08897552652101286, 32'sd0.08598556365698569, 32'sd-0.05201755085790941, 32'sd0.028451082263282225, 32'sd0.0011248287432501867, 32'sd0.025844795689660707, 32'sd-0.02240903047157884, 32'sd-0.056120127580128715, 32'sd0.03258333734975455, 32'sd0.11443813643732356, 32'sd0.1303863372527332, 32'sd0.03186159717734215, 32'sd-0.008352748728133288, 32'sd-0.005872396687388766, 32'sd0.029415220026378506, 32'sd-0.08466208125905247, 32'sd0.04779294600664849, 32'sd0.014273018981696656, 32'sd-0.07329633425693106, 32'sd0.05205429091664836, 32'sd0.09881946497157199, 32'sd-0.09890238267016713, 32'sd-0.04435076969849279, 32'sd-0.13408802967421654, 32'sd-0.024963039534308094, 32'sd0.08301388873793827, 32'sd0.047435297026505896, 32'sd-0.09206697896302796, 32'sd-0.005328223618161716, 32'sd0.09703178396870427, 32'sd-0.08390412684362504, 32'sd-0.022508886575280943, 32'sd-0.06404011389012929, 32'sd-0.05514166111218488, 32'sd-0.014706979749907978, 32'sd0.03939160120480689, 32'sd0.07925615706863491, 32'sd0.05924370295120067, 32'sd-0.006724400467044273, 32'sd-0.006835663398303749, 32'sd-0.02823926787969846, 32'sd0.013078304138228924, 32'sd0.01169929727066606, 32'sd-0.030558175024619844, 32'sd-0.004027807404992045, 32'sd-0.12271350650757346, 32'sd-0.07696182994664777, 32'sd-0.06363886128593793, 32'sd0.062496723286868595, 32'sd0.02299668684670982, 32'sd-0.08396979496297483, 32'sd0.006649083050838913, 32'sd0.04475090840274873, 32'sd0.03514254843052071, 32'sd0.032091313661550915, 32'sd0.08679094153587284, 32'sd0.07405221961334578, 32'sd0.05600980582656658, 32'sd-0.014001371648458553, 32'sd-0.17270640994177447, 32'sd-0.033448110382381505, 32'sd0.10362581415540069, 32'sd-0.01555897342313196, 32'sd-0.054145898047023966, 32'sd0.07688754679071266, 32'sd-0.03704237622533829, 32'sd0.05040579898804562, 32'sd-0.08500749179141055, 32'sd-0.05066737310942437, 32'sd-0.11789661815672807, 32'sd-0.0038581866883511057, 32'sd-0.02026249624080936, 32'sd-0.02215315959783503, 32'sd-0.10282578079028383, 32'sd-0.01858382686825217, 32'sd0.016028217534163836, 32'sd0.03468983375012474, 32'sd-0.04227583603153902, 32'sd0.08850588870969171, 32'sd0.04328572256299292, 32'sd-0.008812249193906128, 32'sd0.13387496429860163, 32'sd0.12097119205408527, 32'sd0.04509503328513687, 32'sd-0.05017875479356222, 32'sd0.05092305053674866, 32'sd-0.05997584364338128, 32'sd-0.2232480280781494, 32'sd-0.16232334424930547, 32'sd-0.0007817649278301155, 32'sd-0.023115706364282545, 32'sd-0.0003411161456927254, 32'sd0.06930181663354615, 32'sd0.06480669096708369, 32'sd0.001326706319931083, 32'sd0.045000572403445585, 32'sd-0.11164314862410947, 32'sd-0.06615376932899364, 32'sd0.07361337655234754, 32'sd-0.056012659420494326, 32'sd0.06766337906218729, 32'sd-0.051338804414374835, 32'sd0.10769273612712471, 32'sd0.07573773260214849, 32'sd0.07599480808593477, 32'sd0.020798295368649466, 32'sd-0.011911638736337493, 32'sd0.061831724499656786, 32'sd0.06659301056779982, 32'sd0.04036419024352352, 32'sd-0.004250454524590034, 32'sd0.10633154302154874, 32'sd0.08102808618833497, 32'sd-0.019416314974083228, 32'sd-0.13061595446652347, 32'sd-0.1460053008401789, 32'sd-0.009151980218795952, 32'sd-0.006206043623460812, 32'sd0.0028369713584095865, 32'sd-0.06449150392283018, 32'sd0.0006436123753025363, 32'sd0.004801511668522615, 32'sd-0.09704481465608895, 32'sd0.036986378441712944, 32'sd-0.027106060953533705, 32'sd0.09550403717726244, 32'sd0.01318361861146278, 32'sd0.024840032234265317, 32'sd-0.04242547046292868, 32'sd-0.07378312973134886, 32'sd0.00846925392432312, 32'sd-0.0716112321386616, 32'sd-0.09092092738357932, 32'sd-0.0283173244725405, 32'sd0.04461326891305167, 32'sd-0.05936985815680893, 32'sd-0.015087513914616631, 32'sd0.01996172312840722, 32'sd0.0642303550198847, 32'sd0.005357881792480952, 32'sd0.07786905547598474, 32'sd0.039772628230875934, 32'sd-0.1608954900327122, 32'sd-0.2133056801488494, 32'sd0.01759271749235941, 32'sd-0.001969627951169157, 32'sd-0.15177100177813116, 32'sd-0.016047685306370026, 32'sd-0.016043985914098547, 32'sd0.006311270003381836, 32'sd-0.0727815086310089, 32'sd0.07969276204022788, 32'sd0.04973024743229888, 32'sd0.05479574209797835, 32'sd0.047603576943757824, 32'sd0.12108719209495918, 32'sd0.0346488903787517, 32'sd0.02245885414826765, 32'sd0.03795683321964515, 32'sd-0.04999567235215034, 32'sd-0.036115272845202356, 32'sd-0.14946883866530403, 32'sd-0.17177698231043814, 32'sd-0.023586203901228422, 32'sd0.017810610279098377, 32'sd0.12423256697150878, 32'sd0.16533007983541492, 32'sd0.06368386723637659, 32'sd-0.003317491144929558, 32'sd0.02755567115031118, 32'sd-0.008503365568669432, 32'sd-0.13447775344326846, 32'sd-0.033533001659020366, 32'sd0.05846761456108817, 32'sd0.10974543860641862, 32'sd0.016797745824936056, 32'sd-0.04213554924102476, 32'sd0.013263085581912849, 32'sd-0.04307790761432425, 32'sd-0.03854139189287664, 32'sd0.05361941923904736, 32'sd0.04549529543867499, 32'sd0.053736469206046494, 32'sd0.07815083746514372, 32'sd0.028418178819522265, 32'sd-0.043334196092746614, 32'sd-0.013679157334353763, 32'sd-0.06585844676890096, 32'sd-0.08959918763962442, 32'sd-0.18164186825817852, 32'sd-0.09558124953999221, 32'sd0.154804083299976, 32'sd-0.03316586805661673, 32'sd0.2131632979861894, 32'sd0.07315056963665852, 32'sd0.14284308504966045, 32'sd0.024429194744505615, 32'sd-0.04370187335687644, 32'sd0.0595251599973576, 32'sd-0.05081387499508818, 32'sd-0.04818718698067966, 32'sd0.04377821595969835, 32'sd-0.02266429242205317, 32'sd0.06893088278253358, 32'sd0.016953270601262182, 32'sd0.013103215963353222, 32'sd-0.092318603774264, 32'sd-0.06148062976820351, 32'sd0.028383027480147687, 32'sd0.06061586802073616, 32'sd0.047309628838375035, 32'sd0.18440877732277655, 32'sd0.17553067228837071, 32'sd-0.019887876864189517, 32'sd-0.004683684513574796, 32'sd-0.006244196551143847, 32'sd0.060277977563319034, 32'sd0.006489201106175072, 32'sd0.04240563942735803, 32'sd-0.008397513356937662, 32'sd-0.036570640177789854, 32'sd0.054998067968879065, 32'sd0.14446508130956126, 32'sd0.06818289876114685, 32'sd0.15627342132589297, 32'sd-0.024990758126988175, 32'sd0.08456278841852943, 32'sd0.006530701750146943, 32'sd-0.13414898338791909, 32'sd0.056954170493619144, 32'sd-0.05755095771883776, 32'sd0.011254693458875562, 32'sd-3.2857670280908083e-121, 32'sd0.03496214918392459, 32'sd-0.005688369275981508, 32'sd0.0018284397903516306, 32'sd-0.041053148126938846, 32'sd0.03108584912454551, 32'sd0.08574061582654172, 32'sd0.054708768064212064, 32'sd0.08130932473730498, 32'sd0.05334024534897686, 32'sd0.08777982457225059, 32'sd0.11049152065942415, 32'sd0.025946963592424793, 32'sd0.04792918778409385, 32'sd-0.023037324561152234, 32'sd0.03584360024124703, 32'sd0.03635507128686777, 32'sd-0.01761311694696679, 32'sd-0.03660520549276853, 32'sd0.06535561919083127, 32'sd-0.03917660364175343, 32'sd-0.07206604364071521, 32'sd-0.08804552539370933, 32'sd-0.11865817921901585, 32'sd-0.20739584836654584, 32'sd0.023306670621533368, 32'sd0.005488437392171334, 32'sd-0.01688562803658759, 32'sd0.018738291457894084, 32'sd-0.021679546340310447, 32'sd-0.04764812193133616, 32'sd-0.08252031767873795, 32'sd-0.07011044958390221, 32'sd-0.07482173111106125, 32'sd-0.06642816879917034, 32'sd0.05538764682020148, 32'sd0.1556999750150184, 32'sd0.1208576705681667, 32'sd0.15199625919603213, 32'sd0.22761312428847638, 32'sd0.10358261279399819, 32'sd0.06905461928214351, 32'sd-0.049602649532583865, 32'sd0.01680261134598738, 32'sd0.0399727160704131, 32'sd0.1093440596605185, 32'sd-0.14855871815043373, 32'sd-0.04216059083823579, 32'sd-0.07354077653847907, 32'sd-0.057163621793396034, 32'sd-0.19386518375728048, 32'sd-0.06068787245111142, 32'sd-0.21834596032952022, 32'sd-0.02386864231555043, 32'sd-0.01955477406299514, 32'sd-0.06529227153162423, 32'sd0.029310469634417625, 32'sd-0.03964349031834066, 32'sd-0.052715850983109346, 32'sd-0.06658948838742233, 32'sd-0.14200529743853146, 32'sd-0.0866019066726326, 32'sd-0.04722066747151128, 32'sd0.07743789345637424, 32'sd0.06218272579358992, 32'sd0.02305180446979639, 32'sd0.15210047178749322, 32'sd0.1807083424303783, 32'sd0.12041066150514232, 32'sd-0.07924742613046104, 32'sd-0.004436951513464381, 32'sd-0.03232491942967859, 32'sd-0.05288814373048246, 32'sd0.023875034927917295, 32'sd-0.14287855316922296, 32'sd-0.11370208653891639, 32'sd-0.05981146034721092, 32'sd-0.07309284981834453, 32'sd-0.18913649011072972, 32'sd-0.08537601825844475, 32'sd-0.12781437158331532, 32'sd0.005187185021280889, 32'sd0.010160741446862827, 32'sd0.05965595797053864, 32'sd3.242860074284386e-116, 32'sd0.03525853857263503, 32'sd-0.08234993382754052, 32'sd-0.04894619642663525, 32'sd0.029629019350242713, 32'sd-0.024146786195663565, 32'sd-0.05596298852948216, 32'sd-0.03979515347601593, 32'sd-0.05085630320482052, 32'sd-0.1198025737169402, 32'sd0.00679245770486491, 32'sd-0.06135984688592035, 32'sd-0.03153625670741523, 32'sd-0.09926506389732076, 32'sd-0.12535930657913041, 32'sd-0.060027427693321055, 32'sd-0.050981838064414774, 32'sd0.009100360606537952, 32'sd-0.038063757441484186, 32'sd0.05223742912357619, 32'sd-0.11309735116852575, 32'sd-0.12897908061974445, 32'sd-0.060251570730694884, 32'sd-0.05262260571180089, 32'sd-0.08952924519193933, 32'sd0.07258123461916725, 32'sd-0.1099551421546161, 32'sd0.042062011825260655, 32'sd-0.014403019329987471, 32'sd-0.041145379743805305, 32'sd-0.020087277024031257, 32'sd-0.03626124427459457, 32'sd0.0019555613754835503, 32'sd-0.02930012358406241, 32'sd-0.0008922059473569326, 32'sd-0.0003153585272896574, 32'sd-0.1533838717352436, 32'sd-0.06881266594358557, 32'sd-0.1929152435277219, 32'sd-0.2141698447830569, 32'sd-0.0966275773528653, 32'sd-0.2232327392971541, 32'sd-0.22295230802914637, 32'sd-0.10731154877238527, 32'sd-0.0525468200412901, 32'sd-0.04710938729595831, 32'sd-0.007819852959085815, 32'sd0.026014639786390424, 32'sd0.0018269754384242498, 32'sd0.024601790539946593, 32'sd0.08200773677127685, 32'sd0.03733373910687482, 32'sd0.04087999801012077, 32'sd0.07007394183279854, 32'sd-0.04936465167276204, 32'sd0.04318788665564341, 32'sd0.05139256239527328, 32'sd-0.003432575325208656, 32'sd0.018622170939955267, 32'sd-0.05499622280086771, 32'sd-0.04174548326615111, 32'sd-0.027008087886468128, 32'sd-0.04884782877843985, 32'sd-0.07513630215640897, 32'sd0.004086309577927473, 32'sd-0.10570419952459335, 32'sd-0.09632591960094466, 32'sd-0.14565883402629534, 32'sd-0.17568905943507981, 32'sd-0.1777572592827484, 32'sd-0.1284720248669234, 32'sd-0.17390535603498894, 32'sd0.036066694948546155, 32'sd-0.1428676143203036, 32'sd0.07410913974937411, 32'sd-0.010401140454204452, 32'sd0.06615524099148254, 32'sd0.04227548265729, 32'sd0.03333868302612617, 32'sd-0.037058464944173065, 32'sd0.016470186652473406, 32'sd0.1020709917144906, 32'sd-0.04448803541052936, 32'sd0.009898979443702022, 32'sd-3.635061449322532e-116, 32'sd0.06699843728941784, 32'sd0.030444112151060496, 32'sd-0.11813174171254386, 32'sd-0.009982058930508634, 32'sd-0.01228261941463906, 32'sd0.07135273590682352, 32'sd0.06561830978459365, 32'sd-0.03312567093954956, 32'sd-0.146416915180993, 32'sd-0.11991344298499192, 32'sd-0.09253904683883139, 32'sd-0.1393212909987566, 32'sd-0.11582417321807319, 32'sd-0.03402079011764414, 32'sd-0.11255840787308986, 32'sd-0.025072288207850207, 32'sd-0.06180443037027695, 32'sd-0.054174116248012834, 32'sd0.030272953387249276, 32'sd-0.0776105627437657, 32'sd0.0371568488122984, 32'sd0.08212502842865951, 32'sd-0.0010494535877715566, 32'sd0.007101343638678131, 32'sd0.016923913895585778, 32'sd0.00714993129913945, 32'sd-2.076111954018769e-117, 32'sd5.291564038586356e-122, 32'sd6.2230745234661415e-124, 32'sd-0.05191982344952169, 32'sd-0.014745358144420082, 32'sd-0.03351657916811555, 32'sd0.11815967483588033, 32'sd0.0017672312124957402, 32'sd0.08656797839322516, 32'sd-0.029729238433320787, 32'sd-0.03505496254931024, 32'sd-0.0958780084639427, 32'sd0.03118078976307222, 32'sd-0.20227810361223247, 32'sd-0.0715134155334972, 32'sd-0.03803815272308299, 32'sd-0.07971184873195616, 32'sd-0.06304332227923873, 32'sd0.033104682671532826, 32'sd-0.05452392707054497, 32'sd0.0352332860923706, 32'sd0.03344048334929849, 32'sd0.09003789674252828, 32'sd-0.03524732658391435, 32'sd0.0578324841002286, 32'sd-0.03913886114831002, 32'sd-0.018660607033576998, 32'sd0.038941519995776816, 32'sd3.655439516415781e-120, 32'sd-3.389132447649952e-122, 32'sd-2.172311169768914e-116, 32'sd0.03804961695057142, 32'sd-0.017711213463519407, 32'sd0.0734593800610684, 32'sd0.13141188785254265, 32'sd-0.04409465588204784, 32'sd0.03955028023222523, 32'sd-0.029119096884520097, 32'sd-0.17393515677967597, 32'sd0.0014185818436928015, 32'sd0.10321603711166982, 32'sd-0.06895555395630562, 32'sd-0.06598815341450211, 32'sd0.01186783639659134, 32'sd-0.1919005859738479, 32'sd-0.01999079435201506, 32'sd0.0575251037887739, 32'sd0.05200512467797321, 32'sd-0.018646361168301585, 32'sd-0.0586558644376864, 32'sd-0.017667431009131814, 32'sd0.09024586922960658, 32'sd0.06747805962024668, 32'sd0.039904606099515585, 32'sd0.025210569474733654, 32'sd-0.0695624334350131, 32'sd1.0528819985209265e-120, 32'sd-1.7946664669899656e-126, 32'sd-4.019665977977168e-122, 32'sd1.807882594095011e-123, 32'sd0.06750379575157087, 32'sd0.07192917980302556, 32'sd0.0698527210417074, 32'sd0.048068519737224605, 32'sd0.0069826020838465105, 32'sd-0.04137347849935707, 32'sd0.03281785313702988, 32'sd-0.027604024369880686, 32'sd-0.021391252910070196, 32'sd-0.10597754312878396, 32'sd-0.08601414369013782, 32'sd-0.008330147968728179, 32'sd-0.08984223140205395, 32'sd0.04352026464664466, 32'sd0.08277522289935754, 32'sd-0.01801521395662446, 32'sd-0.04014504212082275, 32'sd-0.03689010296686895, 32'sd-0.07468756651457328, 32'sd-0.05445635979933978, 32'sd-0.020785691058307756, 32'sd-0.016531418734545163, 32'sd0.03680454954924295, 32'sd4.578487670883947e-126, 32'sd8.633905282697506e-118, 32'sd2.924009960042925e-119, 32'sd-3.8035039260083424e-119, 32'sd3.3488091945252917e-121, 32'sd-6.757660152521116e-115, 32'sd0.030002549536050204, 32'sd0.06215478907840946, 32'sd-0.016302389190777884, 32'sd-0.01661608816335059, 32'sd0.009229228871747099, 32'sd-0.0380034689807648, 32'sd-0.027145622226901568, 32'sd-0.013507989017490748, 32'sd0.020493834386114226, 32'sd0.0017891188429993475, 32'sd0.013002246062437127, 32'sd0.01539886694352129, 32'sd0.01654216421769356, 32'sd0.059535994023114894, 32'sd0.06410128302563484, 32'sd0.04350907072531671, 32'sd0.0014535970983586932, 32'sd-0.07228397455220273, 32'sd0.08283190866088376, 32'sd0.02517930228479502, 32'sd-3.717860978604816e-120, 32'sd3.839771270050688e-122, 32'sd7.447856608067183e-124, 32'sd-1.5795543603269313e-125},
        '{32'sd-4.655041057901574e-126, 32'sd-9.417466222206543e-122, 32'sd-1.1118754478369392e-121, 32'sd-1.0419987801553197e-124, 32'sd-1.9194367740837995e-124, 32'sd-3.474213564534774e-123, 32'sd7.418278782290644e-126, 32'sd-1.5106666588083902e-116, 32'sd1.8074682594861127e-122, 32'sd9.404990421725767e-125, 32'sd1.0840125156964245e-126, 32'sd-7.577938111235674e-122, 32'sd-0.05676190025782758, 32'sd0.05558908280991584, 32'sd0.02417156453487107, 32'sd-0.05664771467663023, 32'sd-1.9876578880868705e-123, 32'sd-1.865858988467354e-126, 32'sd-8.928432449259695e-118, 32'sd-2.517043915800091e-116, 32'sd2.5973344401347237e-125, 32'sd5.761942734426712e-121, 32'sd-1.5475129429629866e-123, 32'sd-2.148697065055423e-120, 32'sd-6.6632303823805365e-115, 32'sd-7.224117755391746e-122, 32'sd1.3720863958536833e-121, 32'sd-8.836605569966104e-122, 32'sd-7.634727045240063e-125, 32'sd-4.082090671630989e-124, 32'sd-1.0680963181983366e-124, 32'sd5.542056375864299e-117, 32'sd0.07206316690538916, 32'sd0.023480779002618583, 32'sd-0.002854055715727577, 32'sd0.10619982974372318, 32'sd0.09112091625868451, 32'sd-0.0030403699816080533, 32'sd-0.0452848836376111, 32'sd0.07840506874871296, 32'sd0.014109609372638306, 32'sd0.023644076041535764, 32'sd-0.049860951926196946, 32'sd-0.010629218204376867, 32'sd0.10715494797332928, 32'sd0.023443427729195082, 32'sd-0.07675036779377109, 32'sd-0.008231241764711641, 32'sd-0.041173551462197776, 32'sd0.020092619730983887, 32'sd-0.012125591479208836, 32'sd-0.00990698862763864, 32'sd3.9860967224050684e-123, 32'sd-1.3729801857181476e-118, 32'sd8.210609562282809e-122, 32'sd2.3384621325447958e-122, 32'sd3.059549845057854e-126, 32'sd-2.0408412683261683e-127, 32'sd0.0009324320671459863, 32'sd-0.000748428438350362, 32'sd-0.0013521804233567168, 32'sd0.09882949769952377, 32'sd0.04106784865642103, 32'sd0.02733184064605897, 32'sd0.020980680986746568, 32'sd0.06163376990857456, 32'sd-0.06487654905977579, 32'sd0.05845830515778319, 32'sd0.05504610979224641, 32'sd-0.06864306576282674, 32'sd0.0002727079390653989, 32'sd-0.10975142899531788, 32'sd0.017103551288453357, 32'sd-0.006520757787513126, 32'sd0.013371348287756248, 32'sd-0.005182590395669708, 32'sd0.02895535162650102, 32'sd-0.06826195977777286, 32'sd0.05100873818407389, 32'sd0.011966858266610638, 32'sd0.0435157568722604, 32'sd-0.035019057583865636, 32'sd1.0900355888529332e-114, 32'sd6.156282930219248e-117, 32'sd-3.1469973353440027e-117, 32'sd-6.603979141384405e-115, 32'sd0.04437496541757087, 32'sd0.01963972964589671, 32'sd-0.038159817583474046, 32'sd-0.015345011144010372, 32'sd0.05889899426133337, 32'sd-0.08212820343704316, 32'sd0.03125507712487726, 32'sd0.03819686545281675, 32'sd-0.09180808165847437, 32'sd0.008751913326329035, 32'sd0.03939339171872628, 32'sd-0.022290715826699094, 32'sd4.0184767008260094e-05, 32'sd-0.06105687503915661, 32'sd-0.003401071687317524, 32'sd0.0846148572314358, 32'sd0.15765264461892234, 32'sd-0.08835302664065049, 32'sd-0.08198747993047732, 32'sd-0.11164982445666304, 32'sd-0.15242635703836369, 32'sd-0.10411739828120467, 32'sd0.019880551457926894, 32'sd0.03801551639936352, 32'sd0.05105133633801373, 32'sd-8.482286158627442e-127, 32'sd2.095872746933349e-124, 32'sd-0.02202421663977825, 32'sd-0.019294831134155737, 32'sd0.036987015552435866, 32'sd0.08761500601150975, 32'sd0.04079853519499237, 32'sd0.10099240031044943, 32'sd0.05482940257171928, 32'sd0.01666680856051097, 32'sd-0.06758441521355636, 32'sd-0.06938142529895919, 32'sd-0.07935201971910226, 32'sd-0.08267549989344761, 32'sd-0.08608264335912201, 32'sd-0.04068774322368433, 32'sd0.0731527957052138, 32'sd-0.03435429907368051, 32'sd0.09178746737682132, 32'sd0.11969623747602769, 32'sd0.017374517595775837, 32'sd0.016745453585261836, 32'sd-0.032167809320017594, 32'sd0.04018843421381866, 32'sd0.02276326558864015, 32'sd-0.0881582010150859, 32'sd0.00630197050125051, 32'sd0.03199159049494438, 32'sd-0.0014918128486001152, 32'sd-9.008600799880973e-121, 32'sd0.01912542654945304, 32'sd0.0148690243463501, 32'sd0.011167780120093621, 32'sd-0.04328068413966314, 32'sd-0.008393272946828222, 32'sd-0.0661421888170361, 32'sd0.025142467438972707, 32'sd0.009133821782006123, 32'sd-0.0347156129181654, 32'sd-0.049849481735350136, 32'sd0.027630246846051566, 32'sd-0.0371342737138677, 32'sd0.053177621539503096, 32'sd0.047970999802930916, 32'sd-0.0974750581168615, 32'sd-0.11874053175086789, 32'sd0.0640723349995479, 32'sd-0.018248804491055433, 32'sd8.255308407997251e-05, 32'sd-0.034451485709229734, 32'sd-0.07052704080881346, 32'sd-0.061652443753160834, 32'sd-0.09107454103327807, 32'sd-0.02758352587293001, 32'sd0.10034304163413077, 32'sd0.09747356846736828, 32'sd-0.038645359750843225, 32'sd-1.3423564792904264e-124, 32'sd0.024796492047952375, 32'sd0.0012884562875659909, 32'sd-0.07657031604362424, 32'sd-0.09072525100728838, 32'sd0.013243265746719461, 32'sd-0.03506533783058024, 32'sd-0.017179074636967977, 32'sd0.04923867555799145, 32'sd-0.07242705528173193, 32'sd0.0480216506501686, 32'sd0.0075406089505920225, 32'sd-0.029022917080158098, 32'sd-0.00026142440604438964, 32'sd-0.03455200944885156, 32'sd-0.01476008659936903, 32'sd-0.006339252120461654, 32'sd0.0614257753368829, 32'sd0.023409832039401893, 32'sd0.05473629044323226, 32'sd0.13281263526804576, 32'sd0.1352895969834887, 32'sd-0.004112799292727499, 32'sd0.026037076335821734, 32'sd0.051411530603804684, 32'sd0.05834575745082208, 32'sd-0.09467990859885594, 32'sd0.008270822313568797, 32'sd0.003695885888877572, 32'sd0.054686760813316665, 32'sd-0.0527993178951362, 32'sd-0.044357941561865205, 32'sd-0.03481694977526158, 32'sd0.05958017207650566, 32'sd-0.08046923548952223, 32'sd-0.06971042499724323, 32'sd0.050224796294009964, 32'sd-0.03411247112873982, 32'sd-0.0375754460978969, 32'sd-0.042740797049417446, 32'sd-0.11748382533694658, 32'sd-0.0010681225670692302, 32'sd-0.03046430227245095, 32'sd0.0730859358780896, 32'sd0.10452872838838087, 32'sd0.11928421717040005, 32'sd0.09206496009579786, 32'sd0.17520969469658057, 32'sd0.1433789429084318, 32'sd0.09484951043380342, 32'sd0.03209226765540391, 32'sd0.008210161270658788, 32'sd0.0333746042594197, 32'sd0.03890055855359206, 32'sd-0.07944203570461332, 32'sd0.01710758182360097, 32'sd0.002887805771629551, 32'sd-0.0702295819593834, 32'sd0.030834948856253777, 32'sd0.06098749832989414, 32'sd-0.0057939817564869826, 32'sd0.01810824153263025, 32'sd-0.00022587526863098288, 32'sd-0.002607179430774949, 32'sd0.05789416160264695, 32'sd-0.010132733327020652, 32'sd-0.03665279050117324, 32'sd-0.04327130477440515, 32'sd-0.027379612177976492, 32'sd-0.08023424688130919, 32'sd-0.001987577187362614, 32'sd0.09865598775458957, 32'sd0.1914939008425941, 32'sd0.13120757122112628, 32'sd0.0613119538741387, 32'sd0.09136797232906504, 32'sd0.05962285914890045, 32'sd0.015527889519614677, 32'sd0.039776447217157604, 32'sd-0.01959781663413602, 32'sd0.02290185888514482, 32'sd-0.08306824323943962, 32'sd-0.04232274095217149, 32'sd0.029285282050826627, 32'sd-0.03329883956115026, 32'sd-0.049790255534209224, 32'sd0.029178329933707885, 32'sd0.07538534322150435, 32'sd-0.04072972250892309, 32'sd-0.09239329991086297, 32'sd0.040630444040992156, 32'sd-0.04591378642611352, 32'sd-0.007182665289319112, 32'sd-0.0070121811498459795, 32'sd-0.09434047240006238, 32'sd0.01073575116208664, 32'sd0.01418445650095648, 32'sd0.025623820707670223, 32'sd-0.06389916472770651, 32'sd-0.13548654203591065, 32'sd-0.05077685277473832, 32'sd0.028766943960415608, 32'sd-0.07477030867271943, 32'sd-0.020438464579399712, 32'sd0.00848737078794702, 32'sd0.08241887052166677, 32'sd-0.03339057380587186, 32'sd0.08406315648545046, 32'sd0.025253067662071974, 32'sd0.048709208636097005, 32'sd0.008342921326870796, 32'sd-0.050372471046759085, 32'sd0.003722506397639053, 32'sd0.004648447374830633, 32'sd0.015876674662593685, 32'sd0.055593679122378885, 32'sd0.008653758425637616, 32'sd-0.021618244950071298, 32'sd-0.08492408232377865, 32'sd-0.1558780035555965, 32'sd-0.12351969062091606, 32'sd-0.00226037822166729, 32'sd-0.015420072546461801, 32'sd-0.015087744854319983, 32'sd0.006886114931025407, 32'sd-0.014663968115798539, 32'sd-0.1690751316586067, 32'sd-0.13602378925971673, 32'sd-0.1785562168756129, 32'sd-0.2553412366444834, 32'sd-0.09430941948908897, 32'sd-0.12934853148061423, 32'sd0.014226820427003796, 32'sd-0.03906866304611865, 32'sd-0.009036273296526705, 32'sd-0.04329944336539744, 32'sd-0.006046830942695742, 32'sd0.038686560293493454, 32'sd0.009150451460171611, 32'sd0.0318971754970124, 32'sd0.04917449403032406, 32'sd-0.06733969557501589, 32'sd-0.05522393414728097, 32'sd-0.11659637078752444, 32'sd-0.07829580459232323, 32'sd-0.04255073777467361, 32'sd-0.05437070520644755, 32'sd-0.0461592826783538, 32'sd0.05686295927304793, 32'sd0.10953144848714523, 32'sd0.06471173176774717, 32'sd0.10211721828505214, 32'sd-0.04676754674547783, 32'sd-0.22236654838086864, 32'sd-0.03893327762097524, 32'sd-0.0667964850257478, 32'sd-0.15557146846918304, 32'sd-0.050219292525556125, 32'sd-0.06767792762465819, 32'sd0.015063291141942443, 32'sd0.09709397297385208, 32'sd0.13591522360914726, 32'sd0.129009969955442, 32'sd0.18231338066019578, 32'sd0.1510258516454807, 32'sd0.07993027602625924, 32'sd-0.016474822753220455, 32'sd0.10197767865018922, 32'sd0.05406198572623628, 32'sd-0.06278241277639783, 32'sd-0.04118024800949986, 32'sd-0.1380825473345117, 32'sd0.0422993129574442, 32'sd0.06904808487903126, 32'sd0.08416560914327056, 32'sd-0.03862448088824808, 32'sd0.05913557074567975, 32'sd0.11948770921610588, 32'sd0.02352395847150254, 32'sd-0.10868625521488665, 32'sd-0.09938970018396275, 32'sd-0.05552363926066664, 32'sd-0.037035450356631514, 32'sd-0.07754193023566608, 32'sd-0.06275152812579032, 32'sd-0.06326961395245957, 32'sd-0.010665242909571713, 32'sd0.005728767621326256, 32'sd0.06304373841660013, 32'sd0.17606727710276995, 32'sd0.07934667388157225, 32'sd0.18241675848017028, 32'sd0.01735751407595442, 32'sd0.09330189608026816, 32'sd0.047922374431088134, 32'sd0.050723193977755654, 32'sd0.04996817411412558, 32'sd-0.056479367389175514, 32'sd0.019988407388956478, 32'sd-0.013552530972015751, 32'sd0.02781767035972657, 32'sd-0.05313086941985004, 32'sd-0.0026792277356056074, 32'sd-0.07362095423987185, 32'sd-0.00046088412502345687, 32'sd0.05763425962076498, 32'sd0.04722813940667721, 32'sd0.05874455599358797, 32'sd-0.005600858132774201, 32'sd0.002985431026077496, 32'sd0.0367585903756927, 32'sd0.005734205849317237, 32'sd0.007982120455631568, 32'sd-0.024855145848096828, 32'sd0.1020702202587804, 32'sd0.06533573533817429, 32'sd-0.035576434148186106, 32'sd0.002526882325978569, 32'sd-0.0809345630154515, 32'sd0.0647505472224134, 32'sd0.05077021143909615, 32'sd0.016230159068582852, 32'sd0.003911333146054996, 32'sd0.04989839109649482, 32'sd0.007666585036707363, 32'sd0.06702605138873789, 32'sd-0.041002062056608155, 32'sd-0.10057427711741582, 32'sd0.03206594482262106, 32'sd0.03400475431270375, 32'sd-0.038718889057212304, 32'sd-0.02904692456776775, 32'sd-0.024882217041807025, 32'sd0.1140586417895382, 32'sd0.09196365844103342, 32'sd0.07731298416748021, 32'sd0.06549266370420448, 32'sd0.09849884984894008, 32'sd0.02083748846627301, 32'sd0.08996214553262841, 32'sd-0.08831252144318126, 32'sd-0.01984649360847011, 32'sd0.00956755108045971, 32'sd-0.08515344380580575, 32'sd-0.04210550666886747, 32'sd-0.03014916599399449, 32'sd-0.1563903658404524, 32'sd-0.06942489766970561, 32'sd0.01183269197305093, 32'sd0.04202650863930786, 32'sd-0.005176267203386118, 32'sd-0.06190421355027791, 32'sd-0.06324432454269184, 32'sd1.4849461392762909e-05, 32'sd-0.054437575639003664, 32'sd-0.1057042360420548, 32'sd-0.023407223769106547, 32'sd0.0830218719947019, 32'sd0.01781024585888526, 32'sd0.024018322623485966, 32'sd0.09034502958571258, 32'sd0.09507993380607752, 32'sd0.16698941901071296, 32'sd0.14413339823016252, 32'sd0.19945647701565908, 32'sd0.08201412165281434, 32'sd0.16608738243223695, 32'sd0.0032663357970418093, 32'sd-0.06311052061074725, 32'sd-0.009748759024030976, 32'sd-0.052760742138282905, 32'sd-0.043642061111166655, 32'sd-0.10344385172940147, 32'sd-0.18140737611581734, 32'sd-0.05849492718525586, 32'sd-0.04757434016284295, 32'sd0.013916147329524398, 32'sd-0.014457135630027733, 32'sd0.08883098798233297, 32'sd-0.039719245342185946, 32'sd0.05066993898879957, 32'sd0.07938617892948185, 32'sd-0.013890364078683812, 32'sd0.02181162851009504, 32'sd-0.04532670962843051, 32'sd-0.044222637082516184, 32'sd0.028169087040822317, 32'sd-0.051543514559911026, 32'sd-0.03352684226635378, 32'sd0.056409537881895545, 32'sd0.2249352604051663, 32'sd0.16745688529784414, 32'sd0.25785453657494084, 32'sd0.1631837714199036, 32'sd0.10829069112156249, 32'sd0.012701947848640451, 32'sd0.04686071477181307, 32'sd0.014804321085107073, 32'sd-0.09515255055430076, 32'sd-0.1836792922915647, 32'sd-0.17405955049205593, 32'sd-0.09587963846305737, 32'sd0.00838055098920278, 32'sd-0.05955397551180642, 32'sd-0.02642976204373354, 32'sd0.024265463849182423, 32'sd0.015410023860104032, 32'sd0.04196350300083775, 32'sd-1.2959876376633807e-115, 32'sd-0.03823782118076059, 32'sd-0.05210690378840306, 32'sd-0.10648446297731222, 32'sd-0.07677504236213392, 32'sd-0.045865548049383156, 32'sd0.013199813391682785, 32'sd-0.05797771504324033, 32'sd-0.06334991731748121, 32'sd-0.11116317266144675, 32'sd0.034373147476930266, 32'sd0.05891795056262056, 32'sd0.08435775148231495, 32'sd0.1770462452430833, 32'sd0.06939175757696096, 32'sd0.16145122052517144, 32'sd-0.025723660066118245, 32'sd-0.03711420213640401, 32'sd-0.01081977449258466, 32'sd-0.22810513460689208, 32'sd-0.03494285397049082, 32'sd-0.11891054531538316, 32'sd-0.12204778345055955, 32'sd-0.14502999061436714, 32'sd0.017930552190136485, 32'sd0.0047771347132186965, 32'sd0.06020799255504277, 32'sd-0.04919845866064808, 32'sd0.031184416836009105, 32'sd-0.011748655822883567, 32'sd-0.11231098991414197, 32'sd-0.06777092173365462, 32'sd-0.1062336677638451, 32'sd-0.1487499974074966, 32'sd-0.07119217972814085, 32'sd-0.005621077849730932, 32'sd-0.045303191654348776, 32'sd-0.22069838051066365, 32'sd-0.06746064292713633, 32'sd-0.08479350853663815, 32'sd-0.08775006650083748, 32'sd0.003955878095561211, 32'sd-0.006010158020487433, 32'sd0.11515103775544297, 32'sd0.07530016329314569, 32'sd-0.0551682153493102, 32'sd-0.09501773207831891, 32'sd0.0004024274034022468, 32'sd-0.06739947500286264, 32'sd0.0018241482768356003, 32'sd-0.06386787256608772, 32'sd-0.1073940836887631, 32'sd-0.10019435033834734, 32'sd-0.01725277567865328, 32'sd0.013014723113302602, 32'sd-0.02599236126314959, 32'sd-0.009113251637129978, 32'sd-0.002738587932906517, 32'sd0.004981763433741377, 32'sd-0.0301591064766396, 32'sd-0.09931016159145467, 32'sd-0.029959395812417123, 32'sd-0.054691115258780516, 32'sd-0.08664848105231358, 32'sd-0.09771871191051959, 32'sd-0.18120845740963912, 32'sd-0.17608908464223652, 32'sd-0.0642867354353727, 32'sd-0.02556165871336583, 32'sd-0.08603609995300286, 32'sd-0.08993546407866446, 32'sd0.0843581506267047, 32'sd0.10641862695905085, 32'sd0.06788866487586766, 32'sd0.0027657489867803186, 32'sd-0.03468215665978269, 32'sd-0.028202490242473028, 32'sd0.006165682171095939, 32'sd-0.11157867663067897, 32'sd-0.12014441519384422, 32'sd0.029871621288389827, 32'sd0.004568360412676428, 32'sd0.02217664364150115, 32'sd-0.034626830922020575, 32'sd-1.1296148547707808e-114, 32'sd-0.0471748006694623, 32'sd0.054734834564686995, 32'sd-0.015499065838296288, 32'sd-0.04298135583686699, 32'sd0.07444190602435252, 32'sd0.09357069123602037, 32'sd0.01259957381481031, 32'sd-0.011444617810544828, 32'sd-0.15809843720957084, 32'sd-0.013559145670908103, 32'sd-0.04882281572325428, 32'sd-0.11026942321712084, 32'sd-0.09008238700138126, 32'sd-0.0011801482474792769, 32'sd-0.015577065392150868, 32'sd-0.019515807328427445, 32'sd0.21272063394317903, 32'sd0.08429414518328991, 32'sd0.049757270343705966, 32'sd0.004945966321515297, 32'sd0.06766235391871062, 32'sd-0.11134848285095289, 32'sd-0.06212344989470724, 32'sd-0.08028258312413936, 32'sd-0.012347241754238852, 32'sd-0.0034681913575479234, 32'sd0.03319894163553272, 32'sd0.005367667705933129, 32'sd0.004999555992022559, 32'sd0.03452143402519631, 32'sd-0.006813522428120445, 32'sd0.057721568804092946, 32'sd-0.015549914120854966, 32'sd0.0381376534566882, 32'sd0.12024755104923573, 32'sd0.03688465093570954, 32'sd0.013464879014923518, 32'sd-0.05260571278468478, 32'sd-0.07335157389759583, 32'sd-0.03317076009432451, 32'sd-0.0203477986336725, 32'sd0.001352439576356356, 32'sd0.08051674325211677, 32'sd0.005496904039250165, 32'sd0.12809653283620312, 32'sd-0.007983337718890829, 32'sd-0.04940670349248486, 32'sd-0.00842346450823681, 32'sd-0.05520666789089265, 32'sd-0.06582827995704658, 32'sd-0.0996414797983015, 32'sd-0.02576770295145386, 32'sd-0.09204970415873934, 32'sd0.011467812117913739, 32'sd0.00045398614992012186, 32'sd-0.015087134389958118, 32'sd0.026839553060196274, 32'sd-0.02544226259882357, 32'sd-0.030773338252979135, 32'sd-0.011120573059736759, 32'sd0.0010757847915736586, 32'sd0.1181550024199394, 32'sd0.11527887486317931, 32'sd0.01623744669413022, 32'sd-0.0023848323279217387, 32'sd0.0541321481522899, 32'sd0.002650677146948292, 32'sd-0.054025991395373174, 32'sd0.04464192304054735, 32'sd0.12699189866207952, 32'sd0.08101824359823759, 32'sd-0.10747926097940418, 32'sd0.016155267096606796, 32'sd-0.10513459620183041, 32'sd-0.027189581102784455, 32'sd0.003950003139409636, 32'sd-0.15374427976975652, 32'sd-0.12461663210290898, 32'sd-0.03830555610742368, 32'sd-0.03224099035712689, 32'sd-0.04604759981794439, 32'sd-0.016267236304489455, 32'sd0.055226443402009565, 32'sd-1.7257860808530014e-117, 32'sd0.03470823964413656, 32'sd0.0030252628463555485, 32'sd-0.04772643634384328, 32'sd-0.028566617747290735, 32'sd-0.03449122408515109, 32'sd-0.073003044243072, 32'sd0.07597812943690374, 32'sd0.11742048189465926, 32'sd0.06831969409700595, 32'sd-0.005598824837472753, 32'sd0.10157451744167, 32'sd0.11819297203875206, 32'sd0.11840709577947219, 32'sd-0.004216503470961259, 32'sd0.05211968212496622, 32'sd-0.05327052942977004, 32'sd-0.04480666612007253, 32'sd-0.019713581057740386, 32'sd-0.020334745646707154, 32'sd0.04421022010029978, 32'sd-0.054076764266486776, 32'sd-0.009638978881113891, 32'sd0.004018053943150214, 32'sd-0.03124362492691941, 32'sd-0.0503606231784257, 32'sd-0.03433411071515983, 32'sd-9.92062256515306e-119, 32'sd2.1256859410454823e-127, 32'sd9.754330154114338e-121, 32'sd0.010876469530667707, 32'sd-0.010836953485945742, 32'sd-0.08595821883361694, 32'sd-0.05111296407798857, 32'sd-0.022730391478125018, 32'sd0.030247498286425187, 32'sd-0.04030686492211355, 32'sd0.09096380286171607, 32'sd0.10405723848550036, 32'sd0.06800808331119162, 32'sd0.08095964729969951, 32'sd0.15090157424953854, 32'sd-0.01847984226282268, 32'sd0.059299903547745635, 32'sd0.027887898266551643, 32'sd-0.09211458939402224, 32'sd-0.09359192733816722, 32'sd-0.01064240629346919, 32'sd0.06510483077822692, 32'sd-0.039167653209241045, 32'sd-0.023918924737380172, 32'sd-0.03275345161353269, 32'sd0.051919404250121065, 32'sd-0.010299288691881126, 32'sd-0.0024230788249871957, 32'sd5.376924936502865e-118, 32'sd-1.0121607685281207e-121, 32'sd1.5148274250210466e-124, 32'sd0.10636014386615447, 32'sd0.04109702173785954, 32'sd-0.10002677223838884, 32'sd-0.09003439244077618, 32'sd-0.0040003307898088284, 32'sd0.05467776500012174, 32'sd0.01957677296279605, 32'sd0.06710636485971536, 32'sd-0.035028837403298464, 32'sd0.061717388415245336, 32'sd0.1253317128351534, 32'sd0.04268443138693751, 32'sd0.013946160140930806, 32'sd-0.05930457875135063, 32'sd-0.013977324009270617, 32'sd0.037394450313399386, 32'sd0.02606111372546715, 32'sd0.13389412178395066, 32'sd0.0011558503460218708, 32'sd0.0997354610811404, 32'sd0.03473070470777256, 32'sd0.02113211695814232, 32'sd0.018311967631361527, 32'sd-0.003233480504187347, 32'sd0.032562026829329196, 32'sd8.894534585995162e-125, 32'sd-4.733963632945428e-123, 32'sd-3.902400692266368e-119, 32'sd-1.4738239978370567e-117, 32'sd0.02266586183893608, 32'sd0.11203157550702365, 32'sd0.02575810530647755, 32'sd0.04695436316001201, 32'sd0.06175735423919435, 32'sd0.06910107502748593, 32'sd0.007405140939241198, 32'sd0.04401275228471439, 32'sd-0.06694350055011371, 32'sd0.13592501753133343, 32'sd0.15388914857422334, 32'sd0.1440197714934266, 32'sd0.02547398740351199, 32'sd0.11947937095039048, 32'sd0.06490198240546909, 32'sd0.1211349745717028, 32'sd0.07282854325688717, 32'sd0.0804319847198573, 32'sd0.02141882186200893, 32'sd0.018161299314845718, 32'sd0.10678265467639464, 32'sd-0.08338789699325758, 32'sd0.0010977346123926107, 32'sd8.01942277767532e-121, 32'sd-1.3019454798252527e-120, 32'sd5.0781610290548495e-121, 32'sd7.35671360232355e-123, 32'sd7.839302675847206e-123, 32'sd1.9766895916607885e-127, 32'sd-0.019071034646151182, 32'sd0.03514557804917832, 32'sd-0.044401186490523985, 32'sd0.023604544906329156, 32'sd-0.027139780169686042, 32'sd0.003491572263018484, 32'sd0.07950951117303287, 32'sd0.060029613186610535, 32'sd-0.005148224770258505, 32'sd0.06617552729100995, 32'sd0.09303508110098117, 32'sd0.006925723626163298, 32'sd0.04643749038216082, 32'sd0.04175172034657269, 32'sd0.04334997611567557, 32'sd0.028851232222500856, 32'sd0.007867966125812963, 32'sd-0.020077605906567885, 32'sd-0.12191676481011711, 32'sd0.014723982946604637, 32'sd1.045340429221356e-115, 32'sd9.625113759314071e-125, 32'sd4.570617869301137e-127, 32'sd6.255691745085706e-121},
        '{32'sd-1.1955744808173492e-118, 32'sd-1.3804391697612988e-120, 32'sd-9.916447130983336e-118, 32'sd7.180589079251574e-115, 32'sd2.414943554190682e-114, 32'sd-1.4150190103638153e-118, 32'sd-1.2304828608725686e-124, 32'sd-3.4209288294476295e-119, 32'sd-3.958715126010271e-119, 32'sd-1.7127331745640808e-114, 32'sd1.2003514431411635e-127, 32'sd-8.232292225653223e-121, 32'sd-0.021572345804548882, 32'sd-0.055554252457535876, 32'sd-0.03225823204307873, 32'sd-0.02783289264271017, 32'sd3.231052295357659e-121, 32'sd-1.0432739272623883e-124, 32'sd6.955040565690662e-124, 32'sd-1.8999300383565378e-126, 32'sd5.130795544265089e-118, 32'sd-2.7424038183881864e-121, 32'sd3.019306080678005e-125, 32'sd6.461688828695993e-116, 32'sd2.340977165024621e-120, 32'sd-6.806232954766468e-124, 32'sd6.969299662763265e-115, 32'sd-1.3126393713242775e-123, 32'sd6.83171852572101e-120, 32'sd-4.671379369058735e-123, 32'sd-1.8341902183719947e-121, 32'sd-1.4359786582975934e-120, 32'sd0.0056392220470043415, 32'sd-0.022661457753897933, 32'sd-0.024931978515655952, 32'sd-0.008591571915436655, 32'sd-0.033648249534237534, 32'sd-0.009638234174015166, 32'sd0.0255891387106325, 32'sd-0.06272912540372952, 32'sd-0.038997850082697, 32'sd-0.03425680864251809, 32'sd-0.08143520997523113, 32'sd-0.011996791721051288, 32'sd0.03494088733779102, 32'sd-0.02516852168222508, 32'sd0.02085309651004703, 32'sd-0.00365322963384213, 32'sd-0.0031100767303393487, 32'sd-0.02318594085133759, 32'sd0.01071033414905557, 32'sd-0.027902571756292748, 32'sd4.7363894480364625e-123, 32'sd1.3262862629314036e-122, 32'sd-2.3228060423702357e-120, 32'sd-9.983444423263993e-115, 32'sd-5.656447939907101e-117, 32'sd2.487706575555724e-121, 32'sd0.004575013870656594, 32'sd0.02771845961489405, 32'sd-0.0005053877699067236, 32'sd-0.023397665022222066, 32'sd0.04239764853940213, 32'sd0.06209759749186782, 32'sd-0.04850704962447961, 32'sd-0.0643193985441612, 32'sd0.05182945342654078, 32'sd-0.06880086897918065, 32'sd-0.11024453376654178, 32'sd0.014135593300335245, 32'sd0.03916000389852444, 32'sd-0.01540546793185683, 32'sd-0.09212149016263754, 32'sd0.00753667934485744, 32'sd-0.05516298782285486, 32'sd-0.129776973121089, 32'sd-0.07010199332292982, 32'sd0.011199659089549618, 32'sd0.0208356773506744, 32'sd-0.05844879819254225, 32'sd0.023704384542022228, 32'sd0.0419227530926517, 32'sd-3.771120462680514e-125, 32'sd-6.886103398787263e-124, 32'sd-4.0471054882283156e-115, 32'sd5.365594112563531e-118, 32'sd-0.05274478650412983, 32'sd-0.057695688702572134, 32'sd0.028226342773217162, 32'sd-0.07970320691355672, 32'sd-0.027361194124086993, 32'sd-0.004844696188103539, 32'sd0.03139454973196645, 32'sd-0.08103502632604526, 32'sd0.0132023996340131, 32'sd0.0019012401623633628, 32'sd-0.06640462398231278, 32'sd-0.0999438129371344, 32'sd-0.07757120652895669, 32'sd-0.05801929665293444, 32'sd-0.10088581458601856, 32'sd-0.17502541491607246, 32'sd-0.07151684756891356, 32'sd-0.18571840419300192, 32'sd-0.04777048559957049, 32'sd-0.1138523961363644, 32'sd-0.01682282193690348, 32'sd0.04952754861656518, 32'sd0.05882755205112101, 32'sd0.044292474263104675, 32'sd-0.008937418609133295, 32'sd2.723975313524344e-120, 32'sd-2.5950200290828704e-122, 32'sd0.004222870896725373, 32'sd-0.015989191725265254, 32'sd0.04148241022572628, 32'sd0.07183918770561493, 32'sd0.012365632847531177, 32'sd-0.050757367084419955, 32'sd0.05776864195683441, 32'sd0.02805934919670736, 32'sd-0.03139836874672836, 32'sd-0.014049202545450478, 32'sd0.04601786673718417, 32'sd0.06750814444639668, 32'sd0.13228358519466477, 32'sd-0.06415646049217673, 32'sd-0.0337492965086409, 32'sd-0.032205309608602684, 32'sd-0.0754985891213367, 32'sd-0.15922780141128454, 32'sd-0.0740985007765182, 32'sd-0.17259071159506548, 32'sd-0.04352046601534031, 32'sd-0.009883881215270595, 32'sd-0.061632726575647306, 32'sd0.008435358280963966, 32'sd-0.04099342780538936, 32'sd-0.017475018736449924, 32'sd-0.028144900719496824, 32'sd-1.6321640286610192e-115, 32'sd-0.0010442924493294214, 32'sd0.00301955745239848, 32'sd0.06416435553012556, 32'sd0.07103921634970312, 32'sd0.06537277093159427, 32'sd0.008574028252800778, 32'sd0.09228150688880946, 32'sd-0.008373994281468749, 32'sd-0.00038673031225471536, 32'sd0.055023199990273, 32'sd0.0064927151973551795, 32'sd0.05222852234981384, 32'sd-0.012516860848349567, 32'sd-0.03318895464966532, 32'sd0.0225615398288152, 32'sd-0.09801749453269945, 32'sd-0.18197216673344355, 32'sd-0.1335699703958091, 32'sd-0.13097910183526557, 32'sd-0.14044355445670362, 32'sd-0.18005074854411754, 32'sd-0.054420223931717, 32'sd0.09421677804779917, 32'sd-0.11652850299246527, 32'sd0.041262016062238505, 32'sd-0.06465830705821424, 32'sd-0.043044493604933606, 32'sd2.036790181250002e-122, 32'sd0.048298485423030384, 32'sd0.005566592307255407, 32'sd0.015956755748988624, 32'sd0.04443241244331067, 32'sd0.051725296332309156, 32'sd0.03192152464206141, 32'sd0.05913259794135315, 32'sd0.05959018079830054, 32'sd0.09092100425956127, 32'sd0.11272651979527652, 32'sd0.053452192985639545, 32'sd-0.029169945202159292, 32'sd0.06101926023505599, 32'sd0.05606894218701604, 32'sd0.07856479448217821, 32'sd-0.07144021739081984, 32'sd-0.01944720802348173, 32'sd-0.01699304494676619, 32'sd-0.07767832197122444, 32'sd-0.07528403994743521, 32'sd-0.01692689062731975, 32'sd0.05992666654255349, 32'sd-0.06566958839770647, 32'sd-0.09094006003976109, 32'sd-0.11536280569029189, 32'sd0.075626560169924, 32'sd-0.08235328819284247, 32'sd-0.016711101436696067, 32'sd-0.06252527404895133, 32'sd0.0014967764712788077, 32'sd0.04395410951400593, 32'sd0.10935080257402328, 32'sd0.0496087670960993, 32'sd0.08495036641849939, 32'sd0.06531978973801043, 32'sd0.08337542712140689, 32'sd0.0050382773549876815, 32'sd0.0008882300233677816, 32'sd-0.06487197856915737, 32'sd0.08087051457467316, 32'sd0.026972380701138, 32'sd0.1630223128795201, 32'sd0.004209530464385776, 32'sd0.046558711089366586, 32'sd-0.06271194874166991, 32'sd-0.06050537537068178, 32'sd-0.05713962299999836, 32'sd-0.04594103743031526, 32'sd-0.09289100632500809, 32'sd-0.1005698278354333, 32'sd-0.1313362994899493, 32'sd-0.02446120703841636, 32'sd0.06806588325968363, 32'sd0.050997580215551834, 32'sd0.02282353331347236, 32'sd0.03894259765456485, 32'sd-0.047196144384504694, 32'sd-0.056962397521676374, 32'sd-0.02018623296475663, 32'sd0.10445940981085189, 32'sd0.09746694442139854, 32'sd0.0003075321300619397, 32'sd-0.13864087880259873, 32'sd0.11697912971912616, 32'sd-0.027704240312973544, 32'sd0.04440603185416801, 32'sd0.04017341699508634, 32'sd-0.04007096104153329, 32'sd0.12283235082382311, 32'sd0.03789327191665708, 32'sd-0.006413602741766383, 32'sd-0.05157539306574688, 32'sd0.008328773828110083, 32'sd-0.02741265456902599, 32'sd-0.004348992254846799, 32'sd-0.05450749434699881, 32'sd-0.08405857444752865, 32'sd0.006116378246795931, 32'sd0.01087349606995898, 32'sd-0.05157347084712041, 32'sd0.08522387184249788, 32'sd-0.005462315216737888, 32'sd-0.08326403663297982, 32'sd0.0631174483261221, 32'sd-0.05211256575659616, 32'sd0.068871660840864, 32'sd-0.008223004217152363, 32'sd-0.007360601371473638, 32'sd-0.017057849890296618, 32'sd-0.10831064907497215, 32'sd0.01961921905963963, 32'sd0.00430789354533718, 32'sd0.008170031827495572, 32'sd-0.02046827431692502, 32'sd-0.02795202855153075, 32'sd0.1071876472826232, 32'sd0.19926967844572127, 32'sd0.22664560247050142, 32'sd0.10897945450241663, 32'sd-0.06907569669221593, 32'sd-0.09636523002307544, 32'sd-0.12365332112283141, 32'sd-0.02183454601758391, 32'sd-0.06335685100306442, 32'sd0.040009326429542476, 32'sd0.09813195987017426, 32'sd0.06550830021611703, 32'sd-0.00010111875518939004, 32'sd-0.012673050259769213, 32'sd0.022118288806313433, 32'sd0.018554206358822857, 32'sd0.020053309360077255, 32'sd-0.011455806164264387, 32'sd-0.014098970945323587, 32'sd0.07562955330443735, 32'sd-0.0791511094923276, 32'sd-0.05891515822377239, 32'sd-0.09646694920977408, 32'sd0.04141478970221798, 32'sd-0.04369062031474589, 32'sd-0.12560029115674792, 32'sd-0.07921959534154052, 32'sd0.12861391568775948, 32'sd0.03076196457081126, 32'sd0.12970811233451437, 32'sd0.07755178940136445, 32'sd-0.039407349953467063, 32'sd-0.05282309121374915, 32'sd-0.09539645514150727, 32'sd-0.05011654310117772, 32'sd-0.08694847695020044, 32'sd0.08476455651757844, 32'sd0.06741992599984938, 32'sd-0.031728012770617244, 32'sd0.13344172906034385, 32'sd0.07090360716727086, 32'sd-0.02415484626363595, 32'sd0.017648717412297083, 32'sd0.07661612119980109, 32'sd-0.042219472018095346, 32'sd-0.08216751649470423, 32'sd0.017903041075955986, 32'sd0.13482922202387113, 32'sd-0.01870909891780536, 32'sd-0.07298911431632979, 32'sd-0.0056745635514829085, 32'sd0.009210381692851153, 32'sd0.014030563974687871, 32'sd-0.09110927620527112, 32'sd0.0956529641221046, 32'sd0.04496704411619266, 32'sd-0.08219339296982194, 32'sd-0.02597784829640566, 32'sd0.009106198968833466, 32'sd-0.05753538820340409, 32'sd-0.07713204774644589, 32'sd-0.03633906092269658, 32'sd-0.08239375263253713, 32'sd0.004182120399482431, 32'sd0.11757246999311638, 32'sd0.04164574733028641, 32'sd-0.03817145707383743, 32'sd0.025558753615321436, 32'sd-0.133384095412877, 32'sd0.04948999096167033, 32'sd0.03228957837544927, 32'sd0.011252348693576254, 32'sd0.029401853792565765, 32'sd-0.025861166811603088, 32'sd0.013657370590257477, 32'sd0.02132686422935735, 32'sd0.048783571902247976, 32'sd-0.01694176589613485, 32'sd0.07349913341536314, 32'sd-0.12209024222050342, 32'sd0.013805224983007817, 32'sd-0.01705613467108978, 32'sd-0.019773877535699758, 32'sd-0.12797348149399435, 32'sd-0.26034923996627884, 32'sd-0.06571634990114253, 32'sd0.035128563276758486, 32'sd0.012625288205076675, 32'sd0.0033184691316355086, 32'sd0.011689062461928091, 32'sd0.05056285183294392, 32'sd0.05250187397489579, 32'sd0.11831930755584243, 32'sd0.01867210811297949, 32'sd-0.0626677301991041, 32'sd0.021743522473163426, 32'sd-0.0061776441975027645, 32'sd0.02960641034327396, 32'sd-0.0700584845364063, 32'sd-0.026700537408158392, 32'sd-0.01699892514931671, 32'sd0.08317381209332465, 32'sd0.07504131559833219, 32'sd0.06639804270331395, 32'sd-0.08508432319942548, 32'sd-0.09570618058606807, 32'sd0.10402253029640927, 32'sd-0.05320520378398339, 32'sd-0.033438525397232036, 32'sd0.010648274601181533, 32'sd-0.1513927477415977, 32'sd-0.20430597616694346, 32'sd-0.14226661625497344, 32'sd0.026223402966764765, 32'sd0.19469297315883688, 32'sd0.12369083901059054, 32'sd0.0896559460263394, 32'sd0.1582480755836737, 32'sd0.17801286704209704, 32'sd0.030208373516253918, 32'sd0.007489383986178762, 32'sd-0.028317327516570075, 32'sd-0.0893551119598063, 32'sd-0.019911871626176858, 32'sd-0.04487579541994053, 32'sd0.009637801655055091, 32'sd-0.034892401087940575, 32'sd-0.022431111061500596, 32'sd-0.026286450102007194, 32'sd-0.045270644295169284, 32'sd0.09999419791505058, 32'sd-0.16028847162851456, 32'sd-0.047579213948432675, 32'sd-0.0961973662607338, 32'sd-0.10429071819281122, 32'sd0.08434463950587334, 32'sd-0.02155949714116666, 32'sd-0.12590706019239412, 32'sd-0.22962402613777774, 32'sd-0.05093286286595222, 32'sd0.11149251112437128, 32'sd0.1265519454325897, 32'sd0.20393740041261235, 32'sd0.19771813570469352, 32'sd0.14983441656018842, 32'sd0.14095351945529397, 32'sd0.016731743825372625, 32'sd0.050317147137524686, 32'sd-0.002405593318248919, 32'sd0.05057595183454154, 32'sd-0.16248382932441152, 32'sd-0.07199749707340382, 32'sd0.011357795257052758, 32'sd0.010981509947297411, 32'sd0.1357841623511353, 32'sd0.027440534990327423, 32'sd-0.05057851635039226, 32'sd0.06418010535807424, 32'sd0.051926819531810706, 32'sd-0.049803853808887716, 32'sd-0.11867271476715295, 32'sd0.0244799555832128, 32'sd-0.030043731830770075, 32'sd-0.11705052452268826, 32'sd-0.12757259701437149, 32'sd-0.17903023918196292, 32'sd-0.08344327842076847, 32'sd-0.0553024980177803, 32'sd0.09710454614343982, 32'sd0.20983981633407334, 32'sd0.2622227313314183, 32'sd0.07448995204489128, 32'sd0.23535597928589364, 32'sd0.13442793290809296, 32'sd-0.07423641447291615, 32'sd0.020629467070648628, 32'sd0.1357053926749871, 32'sd-0.02927492197373988, 32'sd-0.12304977519408025, 32'sd-0.04271105402188148, 32'sd-0.08578870572008732, 32'sd0.03279151960399162, 32'sd0.06709114596818375, 32'sd0.06741163451372546, 32'sd0.003365248632647989, 32'sd-0.05648466956607961, 32'sd0.03810208982675434, 32'sd0.038347771162403954, 32'sd0.11164899684217304, 32'sd0.05493139213587072, 32'sd-0.05851638614946224, 32'sd0.07628783042739622, 32'sd-0.1000319104947971, 32'sd0.020883696952173986, 32'sd0.03435742319051008, 32'sd7.797124053179957e-05, 32'sd0.21385107460367422, 32'sd0.23795282634660522, 32'sd0.08462955872960669, 32'sd0.022176421769164633, 32'sd0.00544862521697099, 32'sd-0.07289025559283321, 32'sd-0.008561125399150887, 32'sd-0.005290717683355978, 32'sd0.04620026407307749, 32'sd0.04383163290563535, 32'sd-0.030334058688393683, 32'sd-0.08098677935016621, 32'sd0.010310528976099473, 32'sd-0.007279203443317541, 32'sd-0.0211392107579285, 32'sd-0.02945610861816702, 32'sd2.5617255308778784e-124, 32'sd0.058276975350197456, 32'sd-0.05709198137080968, 32'sd0.0538227689449882, 32'sd0.0922952759756032, 32'sd0.09907579151983734, 32'sd-0.029269541012803803, 32'sd-0.02292719364269648, 32'sd-0.010165625156131541, 32'sd-0.13595944619941136, 32'sd-0.12157918641543211, 32'sd-0.07891341289953727, 32'sd0.10603644046036789, 32'sd0.0168792052951173, 32'sd0.004916045521696785, 32'sd-0.02065477351470072, 32'sd-0.14887867134181365, 32'sd-0.12351781934656013, 32'sd-0.16015711934946858, 32'sd-0.042411969638642036, 32'sd0.028432367499006232, 32'sd-0.043024242865041876, 32'sd-0.16674431069777285, 32'sd-0.06759077801506688, 32'sd0.03465720636894591, 32'sd0.03695647876671835, 32'sd0.03376299573595385, 32'sd0.009689245520427487, 32'sd-0.06874054700739454, 32'sd-0.010355432731879565, 32'sd0.06367838625006454, 32'sd-0.08915508944360842, 32'sd0.08480475656542268, 32'sd0.04432309703342911, 32'sd-0.07061197478104371, 32'sd-0.05616104167846706, 32'sd-0.12799369234441352, 32'sd-0.12791821078918264, 32'sd-0.15967751795546073, 32'sd-0.03979080487781513, 32'sd-0.04902360379630953, 32'sd-0.0772246715440518, 32'sd-0.09526507709121491, 32'sd-0.10639515803966114, 32'sd-0.03576816689641336, 32'sd-0.1267274524755362, 32'sd-0.07313051455585243, 32'sd-0.07272613656003822, 32'sd-0.04022875234492863, 32'sd-0.04739568247371982, 32'sd-0.0636221965551498, 32'sd0.014740474855041699, 32'sd-0.07097117944601487, 32'sd-0.08179688720808546, 32'sd-0.10881877255842237, 32'sd-0.07807774406123562, 32'sd-0.002717986968880663, 32'sd0.03991268336332833, 32'sd-0.03195893787809609, 32'sd-0.07640403667240046, 32'sd0.09437839988793528, 32'sd0.02563964580832639, 32'sd-0.08601742671889417, 32'sd-0.1401019379208356, 32'sd-0.0565163189773203, 32'sd-0.0191979918843613, 32'sd0.03346142856509628, 32'sd-0.16044012319445808, 32'sd-0.19418371859871977, 32'sd-0.1577812563789415, 32'sd-0.07529762399703428, 32'sd-0.11408102076337391, 32'sd0.05453701486984799, 32'sd-0.08326813355418337, 32'sd-0.036792386052726035, 32'sd-0.014542973982399869, 32'sd-0.060623518978337086, 32'sd0.03995040055963938, 32'sd-0.04977523472692724, 32'sd0.005005872224392512, 32'sd-0.03238802228742794, 32'sd0.04482271815863417, 32'sd-0.09029207651063088, 32'sd0.010237539311732931, 32'sd3.3282919722932196e-121, 32'sd0.05061110906094285, 32'sd-0.01890042152715869, 32'sd0.07546462878802712, 32'sd-0.02420435111915727, 32'sd-0.022543653430561673, 32'sd0.027156307978342047, 32'sd0.04726604736803303, 32'sd-0.023020643544472152, 32'sd0.0015076085884379318, 32'sd-0.13330084718292018, 32'sd-0.10213620422267336, 32'sd-0.058324290913774404, 32'sd-0.08464962376625311, 32'sd0.037875985705142244, 32'sd-0.0948005218136928, 32'sd-0.11600562634087351, 32'sd0.012933787335545678, 32'sd0.06758804767535079, 32'sd0.0004434737533266688, 32'sd0.03263661723405159, 32'sd0.023945156219908396, 32'sd-0.022124527238974668, 32'sd-0.018634938422106707, 32'sd-0.07960357507690581, 32'sd-0.027550223289608683, 32'sd-0.04800682576218368, 32'sd-0.02812016696883314, 32'sd-0.002683241435997796, 32'sd0.04906957120879677, 32'sd-0.05775373520379008, 32'sd0.06754337732373324, 32'sd0.07591278639724529, 32'sd0.120541652577073, 32'sd0.06952917166821104, 32'sd0.06233221414836981, 32'sd0.015236628536518299, 32'sd-0.04615423205530468, 32'sd0.06634618697887858, 32'sd-0.006530279457997609, 32'sd-0.09866726945889381, 32'sd-0.08814701978799976, 32'sd-0.09848850614493344, 32'sd-0.10623615820648172, 32'sd-0.056356290681823566, 32'sd-0.17769315123843235, 32'sd-0.003871537733929642, 32'sd-0.02704497921626529, 32'sd0.03372130944367383, 32'sd-0.07284358048270434, 32'sd-0.06569810562369272, 32'sd-0.0880524155638189, 32'sd-0.1189148803187128, 32'sd-0.0028966748150178806, 32'sd-0.053819304202655814, 32'sd0.07062044910291063, 32'sd-0.026444147946509105, 32'sd0.03173760173987478, 32'sd-0.028942417257638405, 32'sd-0.03325858717418375, 32'sd0.1094160891583452, 32'sd-0.006215457050188997, 32'sd-0.03415528242364407, 32'sd0.05361183549626118, 32'sd0.038497760945668966, 32'sd0.03274888227565472, 32'sd0.007442412217584212, 32'sd-0.10882220932627186, 32'sd-0.024089824266107847, 32'sd-0.040269129132263715, 32'sd0.012474629850425656, 32'sd-0.029777290065588127, 32'sd-0.12010038271715798, 32'sd-0.04234406745063573, 32'sd0.0855919905647103, 32'sd-0.03540404885772595, 32'sd-0.03168147853686104, 32'sd-0.03415467278464997, 32'sd0.026524418805960376, 32'sd-0.08978320725860686, 32'sd0.04907853174222997, 32'sd0.023666468596151586, 32'sd0.04355215547553765, 32'sd0.04660005162216589, 32'sd3.9416820497382416e-119, 32'sd-0.03162074241243593, 32'sd0.02133970783233417, 32'sd0.020296718856906353, 32'sd0.017872727957277987, 32'sd0.044250013101482216, 32'sd0.014387150604078584, 32'sd0.08415189306070434, 32'sd-0.03570047798757759, 32'sd0.02675039341863039, 32'sd-0.05694691321876635, 32'sd-0.056256979822771225, 32'sd0.03250384716073122, 32'sd-0.05334406057482201, 32'sd0.04408376752848541, 32'sd0.05795790568073307, 32'sd-0.028162524848963554, 32'sd-0.03011173007577399, 32'sd0.029530322885534328, 32'sd-0.037605076174052524, 32'sd-0.08865289416046601, 32'sd-0.012270946806135254, 32'sd-0.014189611019830307, 32'sd-0.10687443976918104, 32'sd0.07910971524909792, 32'sd-0.02657693760248451, 32'sd0.07762251418426, 32'sd-3.6047508620751234e-121, 32'sd-5.388553531568572e-118, 32'sd-1.1101260976900462e-121, 32'sd-0.06867412619711652, 32'sd0.024110391656742756, 32'sd-0.0718764319412464, 32'sd0.0114056744775159, 32'sd0.048993681416773995, 32'sd-0.005013911950817165, 32'sd-0.02146885643355341, 32'sd-0.06139852115309946, 32'sd0.0449523235244735, 32'sd-0.04956678077016706, 32'sd-0.16043011628640205, 32'sd-0.025468788516019053, 32'sd0.048901852951714606, 32'sd-0.03729552239611433, 32'sd0.00010202242479346469, 32'sd0.08236636807466005, 32'sd0.12306885455546109, 32'sd0.07552096077689034, 32'sd0.09349703972224738, 32'sd0.005544492180077568, 32'sd0.009968933266875101, 32'sd-0.11879061765854171, 32'sd0.009143803698805044, 32'sd-0.06965828186159713, 32'sd0.05329657509541011, 32'sd8.324021439169438e-125, 32'sd-2.0156091589365606e-124, 32'sd-2.286896949602678e-120, 32'sd0.09046656989907045, 32'sd0.01971540671128419, 32'sd0.001970566793371286, 32'sd0.13084604832697738, 32'sd-0.03414991104879145, 32'sd0.13756632094630014, 32'sd0.10295804584096273, 32'sd0.051291063662356584, 32'sd-0.03692283202651646, 32'sd-0.03690536594125955, 32'sd-0.042069093584375335, 32'sd0.07734047539069355, 32'sd0.04203277387937235, 32'sd-0.05571315032762498, 32'sd-0.008749771044331058, 32'sd-0.007739558843611237, 32'sd-0.07893395374245206, 32'sd-0.044531750810158484, 32'sd0.05019987214857459, 32'sd0.09793736781152651, 32'sd-0.0516316662157678, 32'sd0.03297438481389421, 32'sd-0.028035941011842543, 32'sd-0.0063205564676828115, 32'sd0.02160509781869719, 32'sd1.9071383675381928e-126, 32'sd1.50982617252327e-124, 32'sd1.4021392413058092e-124, 32'sd-1.8674884669266492e-126, 32'sd0.031946459719862895, 32'sd0.10305563879975832, 32'sd0.0926417035707672, 32'sd-0.013973178469875778, 32'sd0.1769673405056412, 32'sd0.0460777758033736, 32'sd0.10963125686406577, 32'sd0.052013567526027385, 32'sd0.09735084224018008, 32'sd0.08534178622306594, 32'sd-0.020158955631023087, 32'sd-0.008306983861876293, 32'sd-0.11994179629830393, 32'sd-0.02248170692047495, 32'sd0.045971087008088746, 32'sd-0.04453322952156389, 32'sd-0.02283191677866022, 32'sd0.031550527758592066, 32'sd0.05418031086468865, 32'sd0.03155148757506733, 32'sd-0.001234236367773196, 32'sd-0.051446773173535035, 32'sd0.0028766610726325328, 32'sd-2.71604688378167e-124, 32'sd-2.6746779047193187e-125, 32'sd1.1958497743541823e-117, 32'sd6.38316119029028e-117, 32'sd-3.1727220195552284e-121, 32'sd7.285807243013368e-122, 32'sd0.04354825251297372, 32'sd-0.022758770382038516, 32'sd-0.036581319867661874, 32'sd-0.009144743141209402, 32'sd0.005545134177004634, 32'sd-0.04613134100763993, 32'sd0.07699604213997675, 32'sd-0.03632054359845549, 32'sd0.06093569411933077, 32'sd-0.005230565024819841, 32'sd0.10697806456853187, 32'sd-0.017694350180687768, 32'sd-0.006969087536975582, 32'sd0.04821396732730659, 32'sd0.04949587721256558, 32'sd-0.08846822605296503, 32'sd0.049267343890896875, 32'sd-0.046348348365921097, 32'sd-0.08551608862797486, 32'sd-0.011030797812073993, 32'sd-1.0463732211414846e-120, 32'sd-7.554149086045057e-115, 32'sd1.1737099278256256e-118, 32'sd3.277024466530463e-125},
        '{32'sd3.3470534275471847e-128, 32'sd-1.8037464127818962e-121, 32'sd-6.532412508067952e-121, 32'sd-4.0325523454031266e-127, 32'sd2.0654722091186685e-127, 32'sd-1.8665585135427824e-126, 32'sd2.206710674673478e-124, 32'sd-5.523830824378826e-115, 32'sd5.7817824788173924e-126, 32'sd-8.21411910919725e-128, 32'sd3.3795344826398094e-125, 32'sd1.0945595504042873e-115, 32'sd-0.00495094678980464, 32'sd0.06689092435182675, 32'sd0.04307101980900563, 32'sd0.10722185120621369, 32'sd3.875429627845417e-117, 32'sd-3.3395774384709175e-123, 32'sd1.32731017008827e-126, 32'sd3.4336973631302216e-125, 32'sd5.3467434000394575e-121, 32'sd9.23191745280038e-124, 32'sd-7.677331993476898e-125, 32'sd-2.431455642771972e-120, 32'sd4.8924823365147955e-115, 32'sd9.418355075550487e-120, 32'sd-3.704627027290137e-123, 32'sd-4.536229030794485e-127, 32'sd8.16548114764692e-127, 32'sd1.0779616964630822e-124, 32'sd9.680371466958613e-122, 32'sd2.0531279501420537e-121, 32'sd0.04318319323414228, 32'sd-0.008541567192018358, 32'sd-0.03295716615064897, 32'sd-0.054894872549347676, 32'sd-0.06278067877740223, 32'sd-0.0385921690802835, 32'sd0.04244497175378259, 32'sd0.10150260559660226, 32'sd-0.036387385454678726, 32'sd-0.022001816538022568, 32'sd-0.028568743308476745, 32'sd0.07714180901526717, 32'sd0.0379167820077881, 32'sd0.046694470025781476, 32'sd-0.04947830695716888, 32'sd-0.016273519136542132, 32'sd0.06518194192311694, 32'sd0.06746027200398634, 32'sd-0.06675771861444099, 32'sd0.08162277044878108, 32'sd-6.4318249306844065e-124, 32'sd7.9395034218318e-122, 32'sd-3.4319897862650522e-121, 32'sd-3.0563359230871525e-120, 32'sd-4.1984343911059805e-118, 32'sd-2.0614110062825848e-116, 32'sd0.08688532248955971, 32'sd-0.016276092452576326, 32'sd-0.093306251496852, 32'sd0.010966925527511018, 32'sd-0.01222773908232416, 32'sd0.0456559643736943, 32'sd0.028330425421851588, 32'sd0.0027748268172919357, 32'sd0.14599263713073923, 32'sd0.04645282549331277, 32'sd0.04277733431328815, 32'sd0.027108991283186532, 32'sd0.045243431126946065, 32'sd0.04200533407522044, 32'sd0.1174949154544889, 32'sd-0.007077187701108821, 32'sd0.05796596175222605, 32'sd0.13872544094759992, 32'sd0.1240958042892906, 32'sd0.033685976652896035, 32'sd0.01310892004068219, 32'sd-0.057349988863480424, 32'sd0.0687491239544077, 32'sd0.05540522585222774, 32'sd2.675897828644405e-122, 32'sd1.9996267516710336e-116, 32'sd9.78071704945996e-121, 32'sd3.327569992469291e-122, 32'sd-0.05849692657021756, 32'sd0.021777541769064154, 32'sd0.07184506108361892, 32'sd0.025928631991473352, 32'sd0.07033217820180225, 32'sd0.04637936298796525, 32'sd0.009555459492075188, 32'sd0.0619533945187174, 32'sd-0.002682761676255712, 32'sd0.0008420569115231725, 32'sd0.07206891883827028, 32'sd0.020107674409521034, 32'sd-0.019523598278160016, 32'sd0.1270210292364665, 32'sd0.008089174396592637, 32'sd0.05002210844256945, 32'sd0.2326159824551825, 32'sd0.12985851374535617, 32'sd-0.04311289763358721, 32'sd0.053590676230539945, 32'sd0.13880022637640416, 32'sd0.01699802222412285, 32'sd0.05329479754384074, 32'sd0.032552061206827264, 32'sd0.013045443283428451, 32'sd1.3032158504117787e-118, 32'sd8.424609692380856e-123, 32'sd0.011952804683166946, 32'sd0.04620011579377956, 32'sd0.08957797501654152, 32'sd0.006927452510458702, 32'sd-0.04189446716129335, 32'sd0.035833180184132785, 32'sd-0.00020701362822057547, 32'sd0.1315539283043283, 32'sd0.06719185994900904, 32'sd0.08213978499011962, 32'sd0.014933798238910393, 32'sd0.010706372299833834, 32'sd0.09035529879580254, 32'sd-0.016834286440489257, 32'sd0.09491493258682787, 32'sd0.12629088451249212, 32'sd0.052087407622554156, 32'sd0.14453185509033778, 32'sd0.10519076022997426, 32'sd0.02934871562306065, 32'sd0.08058676103303727, 32'sd-0.02060581625262678, 32'sd-0.1620210796738838, 32'sd0.047301033287455024, 32'sd0.07839544278880517, 32'sd-0.029346028080136952, 32'sd0.03493065625735789, 32'sd1.2582357217735849e-123, 32'sd0.07739201982354599, 32'sd0.06580509017244537, 32'sd0.07669123253467511, 32'sd-0.04320277341227935, 32'sd0.14373707390570895, 32'sd-0.01757724929675501, 32'sd0.03832988879220393, 32'sd0.11217832226867884, 32'sd0.12616160621763345, 32'sd0.11280484995936946, 32'sd-0.04136073069654129, 32'sd-0.06404101242928832, 32'sd-0.003804851471545228, 32'sd-0.018340483729553637, 32'sd0.037022260637959416, 32'sd0.05230146661682794, 32'sd0.06754064589416531, 32'sd0.20176431690397417, 32'sd0.01686956197043422, 32'sd0.08874637850248818, 32'sd0.012441686121424274, 32'sd0.005508219312905642, 32'sd0.10422907660410102, 32'sd0.06351641813547974, 32'sd-0.05541818405863719, 32'sd-0.08133670144720855, 32'sd0.024139986840033566, 32'sd-1.189923547692493e-117, 32'sd0.022955961032251396, 32'sd0.018559253250244788, 32'sd0.05560693798868685, 32'sd0.01969579750380952, 32'sd-0.044288108989984296, 32'sd-0.007247139150669879, 32'sd0.08809746623587329, 32'sd0.03883687294257065, 32'sd0.15733582525591985, 32'sd0.1991604310921123, 32'sd0.006570932721419685, 32'sd0.08893247313989842, 32'sd0.07182757021032879, 32'sd0.047967005602295686, 32'sd0.08878340949351356, 32'sd-0.03835124565043107, 32'sd-0.03314615448494581, 32'sd0.059948769031084446, 32'sd0.10803209130099008, 32'sd-0.05064874929248539, 32'sd0.05475567432137409, 32'sd0.039794878753253306, 32'sd-0.027623098666307393, 32'sd0.03455028014216979, 32'sd0.042567604004264056, 32'sd0.0482923358952249, 32'sd-0.08086037112535623, 32'sd0.09014058644521616, 32'sd0.06446611669261766, 32'sd0.0018283917902867713, 32'sd0.08124234065956472, 32'sd-0.010643166790937918, 32'sd-0.07170283579809064, 32'sd-0.004826294150058411, 32'sd0.026576682871737804, 32'sd-5.979812382837525e-05, 32'sd0.01847632797634954, 32'sd0.02529227200701314, 32'sd0.01302986015631534, 32'sd0.04312368916518459, 32'sd0.055228489298218324, 32'sd0.07399228634577704, 32'sd-0.035205759327434485, 32'sd0.011837689460819303, 32'sd0.048545801272010254, 32'sd0.07477410142837364, 32'sd0.1789496211519148, 32'sd0.056337683122264295, 32'sd0.13502944589622992, 32'sd0.03232078175330806, 32'sd0.11911888900918353, 32'sd-0.05484132888358493, 32'sd0.10349504480171255, 32'sd0.007405115832871316, 32'sd0.04579542559021221, 32'sd0.038801640738630856, 32'sd0.051846551050657774, 32'sd0.024504494337360194, 32'sd-0.014575107433661843, 32'sd-0.0024962156380128305, 32'sd-0.02451842251507084, 32'sd-0.057189060927889654, 32'sd0.04817366852800772, 32'sd-0.0662192305358108, 32'sd-0.04623693040754164, 32'sd-0.0716130380500961, 32'sd-0.04067847665773702, 32'sd0.007725854353174432, 32'sd-0.09402526033312956, 32'sd-0.0963082813408768, 32'sd-0.07817357465265719, 32'sd0.06540285130313768, 32'sd0.10701867792083437, 32'sd0.011627921441326159, 32'sd0.21903595328491185, 32'sd0.006456449105814875, 32'sd0.041677500875199634, 32'sd-0.005647462762541056, 32'sd0.0052691225005066945, 32'sd-0.037577145832706826, 32'sd0.008626415516545518, 32'sd0.1328300829213088, 32'sd0.06591301995123491, 32'sd-0.009407869958302749, 32'sd-0.02801231673685134, 32'sd-0.05878693363466722, 32'sd0.04221779564316285, 32'sd0.08118788809137308, 32'sd0.005735153421752521, 32'sd0.046115118688876855, 32'sd0.023784484842811912, 32'sd-0.028734222327267845, 32'sd0.0015089468166861954, 32'sd-0.09168058676949481, 32'sd-0.21685952972287006, 32'sd-0.12969051449849744, 32'sd-0.20102006570631048, 32'sd-0.2531333093475911, 32'sd-0.16566816805158244, 32'sd0.04746948707583832, 32'sd0.18887090537801296, 32'sd0.03742175102552839, 32'sd0.08999888895074366, 32'sd-0.03291740017098026, 32'sd-0.10919411707205136, 32'sd0.06480116163851973, 32'sd0.025646123292180772, 32'sd-0.12005095549394472, 32'sd-0.0604520559137555, 32'sd-0.0038076676390656045, 32'sd0.03192177882960009, 32'sd0.05230460532464053, 32'sd0.01035856349783797, 32'sd0.0378148021778552, 32'sd0.05114932434890153, 32'sd0.10496246890886483, 32'sd-0.15952519001667706, 32'sd-0.10277481731346748, 32'sd-0.18848355097248384, 32'sd-0.0526951037317315, 32'sd-0.09149678928548823, 32'sd-0.26522487603221956, 32'sd-0.30093137884505894, 32'sd-0.22860439568231425, 32'sd-0.3420031366228468, 32'sd-0.26567427180394004, 32'sd-0.17332083413966348, 32'sd0.21628831048359676, 32'sd0.15002565762141468, 32'sd0.0412681719279732, 32'sd0.0949402200164214, 32'sd-0.03320195534735397, 32'sd-0.04467397640274788, 32'sd0.009831063880737432, 32'sd-0.08715355169586068, 32'sd-0.04615120599134783, 32'sd0.02441584299741593, 32'sd0.08686973380885282, 32'sd0.04394597984136144, 32'sd-0.014912867835736242, 32'sd-0.044846075398327974, 32'sd0.03193647351289634, 32'sd-0.009290776010080489, 32'sd-0.07831905995213029, 32'sd-0.14676807306739587, 32'sd-0.1456655503657011, 32'sd-0.2205972816202038, 32'sd-0.2842230107567359, 32'sd-0.2361770942661458, 32'sd-0.2178545486447721, 32'sd-0.250791075001889, 32'sd-0.16457355337993787, 32'sd-0.2316704448421733, 32'sd-0.22793568532391045, 32'sd-0.020848991715874194, 32'sd0.1443263927535078, 32'sd0.09340342050618931, 32'sd0.09377814403137097, 32'sd0.05807577755629129, 32'sd-0.009646151171372526, 32'sd0.028360020330576836, 32'sd-0.02822885640840082, 32'sd-0.002917750421068995, 32'sd-0.03909133883480648, 32'sd0.05259681893756604, 32'sd0.0141397983416312, 32'sd-0.006994791442477023, 32'sd0.048761956931148535, 32'sd-0.0008040431360415851, 32'sd-0.05615838963226585, 32'sd0.021965664591407807, 32'sd-0.08393341666444312, 32'sd-0.1024214544089101, 32'sd-0.20767892185035683, 32'sd-0.2448620515500913, 32'sd-0.19819391578035284, 32'sd-0.1533105186214421, 32'sd0.027519626406584074, 32'sd-0.015599790020559431, 32'sd-0.1046272861396986, 32'sd-0.03541928726325722, 32'sd-0.0036837180289336635, 32'sd0.20452751976430267, 32'sd0.18111655943303576, 32'sd0.004640053030877061, 32'sd0.11421049086269994, 32'sd0.005514901849816547, 32'sd-0.10130216673049561, 32'sd0.0018580155542138885, 32'sd-0.02371837720110829, 32'sd0.047583309792445495, 32'sd-0.13256170806605086, 32'sd0.007041567610723021, 32'sd0.0189067285596702, 32'sd0.005539876977700575, 32'sd0.07655227270554589, 32'sd-0.02073323405832607, 32'sd-0.034982473742329524, 32'sd-0.10329191166161047, 32'sd0.03539587329053228, 32'sd-0.05366292540718088, 32'sd0.017943188271914153, 32'sd0.0029990019114015335, 32'sd0.04375094512216948, 32'sd-0.04001338584376782, 32'sd0.049656631306077906, 32'sd-0.02441139005402656, 32'sd0.006120599094559104, 32'sd0.02965421389809966, 32'sd0.046600733278398934, 32'sd0.06592283274794501, 32'sd0.10140613074561657, 32'sd0.09072378086834841, 32'sd0.034396008510936785, 32'sd0.02656845734615503, 32'sd-0.03676339954577073, 32'sd-0.005621084476045043, 32'sd-0.07553347134317674, 32'sd-0.0783112344881606, 32'sd-0.03456177848984917, 32'sd0.008007419528823048, 32'sd-0.015290374261407778, 32'sd0.0682624817238048, 32'sd0.053925306242006185, 32'sd-0.03869243723416764, 32'sd-0.01661409243379029, 32'sd0.012200023649735327, 32'sd0.08306115363232286, 32'sd0.05571323775302557, 32'sd0.15158943802721211, 32'sd0.05086106643192613, 32'sd0.019226026173920645, 32'sd0.11227158309579896, 32'sd0.09043121628311704, 32'sd0.003935289870970561, 32'sd-0.037319039993122645, 32'sd-0.016368256433655297, 32'sd0.09145062209433615, 32'sd0.1584941969385804, 32'sd0.20354423293343465, 32'sd0.1761942157505176, 32'sd0.13077298712020632, 32'sd-0.13132692339332622, 32'sd-0.09194301891874422, 32'sd-0.019743423420048173, 32'sd0.05235790795329144, 32'sd-0.0696578122718478, 32'sd-0.030336843301147467, 32'sd-0.04611865626634476, 32'sd0.015291388494258604, 32'sd0.07305208648463671, 32'sd0.04867970226310544, 32'sd0.05124782733544139, 32'sd-0.02917734109404703, 32'sd0.0858820029798836, 32'sd0.017352935132532936, 32'sd0.09364773415381947, 32'sd0.09548443493241071, 32'sd-0.09894620641123578, 32'sd-0.02702081806855219, 32'sd0.04758433361694471, 32'sd0.017738696014818832, 32'sd-0.1015150370334301, 32'sd-0.09860444478673525, 32'sd-0.08115858955596891, 32'sd0.010661727682877436, 32'sd0.16879129177725152, 32'sd0.04513855170377417, 32'sd0.044332246134816865, 32'sd0.09450712609120092, 32'sd-0.0905381979394183, 32'sd-0.11372328283169626, 32'sd-0.13306819578196827, 32'sd-0.06015924818183304, 32'sd-0.035118302824383066, 32'sd-0.047719490802638306, 32'sd0.011447794005947087, 32'sd-0.03373720361088225, 32'sd0.05869904072737951, 32'sd0.06864060072394759, 32'sd0.01576656808275729, 32'sd-0.06003257730617997, 32'sd0.022916590271431912, 32'sd0.05439396311973364, 32'sd0.055060882162247186, 32'sd-0.04499459744527842, 32'sd-0.04980660734406704, 32'sd-0.2568988514185878, 32'sd-0.040353740234033326, 32'sd-0.05963577590966484, 32'sd-0.021643296036547525, 32'sd-0.16586914704770672, 32'sd-0.0795708747712825, 32'sd0.0024593229966385585, 32'sd0.19273441006572845, 32'sd0.0631515191953964, 32'sd-0.03824680337467241, 32'sd0.0861518044454647, 32'sd-0.08870429955691594, 32'sd0.023650174110619464, 32'sd-0.01035483530749568, 32'sd-0.07673463079372167, 32'sd-0.04277176028214369, 32'sd0.03758993780844382, 32'sd0.06079349864158174, 32'sd-0.03957017775605904, 32'sd-0.02271936795330765, 32'sd-2.0914958280766827e-121, 32'sd0.1081466791029662, 32'sd-0.003548550407198465, 32'sd-0.010689303030311481, 32'sd-0.02726377388224763, 32'sd0.008427069277387508, 32'sd-0.134527742730021, 32'sd-0.033495922167189975, 32'sd-0.16991754824830474, 32'sd-0.14872878197767261, 32'sd-0.03511969040408723, 32'sd0.06798150841371017, 32'sd-0.06368547351109125, 32'sd-0.021397754262966154, 32'sd0.12972577119249126, 32'sd0.1633428386246603, 32'sd0.028039684325682535, 32'sd0.0171291088777848, 32'sd-0.02125614564092623, 32'sd0.02687123530345985, 32'sd-0.07638126610977962, 32'sd-0.006160040860794544, 32'sd-0.04280773067746109, 32'sd-0.028006533847309455, 32'sd0.05522026618348411, 32'sd0.0790440661591222, 32'sd0.14006590823145404, 32'sd0.046306136275341435, 32'sd-0.035779427918993474, 32'sd-0.04865682645311548, 32'sd0.052851530920808396, 32'sd0.06167870381928641, 32'sd-0.09663717184725495, 32'sd-0.05834469327293161, 32'sd-0.07296398900713684, 32'sd-0.06193108672162514, 32'sd-0.0719106475409907, 32'sd-0.007451919411891008, 32'sd-0.05929896068633255, 32'sd0.1035613955959336, 32'sd-0.026694824854493912, 32'sd-0.03900932683039579, 32'sd0.05397658419838662, 32'sd0.007106370363148047, 32'sd0.1056563338150273, 32'sd0.08793684271795332, 32'sd0.07888852611459278, 32'sd0.007373905871408724, 32'sd-0.12325872274871347, 32'sd-0.11394779513208837, 32'sd-0.046933140496457075, 32'sd0.09053403681413728, 32'sd0.10149187573321823, 32'sd0.044258326724289525, 32'sd0.04800981348296075, 32'sd0.06505178235461839, 32'sd0.09719017205817776, 32'sd0.06032066551216724, 32'sd0.028569375515231844, 32'sd0.09188433520535241, 32'sd0.03543798502660971, 32'sd-0.07163731880598997, 32'sd0.026918207142610215, 32'sd0.12668059958136108, 32'sd0.03838637477270072, 32'sd0.0827049197564788, 32'sd0.068702334774877, 32'sd0.16090509103488765, 32'sd0.10562227337203499, 32'sd-0.016084546780225084, 32'sd-0.006034415751615454, 32'sd0.03309591965696253, 32'sd0.09180751686684002, 32'sd0.054660789810638176, 32'sd-0.07829043369416139, 32'sd0.05294565989434902, 32'sd-0.01256043848240676, 32'sd-0.00806652563011681, 32'sd-0.02884390429775145, 32'sd-0.009752196290097997, 32'sd0.05426309583823925, 32'sd0.09458812790054837, 32'sd0.11989307455216132, 32'sd0.0672757334729064, 32'sd-2.7799485829261563e-124, 32'sd-0.05154651345835339, 32'sd0.012208373662649617, 32'sd-0.007418259077473475, 32'sd-0.02313771147983223, 32'sd0.04179163590586129, 32'sd-0.01308540310372919, 32'sd0.0166298478021905, 32'sd0.04793952484919267, 32'sd-0.0007738785606677787, 32'sd0.14169431093673712, 32'sd0.04793711776261774, 32'sd0.18202583927434254, 32'sd-0.04150848980950923, 32'sd-0.007026092811223752, 32'sd-0.07070065864611401, 32'sd0.13269424345966666, 32'sd0.04223602015798581, 32'sd-0.019113564555704995, 32'sd-0.006673351173224636, 32'sd-0.0030734100645359247, 32'sd0.12130354189269482, 32'sd-0.061306767129279384, 32'sd-0.023447726180943224, 32'sd-0.010814113269289183, 32'sd0.06952244139829315, 32'sd0.15120569275804985, 32'sd0.06135429287032488, 32'sd0.024477882421051065, 32'sd0.07998193187059072, 32'sd0.0454252804988085, 32'sd0.0936454284464823, 32'sd0.04883994060570826, 32'sd-0.061181585013457516, 32'sd0.044077848418256856, 32'sd0.14273139831071865, 32'sd0.04910482166760544, 32'sd-0.0030153284660502746, 32'sd0.13154385647261652, 32'sd0.13677894409498745, 32'sd0.01597476923617092, 32'sd-0.017573084827490124, 32'sd-0.02336307436189686, 32'sd-0.12327863186586403, 32'sd0.054549073424710284, 32'sd0.001510503408704984, 32'sd0.021553119777965906, 32'sd0.03345309147279853, 32'sd-0.03367393710232236, 32'sd0.12792224821661466, 32'sd-0.061098267930731205, 32'sd0.046306495291869365, 32'sd0.053055440133403915, 32'sd0.03936616965384884, 32'sd0.04340851508759348, 32'sd0.0355511075506708, 32'sd0.11558582988636085, 32'sd-0.02516038103835359, 32'sd0.04158736073895871, 32'sd0.04115919882984011, 32'sd-0.06380930728701224, 32'sd0.08991292522908563, 32'sd-0.02829985302130968, 32'sd0.09297028382860811, 32'sd0.1245332518326794, 32'sd-0.026351904515553706, 32'sd0.01998779483553577, 32'sd-0.06336442438051891, 32'sd0.0008681213054126358, 32'sd-0.062355535266812326, 32'sd-0.05430456600376289, 32'sd0.06607061360935611, 32'sd0.07913651516967084, 32'sd-0.05118126526382679, 32'sd-0.01187774222267526, 32'sd-0.05050716901865948, 32'sd-0.02690651549195678, 32'sd0.0010251914894104813, 32'sd0.04265971710108273, 32'sd0.10258456556230883, 32'sd0.015001877049064466, 32'sd-0.008193488598541266, 32'sd-0.06604320373231659, 32'sd0.09598789836221765, 32'sd-6.464573829707675e-121, 32'sd0.0474135780397248, 32'sd-0.058080940251532855, 32'sd0.037250697203864466, 32'sd-0.01781829730995304, 32'sd0.1043605610491846, 32'sd-0.0006762068141700181, 32'sd0.029776407744499835, 32'sd-0.08881070657479888, 32'sd0.08497389689311236, 32'sd-0.10257644495962266, 32'sd-0.015243236963703282, 32'sd-0.08758522073177587, 32'sd0.09971745773438233, 32'sd-0.04969146980929494, 32'sd-0.0433883506616715, 32'sd0.05801389695076635, 32'sd0.01604326506330146, 32'sd-0.09069950603147849, 32'sd0.009713839382529949, 32'sd-0.0651100961036758, 32'sd-0.029609633918277374, 32'sd-0.004050232077999178, 32'sd0.009550001992088008, 32'sd0.056831644449441006, 32'sd0.0949937374006772, 32'sd-0.06876187573881425, 32'sd-6.450163763464977e-122, 32'sd1.8173885766737615e-123, 32'sd7.2590113921145365e-115, 32'sd0.13330084811055373, 32'sd-0.023265306154445952, 32'sd0.11737843628682176, 32'sd0.015287494357232673, 32'sd-0.0017426890018229497, 32'sd-0.04418240135797799, 32'sd0.09094333221002769, 32'sd-0.04484108318316263, 32'sd-0.11560584203218154, 32'sd-0.10690345394241657, 32'sd-0.04233530644664049, 32'sd-0.0037652511410951927, 32'sd0.02611414469854227, 32'sd0.06769991614637606, 32'sd-0.08387637045741764, 32'sd-0.025734602664705904, 32'sd-0.12316934250120742, 32'sd-0.23351767838856866, 32'sd-0.09885153597962756, 32'sd-0.014656082625711424, 32'sd-0.12398608720266627, 32'sd-0.006731673353307548, 32'sd0.07821338719857918, 32'sd-0.02025291726122407, 32'sd0.009716160232467458, 32'sd-3.4688655016419963e-116, 32'sd-7.860085335829358e-121, 32'sd-2.341252717828242e-124, 32'sd0.05577958824786365, 32'sd0.018969630741499956, 32'sd0.13886925423338312, 32'sd0.06544921721646832, 32'sd0.03601952315667887, 32'sd0.14949803396344422, 32'sd0.1015415623463565, 32'sd-0.01761876223761603, 32'sd-0.12016695913533608, 32'sd0.01741537523462712, 32'sd-0.014459765826228916, 32'sd0.03389176538552483, 32'sd0.041305020998054914, 32'sd-0.14554867251855041, 32'sd0.009147682567513452, 32'sd0.07078037205479697, 32'sd-0.07041310291774512, 32'sd-0.09849416151509977, 32'sd-0.06025954740872646, 32'sd-0.006166249148557464, 32'sd0.013836914529576924, 32'sd0.045853006836012615, 32'sd-0.01511011718126204, 32'sd-0.020120840753202307, 32'sd-0.0036450624010978348, 32'sd6.881660852024408e-126, 32'sd1.6831763107363274e-123, 32'sd3.2957548168048476e-125, 32'sd-3.6677324222084895e-118, 32'sd0.0927787920390924, 32'sd-0.000266200706327812, 32'sd-0.027395728551936498, 32'sd0.0034584110627078443, 32'sd0.1066830237178431, 32'sd0.10935022948536126, 32'sd-0.008940651863523582, 32'sd0.025817715393710892, 32'sd0.20098591001442778, 32'sd0.04906740498173139, 32'sd-0.0401249645446968, 32'sd0.1648463478756988, 32'sd0.01355891027743626, 32'sd0.0659399637207607, 32'sd0.15189045328312345, 32'sd0.047858837443759704, 32'sd-0.04595440261533774, 32'sd0.015349198424241003, 32'sd-0.020674779588759722, 32'sd-0.0933389313213451, 32'sd-0.043518572139627364, 32'sd0.048844616607391096, 32'sd0.07773150281407126, 32'sd6.882299162108198e-124, 32'sd5.093366118727582e-126, 32'sd-8.854201962383452e-120, 32'sd7.727541910548805e-117, 32'sd-1.3122366843506632e-119, 32'sd-9.309903370415724e-119, 32'sd0.08106143126041926, 32'sd0.04711013983163249, 32'sd0.09529766164863834, 32'sd0.1162603612933563, 32'sd0.059662267516054676, 32'sd0.058482189639867836, 32'sd0.14046107329125235, 32'sd0.05769246496375255, 32'sd0.08600341775129046, 32'sd0.1252217672876216, 32'sd0.13550111400596618, 32'sd0.03801852972218326, 32'sd0.0771335012965629, 32'sd0.13861214168597863, 32'sd0.06252581800507688, 32'sd0.014733854798931545, 32'sd0.043923550225452905, 32'sd0.007587236296814792, 32'sd-0.009289809025813544, 32'sd0.05272718406434466, 32'sd-4.904619166958554e-122, 32'sd1.5846511246815342e-122, 32'sd-1.0345165126300541e-120, 32'sd-1.6582499297582674e-114},
        '{32'sd6.480278010960618e-123, 32'sd1.5776519272696328e-124, 32'sd-1.9150652194991042e-129, 32'sd3.0920312703830346e-114, 32'sd1.3005806859338882e-118, 32'sd-1.2982282571690763e-123, 32'sd-2.13885864008648e-116, 32'sd-3.819949740469736e-118, 32'sd-1.4289490649939346e-118, 32'sd8.199281315769111e-120, 32'sd9.898838952087146e-124, 32'sd7.75275292841249e-115, 32'sd0.05607763679002849, 32'sd0.07929464067518088, 32'sd0.06565320902182166, 32'sd0.0011634615243523454, 32'sd1.0328026459283221e-120, 32'sd-2.616222739182131e-124, 32'sd9.222608597710647e-119, 32'sd-1.3226165533504095e-118, 32'sd-9.145864715171459e-125, 32'sd-2.81836153923611e-120, 32'sd-4.094371325294121e-124, 32'sd7.240309290378014e-115, 32'sd7.101138343291426e-122, 32'sd-4.1545009498844765e-117, 32'sd-1.2306453657410407e-123, 32'sd2.3174325857281585e-121, 32'sd9.126537977965947e-122, 32'sd7.251946703652433e-115, 32'sd-1.6290597262691164e-115, 32'sd-8.970692589315852e-127, 32'sd-0.09768292955105219, 32'sd0.044221654522539115, 32'sd0.0801203305773085, 32'sd0.04576815976709667, 32'sd-0.0055188601201979935, 32'sd-0.030983196608189108, 32'sd0.09830315751150748, 32'sd0.07577523416215447, 32'sd0.11915890526727382, 32'sd0.06905248144821631, 32'sd0.004419388300400283, 32'sd-0.03435789588878651, 32'sd0.020799711043020676, 32'sd0.06730061701069176, 32'sd0.05731727636653924, 32'sd-0.012933114759356983, 32'sd0.09053234809217664, 32'sd-0.0016214431787829288, 32'sd0.07871565523919045, 32'sd0.032164501843339896, 32'sd7.440224253596854e-117, 32'sd-4.663584196139049e-126, 32'sd6.218687728234296e-125, 32'sd-8.044593225494512e-122, 32'sd1.2792163255542683e-122, 32'sd-1.0473082529735779e-121, 32'sd0.03469487464813241, 32'sd0.029029244618639642, 32'sd0.008603375239057553, 32'sd0.00582999284380153, 32'sd0.03403050367767374, 32'sd0.05801766278548225, 32'sd0.09109051404306669, 32'sd0.09680130956036166, 32'sd0.16313854489430468, 32'sd0.0891561960344003, 32'sd-0.03389367309941309, 32'sd-0.007169265131701112, 32'sd0.03149706004723385, 32'sd-0.0014294146056837444, 32'sd0.00930166770073328, 32'sd-0.003918056971596325, 32'sd0.0580835156055252, 32'sd0.044236715763867465, 32'sd-0.04219196723008368, 32'sd0.08969593000191768, 32'sd0.04410820497610219, 32'sd-0.08139736672970024, 32'sd0.03628343890032566, 32'sd0.024011899006301185, 32'sd-6.93529064207222e-123, 32'sd2.252650655133562e-126, 32'sd1.3854442731145362e-118, 32'sd1.3190110062296703e-123, 32'sd0.07948163520710784, 32'sd0.05168596332285389, 32'sd0.040905053604234, 32'sd-0.005269352163696072, 32'sd0.12901167214717352, 32'sd0.0334980210304087, 32'sd-0.03694649780465859, 32'sd0.06343446581650114, 32'sd0.062242134927403193, 32'sd-0.030615036716751514, 32'sd-0.16888113102011254, 32'sd-0.018389397145270305, 32'sd-0.029065300295076056, 32'sd0.02845354875425864, 32'sd0.07766012785772758, 32'sd0.08330399016431768, 32'sd-0.08853884944513098, 32'sd-0.03818746566549584, 32'sd-0.1628106942417013, 32'sd-0.045169288616542326, 32'sd0.0523515971079478, 32'sd0.036338702398973646, 32'sd-0.025311008227986345, 32'sd-0.03749599489841217, 32'sd-0.007024170522961522, 32'sd2.277183101656646e-121, 32'sd1.7882350375537608e-126, 32'sd-0.007363632140698072, 32'sd0.013663558433593815, 32'sd-0.028271788293796053, 32'sd-0.03328701934945818, 32'sd-0.026256682655125218, 32'sd0.03211118845845757, 32'sd-0.12187070792221767, 32'sd-0.0021381628671615607, 32'sd0.001185431595942638, 32'sd-0.0014005641948364044, 32'sd-0.03529664763349785, 32'sd-0.12814358570564438, 32'sd-0.08805482011886095, 32'sd-0.07858880128279717, 32'sd-0.0906159841610138, 32'sd0.11488020143388597, 32'sd0.04315879631973433, 32'sd-0.09347652324522887, 32'sd-0.025317790153135296, 32'sd-0.08785054850217554, 32'sd-0.11561229919292569, 32'sd-0.1735157520616246, 32'sd-0.11649615968025416, 32'sd0.06376480205677688, 32'sd0.03330483795429553, 32'sd0.0062367597986250295, 32'sd-0.01722417628289756, 32'sd2.4419910892172875e-122, 32'sd0.07239876678945861, 32'sd0.06748152166878137, 32'sd0.020752789714148005, 32'sd0.05596670083663341, 32'sd-0.11209329489584365, 32'sd0.009037911967916503, 32'sd0.068668946683482, 32'sd0.05762361037632384, 32'sd0.05656198817277984, 32'sd0.050341383641043784, 32'sd0.045612666817712, 32'sd0.04819484513181987, 32'sd-0.07357471100489067, 32'sd-0.12722343926116034, 32'sd-0.11676553022705576, 32'sd0.05234496111828511, 32'sd-0.0018307269639565497, 32'sd-0.11472847538298442, 32'sd-0.0465962512789293, 32'sd-0.0349749777082646, 32'sd-0.025252091509946693, 32'sd0.09480407337493942, 32'sd-0.01962039237780348, 32'sd0.052961884138339174, 32'sd-0.03288150911992996, 32'sd-0.08922234897087568, 32'sd0.04818209364618019, 32'sd2.1117010416729806e-124, 32'sd0.017797578056544732, 32'sd-0.05385641600420499, 32'sd0.031743647718341456, 32'sd-0.032147451482975146, 32'sd-0.09893351795124303, 32'sd0.05581674849505855, 32'sd0.08597691395172247, 32'sd0.1630708599930282, 32'sd0.09269526244847345, 32'sd-0.07309247549534038, 32'sd-0.06291617378143027, 32'sd-0.03965154325004671, 32'sd-0.08959799389964886, 32'sd0.03342405348703543, 32'sd-0.040871264334090815, 32'sd-0.08234818163803793, 32'sd-0.05103190205773396, 32'sd-0.03663561201735367, 32'sd-0.07268038516972443, 32'sd-0.04157916876154467, 32'sd0.049471800259058764, 32'sd0.03662622615875984, 32'sd-0.04664740882830409, 32'sd-0.1717059806365714, 32'sd0.01090566247490743, 32'sd0.0011478836318600364, 32'sd0.05737985258454392, 32'sd0.033946167902823836, 32'sd0.11614147940215537, 32'sd-0.06502718370395671, 32'sd-0.01788559454630603, 32'sd0.0551033211102261, 32'sd-0.019003099135629316, 32'sd-0.017633302626529578, 32'sd0.10155780958658733, 32'sd0.17248558174872203, 32'sd0.09875434482854299, 32'sd-0.07796226709618347, 32'sd-0.06170448610860895, 32'sd-0.0864687399126435, 32'sd-0.02447273324039994, 32'sd0.0015765084668249447, 32'sd0.014229964974806483, 32'sd-0.12353160951702725, 32'sd0.03835336282439082, 32'sd-0.0801915124645699, 32'sd0.08544133816568562, 32'sd0.01760974935047685, 32'sd-0.03444258837424348, 32'sd-0.15106254823962173, 32'sd-0.15143382932654603, 32'sd-0.08287691668472837, 32'sd0.016138706912466442, 32'sd0.02437919814268238, 32'sd-0.0032733526469416307, 32'sd0.08579528563014768, 32'sd0.04967840232346019, 32'sd-0.06560611282998033, 32'sd-0.026719777098174767, 32'sd0.11917024960846095, 32'sd-0.08154589421858296, 32'sd0.09979876801533565, 32'sd0.191244634740913, 32'sd0.0075103214827251874, 32'sd0.13218768508310832, 32'sd-0.04864205424057531, 32'sd-0.14061092046547605, 32'sd-0.0992807800350416, 32'sd0.08843298887401489, 32'sd0.001019560724640867, 32'sd-0.045696330375480515, 32'sd0.05915721833041058, 32'sd-0.04733056703083092, 32'sd-0.08185233514635969, 32'sd0.07648138308617186, 32'sd0.07013221663272985, 32'sd0.09365542603414696, 32'sd-0.09871731951863108, 32'sd-0.08354795731830131, 32'sd0.058442208673447564, 32'sd-0.025085605589361504, 32'sd0.006456670094318801, 32'sd-0.016593029202515524, 32'sd0.08324972747298466, 32'sd-0.03690453934003031, 32'sd-0.10569320533847916, 32'sd0.021299611991359206, 32'sd0.1538431337355152, 32'sd0.02598563881569909, 32'sd-0.04992624040130247, 32'sd0.040756058585246835, 32'sd0.055791617161391596, 32'sd0.020814478281468436, 32'sd0.059158565478704406, 32'sd-0.10206648921870955, 32'sd0.02780681531354479, 32'sd-0.021696513342584253, 32'sd-0.05253926318646944, 32'sd-0.0014144867137852678, 32'sd0.12491475108361144, 32'sd0.12093137471173954, 32'sd-0.07128366970909042, 32'sd-0.007828155297182513, 32'sd0.1033133916949772, 32'sd-0.04916599295293315, 32'sd-0.024850105313481568, 32'sd-0.08517991311930934, 32'sd-0.06097624707730467, 32'sd-0.06028040830067601, 32'sd-0.04418689516163305, 32'sd0.00929694888134564, 32'sd0.04400727937415579, 32'sd0.0728147874249501, 32'sd0.03166555130025834, 32'sd-0.013666322248057939, 32'sd-0.0320270039064706, 32'sd0.015824211039991983, 32'sd0.04293516890407716, 32'sd0.043697470754783085, 32'sd0.0999943088246204, 32'sd0.08195605286396963, 32'sd-0.008245228656585831, 32'sd-0.0017809062545785432, 32'sd-0.0671757665581098, 32'sd-0.0381584493626258, 32'sd-0.09480494696382427, 32'sd0.01738599613066494, 32'sd0.04279311536645581, 32'sd-0.0059556750725282106, 32'sd-0.0852801854440558, 32'sd-0.0982752007241572, 32'sd0.013053782359967814, 32'sd-0.05977842997969982, 32'sd-0.017845384478381035, 32'sd-0.16363184183033647, 32'sd0.009269544456917267, 32'sd-0.07703493365205641, 32'sd0.006246384106536444, 32'sd-0.09129590006647584, 32'sd-0.025969753579381073, 32'sd-0.07699699598599487, 32'sd0.006541177966968409, 32'sd0.05122942569027991, 32'sd0.06545380045192169, 32'sd0.08639710034139514, 32'sd0.0005307559230625122, 32'sd0.031466969457243796, 32'sd0.055804492649064126, 32'sd0.07194301180632796, 32'sd0.019509774525211184, 32'sd-0.0720204067027418, 32'sd-0.08101144865783162, 32'sd-0.05527807523408051, 32'sd0.018425763390604033, 32'sd0.09302168095683384, 32'sd0.13245019936855532, 32'sd0.020650707905316187, 32'sd-0.04472850432624708, 32'sd0.0114894086286432, 32'sd0.03757268132635902, 32'sd-0.04236190779768258, 32'sd-0.001111561329735646, 32'sd-0.16155974719529917, 32'sd-0.18146453101032464, 32'sd0.0762872380723122, 32'sd0.012969413249206384, 32'sd-0.09912895836017915, 32'sd0.09002139384209688, 32'sd-0.05401983966308833, 32'sd0.06616302772938104, 32'sd-0.03999918010753944, 32'sd0.10919726023596125, 32'sd-0.0020498379305522196, 32'sd-0.15965563391751833, 32'sd0.022935301085815978, 32'sd0.07619840242178287, 32'sd0.026801503343339694, 32'sd-0.08819535135806009, 32'sd-0.032701906758670164, 32'sd-0.18242470156245003, 32'sd0.048618502972705556, 32'sd0.0249708268164429, 32'sd0.20730447810805078, 32'sd0.018975007327235466, 32'sd-0.040111388281800164, 32'sd0.006834887928059699, 32'sd-0.046517854747186255, 32'sd0.01580147711113508, 32'sd0.04441207527371376, 32'sd-0.014112703403701651, 32'sd-0.1838149342151077, 32'sd-0.0937868588122987, 32'sd0.05977254600614324, 32'sd-0.03590248811080236, 32'sd-0.020795716142796156, 32'sd0.03969902643603709, 32'sd-0.07077533997807972, 32'sd0.04971466041649405, 32'sd0.10900671988468125, 32'sd0.023681765943391442, 32'sd0.07823442753148895, 32'sd-0.0289319003670577, 32'sd-0.04822508566803308, 32'sd0.019616941298317654, 32'sd-0.07715160434000146, 32'sd-0.07099155956139594, 32'sd-0.017764110510802365, 32'sd-0.009084676029745197, 32'sd0.1349213573399957, 32'sd0.024081639618007317, 32'sd0.15857165481453778, 32'sd-0.08045146405898276, 32'sd-0.07111320627837127, 32'sd0.07043670989763307, 32'sd0.009341887035312073, 32'sd0.018797032838168526, 32'sd0.03486780352685896, 32'sd0.04022347406439636, 32'sd-0.01807972176715786, 32'sd-0.09963758189408865, 32'sd0.05854101746777814, 32'sd0.00890317059616005, 32'sd0.030194370772080294, 32'sd-0.011081570498401642, 32'sd0.0046280211335856195, 32'sd-0.05060261336130791, 32'sd0.0504505284952816, 32'sd0.12369835158279772, 32'sd0.026180876826401814, 32'sd0.01424244238544728, 32'sd-0.13879359657159746, 32'sd-0.03958218826605395, 32'sd-0.05361281602488856, 32'sd-0.15428494335653262, 32'sd-0.044381524543058895, 32'sd0.009376241074931168, 32'sd0.17769694760625881, 32'sd0.145759338797103, 32'sd-0.06983073121777303, 32'sd-0.1236909019883956, 32'sd0.05529912109237637, 32'sd0.12870993440691889, 32'sd0.16040609158965466, 32'sd0.038546662209988015, 32'sd-0.08204869850948336, 32'sd-0.08380720574360401, 32'sd0.11322834428426587, 32'sd-0.03832912696498331, 32'sd0.010779761971258172, 32'sd0.05491517258231123, 32'sd0.0469574412709802, 32'sd-0.002506216160871287, 32'sd0.030273235583765344, 32'sd-0.03674634860951219, 32'sd0.009166180011222257, 32'sd-0.038269225070590975, 32'sd-0.12391176395055926, 32'sd-0.02385293062839955, 32'sd-0.07349026833049474, 32'sd-0.08154987246571667, 32'sd-0.1158762319482362, 32'sd-0.10721757843428427, 32'sd0.08623442551028143, 32'sd0.07302621923457252, 32'sd0.19788729377015005, 32'sd0.1288940345539188, 32'sd-0.016304177998655574, 32'sd-0.09087238468907716, 32'sd-0.12455940523948904, 32'sd0.027762278125513424, 32'sd0.05017360901143535, 32'sd0.07745661313208817, 32'sd0.012006356408182591, 32'sd-0.022908093793103327, 32'sd0.12659069098064607, 32'sd0.07904340928926201, 32'sd-0.04296443362441256, 32'sd0.03843126748462523, 32'sd0.019660760541133648, 32'sd0.06283213027868344, 32'sd0.07768958900699681, 32'sd-0.04559486730900061, 32'sd0.0805373229415446, 32'sd-0.0911288983638181, 32'sd0.041386458578140724, 32'sd0.012553164268439053, 32'sd-0.06796946894471906, 32'sd-0.14110769896212294, 32'sd-0.2450252801262606, 32'sd-0.10510592212944259, 32'sd0.14047342167399587, 32'sd0.1217096313036365, 32'sd0.10494098658875729, 32'sd0.13552491597118174, 32'sd0.033364165738057866, 32'sd-0.0034230495178841944, 32'sd-0.05660070687348498, 32'sd-0.09333491550005729, 32'sd0.057239884902360226, 32'sd0.07095337642143669, 32'sd-0.0669717544919832, 32'sd0.11711653711677161, 32'sd0.1790908756746328, 32'sd0.041301446957174005, 32'sd0.011351812984197787, 32'sd-0.03831719163332713, 32'sd-0.021655241285962353, 32'sd-1.099657523609797e-127, 32'sd-0.06650962250635326, 32'sd0.03903290721955047, 32'sd0.0570436972400488, 32'sd0.022655830620748142, 32'sd-0.06837171745990944, 32'sd-0.11730352176531691, 32'sd-0.08009535561240291, 32'sd-0.3052722445397893, 32'sd-0.18922401915154588, 32'sd0.11376540334686443, 32'sd0.13442263806903412, 32'sd0.23925061786055865, 32'sd0.066527578718622, 32'sd-0.022313211236027888, 32'sd0.04134972537579498, 32'sd0.026493939551246258, 32'sd0.11763956473785539, 32'sd0.05866140544625845, 32'sd0.11322008045487536, 32'sd0.041723024365392075, 32'sd0.0031468879645459628, 32'sd-0.044241271323654914, 32'sd0.04029897254388587, 32'sd-0.04154342396459207, 32'sd-0.027753506871194288, 32'sd-0.05515752567846489, 32'sd-0.018575019192492073, 32'sd0.025464359567447376, 32'sd0.014680371067032516, 32'sd-0.010197415203605918, 32'sd-0.016814716953186405, 32'sd-0.06917974642335888, 32'sd-0.014453596032769815, 32'sd-0.1448766725435149, 32'sd-0.16846662451005207, 32'sd-0.20451959083576704, 32'sd-0.01874639520834133, 32'sd0.1607197601090079, 32'sd0.18630821712299092, 32'sd0.24838907849355654, 32'sd0.21698925975716518, 32'sd-0.03341070746482677, 32'sd0.02757364596983926, 32'sd-0.041032847131616215, 32'sd-0.005797945264427469, 32'sd0.0938817359404101, 32'sd-0.0029315254417901205, 32'sd-0.02947341717409361, 32'sd0.006000603293763341, 32'sd-0.03309644893341903, 32'sd-0.19936367693542242, 32'sd-0.009585826710411789, 32'sd-0.03384673886754457, 32'sd-0.04200741656241181, 32'sd-0.023415316523553182, 32'sd0.058884450286709696, 32'sd0.01374548861655017, 32'sd-0.10128985219993983, 32'sd-0.05005365473306061, 32'sd0.012649239711454483, 32'sd-0.033617645656522206, 32'sd-0.07913311862143614, 32'sd-0.16711480708107546, 32'sd-0.2091374565539352, 32'sd-0.06964562865415794, 32'sd0.11053781892997515, 32'sd0.057287744099388985, 32'sd0.08761216592925987, 32'sd0.16610135623410274, 32'sd0.004808569607432593, 32'sd-0.05307514183371764, 32'sd0.09157601077732258, 32'sd0.03320782153010548, 32'sd-0.061523352103269854, 32'sd0.03499276079311673, 32'sd-0.022052894025152064, 32'sd-0.0268368818139888, 32'sd-0.12078416650953677, 32'sd-0.05416653580617696, 32'sd-0.08870532393783687, 32'sd-0.03375233744785365, 32'sd-0.012879755277469205, 32'sd0.00325115003825893, 32'sd-1.4234178570985371e-127, 32'sd0.029882418161636753, 32'sd-0.07195367089720599, 32'sd-0.022645384432704634, 32'sd0.0025358879813701727, 32'sd-0.13596202038910318, 32'sd-0.08128630839958075, 32'sd-0.17993400545945448, 32'sd-0.17027544360188457, 32'sd-0.1600597871420189, 32'sd-0.021240739730264427, 32'sd0.14654408090535403, 32'sd0.06332663072143575, 32'sd0.10494060771212244, 32'sd0.04454122811197373, 32'sd0.08325423091935029, 32'sd0.0010954972789713198, 32'sd0.06919284229299744, 32'sd0.02173712034502207, 32'sd-0.06290121550673848, 32'sd0.05229997387058548, 32'sd-0.004568006122004472, 32'sd-0.15800401780171774, 32'sd-0.15396736011681705, 32'sd0.04651966096195986, 32'sd0.041394689812874925, 32'sd0.0230009628983981, 32'sd0.0025513294690524897, 32'sd0.0022233027088917772, 32'sd-0.0673659882003935, 32'sd-0.00999803537357812, 32'sd0.011093992130356287, 32'sd-0.059349182263255376, 32'sd-0.08715957783854815, 32'sd-0.013133825044464954, 32'sd-0.0583331162049323, 32'sd-0.14958285350679074, 32'sd-0.17596745698263433, 32'sd-0.07104011622586703, 32'sd-0.06644275722812572, 32'sd0.06406004635290123, 32'sd0.19447000181993557, 32'sd0.173329031080618, 32'sd0.09639029680822142, 32'sd0.13689597300727943, 32'sd-0.026218810669054828, 32'sd-0.0639870723862135, 32'sd0.026274523628693185, 32'sd-0.1121589991865418, 32'sd-0.11001383562249616, 32'sd-0.040206293645915596, 32'sd0.08561676557695788, 32'sd-0.07841270124277343, 32'sd0.008163126299448554, 32'sd-0.046277528098944816, 32'sd0.02126964131411776, 32'sd-0.008877753890227713, 32'sd-0.044204253178044765, 32'sd0.015706182524256124, 32'sd-0.0349815561143032, 32'sd-0.007259006216503254, 32'sd0.035193729933483776, 32'sd-0.02656248525399463, 32'sd-0.11414912719451054, 32'sd-0.11333435458299132, 32'sd-0.18220720271546925, 32'sd-0.1606729552949202, 32'sd-0.030605363888288804, 32'sd0.1449287657899294, 32'sd0.04557455839639896, 32'sd0.07102931492877212, 32'sd0.059687981718748805, 32'sd0.08049644795951075, 32'sd0.08571672924772056, 32'sd-0.10608207629609935, 32'sd-0.03695072622934619, 32'sd-0.12242625854336237, 32'sd-0.14645390971923514, 32'sd-0.008773915682304775, 32'sd0.0332054065592351, 32'sd-0.15779444974681384, 32'sd-0.053608135515563045, 32'sd-0.10260975573923098, 32'sd0.05573844280109228, 32'sd3.1659316605117834e-122, 32'sd0.01587578443086035, 32'sd-0.021725526922014272, 32'sd-0.039940802519318024, 32'sd-0.10890065919989038, 32'sd-0.06980911438482194, 32'sd-0.0768934552206965, 32'sd-0.09712214567726409, 32'sd-0.09663905763456794, 32'sd-0.12002367007051278, 32'sd-0.12737370759387823, 32'sd-0.06384446142324923, 32'sd0.04409623576922393, 32'sd0.06530318632203219, 32'sd0.11605768961708465, 32'sd0.0826473751654443, 32'sd0.11713531918505606, 32'sd-0.0016679904951045791, 32'sd-0.09494812299654391, 32'sd-0.009728798861417105, 32'sd-0.054747552723988846, 32'sd0.03815854056777155, 32'sd-0.00878872456117725, 32'sd0.015976869686610256, 32'sd0.0002748501102366266, 32'sd0.014870860105172875, 32'sd0.029241941701650006, 32'sd3.938220757612401e-129, 32'sd-4.705914219963964e-123, 32'sd3.74687645481902e-122, 32'sd0.012098207852310583, 32'sd-0.0488194958418004, 32'sd-0.04309697228558416, 32'sd-0.016355320751420276, 32'sd-0.10268098982488938, 32'sd-0.06832684063400829, 32'sd-0.09430206065157772, 32'sd-0.07987810745390603, 32'sd-0.11023395722536579, 32'sd-0.07866949285486047, 32'sd-0.10506123103740782, 32'sd-0.036803609967516575, 32'sd0.11034935642957447, 32'sd-0.02892306812255057, 32'sd-0.025901939685985094, 32'sd-0.08482571577258384, 32'sd-0.09415362811626114, 32'sd-0.04724054026511464, 32'sd-0.004475017493082357, 32'sd-0.10755214500384434, 32'sd-0.014494026855702256, 32'sd0.03736527474744844, 32'sd-0.06716008445131007, 32'sd-0.07114459525875577, 32'sd-0.004383817636024338, 32'sd1.6574352269031014e-126, 32'sd9.042081821300258e-126, 32'sd-2.289364373769216e-119, 32'sd-0.003304139789724726, 32'sd0.013247886133772807, 32'sd-0.01880449511286397, 32'sd0.03105622461473567, 32'sd-0.10074042222550714, 32'sd0.027891278858665873, 32'sd-0.03028712909178015, 32'sd-0.07232432904802873, 32'sd-0.12103765003652503, 32'sd-0.11949666865297671, 32'sd-0.1181827073367316, 32'sd-0.1681792727897346, 32'sd-0.047279644638479064, 32'sd0.002290210528062497, 32'sd-0.11719422116673174, 32'sd-0.025639919670138924, 32'sd-0.19397004864511633, 32'sd0.011893466284854796, 32'sd0.05142810501774786, 32'sd-0.08468824563235773, 32'sd-0.1308679606935281, 32'sd-0.0008640158596411525, 32'sd0.03878910142728177, 32'sd0.035075462068033414, 32'sd0.057321135527067926, 32'sd-2.4980112539132454e-124, 32'sd2.8695232590413897e-125, 32'sd-9.421408869040804e-122, 32'sd3.148765852785346e-121, 32'sd0.06900525432479097, 32'sd-0.005594650274356237, 32'sd-0.053343469155855756, 32'sd0.04978595698352775, 32'sd0.07846661889287197, 32'sd0.06799948766437167, 32'sd-0.03415564292752838, 32'sd-0.04895576119110068, 32'sd0.009763820184686625, 32'sd-0.044611546699303145, 32'sd-0.11128011159626774, 32'sd-0.11514676151349855, 32'sd-0.08537814317247892, 32'sd-0.0061374816275061245, 32'sd0.037061218551509484, 32'sd-0.03243604136544196, 32'sd-0.10673768839890446, 32'sd0.002382181656656127, 32'sd-0.11155094004433247, 32'sd-0.09323365956400824, 32'sd-0.014031929607712755, 32'sd0.020011660008627776, 32'sd0.06065483840694139, 32'sd6.963960244099767e-126, 32'sd1.7802761998652084e-127, 32'sd2.5413309327392826e-118, 32'sd2.1511799900288445e-116, 32'sd3.0956363764523803e-116, 32'sd-5.952140352985278e-126, 32'sd0.05257913325913852, 32'sd0.015545315677114811, 32'sd0.08578294512886799, 32'sd0.10262600471369761, 32'sd0.009338636895224715, 32'sd-0.02883964986052566, 32'sd-0.013571672578931382, 32'sd0.0693762968356901, 32'sd-0.0630157592487469, 32'sd0.026223398683342822, 32'sd-0.04555788143704304, 32'sd-0.0231011400229173, 32'sd0.04161492076888192, 32'sd0.06790140714627421, 32'sd-0.0239355286781085, 32'sd0.1970015641591663, 32'sd0.12932187179846977, 32'sd-0.05813659330376422, 32'sd-0.04450174405827197, 32'sd0.07625048997812109, 32'sd6.712051827093395e-122, 32'sd1.484135368781419e-115, 32'sd-2.3295015544810965e-124, 32'sd1.0591996016425507e-121},
        '{32'sd-2.0833888229681025e-117, 32'sd4.703814493775803e-127, 32'sd-2.7053243466751386e-122, 32'sd-8.964754272153029e-116, 32'sd-1.9521479897008922e-119, 32'sd-8.697281018994053e-119, 32'sd2.3162388320819008e-124, 32'sd-6.8952474424478695e-124, 32'sd-4.675824706664407e-121, 32'sd-3.0245573005047515e-117, 32'sd-4.63448759017804e-124, 32'sd1.4263313583379392e-127, 32'sd0.09932662430778043, 32'sd0.02060761376932684, 32'sd-0.0019137211974365842, 32'sd-0.0018840269270589034, 32'sd3.184796359236657e-123, 32'sd-6.494018765093338e-126, 32'sd-1.0663177425479179e-125, 32'sd-2.5875261351585503e-122, 32'sd-1.0148905479689235e-124, 32'sd1.5551940438653719e-115, 32'sd3.202276437247793e-120, 32'sd-1.4623341718426228e-115, 32'sd3.1656452572730955e-114, 32'sd-8.6375417358767e-117, 32'sd1.3415550238127067e-122, 32'sd-3.237177993562621e-122, 32'sd-1.9277480986469746e-120, 32'sd-1.9379138584693677e-118, 32'sd6.094334229773718e-115, 32'sd-1.0443681147644408e-122, 32'sd0.05966924147882617, 32'sd0.03940066646590148, 32'sd-0.027860620466874274, 32'sd-0.0813940800864401, 32'sd-0.044911479142896595, 32'sd-0.11070096276826831, 32'sd0.04041062893801814, 32'sd-0.03941694529931141, 32'sd0.09077787744171413, 32'sd0.008648772408911713, 32'sd0.060835452763813566, 32'sd-0.03344682855375985, 32'sd0.028981627306248144, 32'sd0.008041228778502775, 32'sd-0.002353841213813222, 32'sd0.05278126982690117, 32'sd0.08999588034957966, 32'sd0.06136526181137241, 32'sd0.029998622989539262, 32'sd-0.009121785627400429, 32'sd1.1960692457254133e-122, 32'sd-8.773300540277626e-125, 32'sd-7.438431804939152e-123, 32'sd-1.3134460792503792e-115, 32'sd-8.485845306138602e-122, 32'sd2.0577653791421774e-118, 32'sd0.005353896119193479, 32'sd0.04816176022266782, 32'sd0.09674058440913663, 32'sd-0.040256874042659554, 32'sd-0.018088230443307395, 32'sd-0.11136928828546044, 32'sd0.055749254276292355, 32'sd0.04164608926992634, 32'sd0.06472849033391008, 32'sd-0.040470583949332006, 32'sd0.005495202901315366, 32'sd0.03219746772033095, 32'sd-0.07179096582092909, 32'sd0.03757744401659058, 32'sd0.006188005429463503, 32'sd0.035489935480524135, 32'sd-0.03544333567249435, 32'sd0.02405591933650528, 32'sd-0.061758041640455855, 32'sd-0.0941796545516765, 32'sd-0.05908447885180401, 32'sd0.03547229617865126, 32'sd0.06382417006537021, 32'sd0.011192995222728134, 32'sd2.729847925650699e-127, 32'sd-9.960373846911969e-118, 32'sd1.0348264902003473e-118, 32'sd-1.156769338189571e-127, 32'sd-0.04924027816051629, 32'sd0.015966515453224174, 32'sd-0.05005759214035756, 32'sd-0.09062039412128314, 32'sd0.040492154430381115, 32'sd-0.02405284437530262, 32'sd0.05420589834920314, 32'sd-0.05339952268898949, 32'sd0.005041551473990882, 32'sd0.040495231926412814, 32'sd0.07266634352162815, 32'sd0.02829521701161885, 32'sd0.08213864238468445, 32'sd0.0471113861723957, 32'sd-0.1069625289429854, 32'sd-0.015763341197820024, 32'sd-0.09239639026398877, 32'sd-0.041618982211008855, 32'sd0.001855263567353354, 32'sd0.04054227244225302, 32'sd0.09200241793587367, 32'sd0.03226861810000939, 32'sd-0.019216956268578823, 32'sd0.05231168927931542, 32'sd0.002186167615436492, 32'sd3.774753840557497e-122, 32'sd-7.337712829787349e-117, 32'sd0.018479544527190514, 32'sd0.05387051643856977, 32'sd-0.05788471723669106, 32'sd-0.023737084160608046, 32'sd0.0071617788460595685, 32'sd-0.054334464613696995, 32'sd-0.06909449697372179, 32'sd-0.059241173627285384, 32'sd-0.056138388054393897, 32'sd-0.17199767086102305, 32'sd0.00620920533495017, 32'sd0.052462783488009326, 32'sd-0.026872838999100788, 32'sd-0.12098520644009353, 32'sd-0.05377775040457659, 32'sd-0.13550788860224797, 32'sd-0.10837780565952063, 32'sd-0.1655266166093338, 32'sd-0.004541594252736292, 32'sd-0.03524894682357966, 32'sd0.13700017892619928, 32'sd0.09193981323533229, 32'sd0.10241365550044143, 32'sd0.04396629531875377, 32'sd0.04953071001228952, 32'sd0.04460907962324177, 32'sd0.04862747871272898, 32'sd-2.3760961628370488e-122, 32'sd0.028709392720083066, 32'sd0.04678382621303726, 32'sd0.02573169769629483, 32'sd-0.08752702028389248, 32'sd-0.06797679796781263, 32'sd0.12406147761818798, 32'sd0.06328094144964284, 32'sd-0.022432427062224095, 32'sd-0.05451565376487725, 32'sd-0.09534386298464226, 32'sd-0.12772486400143834, 32'sd-0.008758478328347762, 32'sd-0.06923262291591091, 32'sd0.05180692232462754, 32'sd-0.07123027700076785, 32'sd-0.12246076493532562, 32'sd-0.07917406753659649, 32'sd0.029552991285032235, 32'sd0.004317355161253212, 32'sd-0.008345294610768514, 32'sd0.04021008555095967, 32'sd0.1316295410339298, 32'sd0.1701975065649439, 32'sd0.0827958360188624, 32'sd0.07013728712452097, 32'sd0.010945985970045952, 32'sd0.06239906609113566, 32'sd-1.1226699435455717e-118, 32'sd0.0612060799044821, 32'sd-0.008845573119465312, 32'sd-0.013730549015456112, 32'sd0.029244201357348384, 32'sd0.0645968192660933, 32'sd0.00606729852150859, 32'sd-0.10248984180247446, 32'sd0.011510339573730748, 32'sd-0.24779365074289728, 32'sd-0.08533630369914763, 32'sd0.03439038999035748, 32'sd-0.01944807826867447, 32'sd-0.006087985269992837, 32'sd0.021599238862578064, 32'sd-0.05819475744885454, 32'sd-0.201525272468417, 32'sd-0.08708157847284262, 32'sd0.0516870615073525, 32'sd-0.07867130004717646, 32'sd0.050778541491042, 32'sd-0.0258891812575817, 32'sd0.006473794891080467, 32'sd0.12722029853905706, 32'sd0.07899141245160207, 32'sd0.04811979017438796, 32'sd-0.0806417316838082, 32'sd0.007037931466851403, 32'sd0.06109357113116166, 32'sd-0.004082717875820084, 32'sd-0.0018990313099755101, 32'sd0.023945306954971313, 32'sd0.0011116482458624916, 32'sd0.13277789256147499, 32'sd-0.11437715327010377, 32'sd-0.019770535058471043, 32'sd-0.022447547836959438, 32'sd-0.16054951637199574, 32'sd-0.027340435465494, 32'sd0.07395367507492011, 32'sd0.08386921239675758, 32'sd0.0987825728500471, 32'sd0.02695063922996735, 32'sd-0.0652101757858145, 32'sd-0.14832421656824382, 32'sd-0.02456672023093355, 32'sd-0.016384613883124986, 32'sd0.003298020455664609, 32'sd-0.15549892520816277, 32'sd-0.1853983393259743, 32'sd-0.01787096908661552, 32'sd-0.017873857713539932, 32'sd-0.027761273068023652, 32'sd-0.03799874265424151, 32'sd0.008541132828020251, 32'sd0.03618250344773691, 32'sd0.07795912272714915, 32'sd-0.05009516693329351, 32'sd-0.01704450660796878, 32'sd0.06674934728700292, 32'sd0.06799480287479713, 32'sd-0.08124316239170919, 32'sd0.007142331640717556, 32'sd-0.044120890950538706, 32'sd-0.16305933990105062, 32'sd-0.15346251476541525, 32'sd-0.019652223705086715, 32'sd-0.07454437443124186, 32'sd0.0861189187411103, 32'sd0.067231687974918, 32'sd0.015067479474200108, 32'sd-0.1918011913001384, 32'sd-0.18686511223475222, 32'sd-0.15366413461015688, 32'sd-0.035381091440461004, 32'sd-0.098681514035587, 32'sd-0.0797584901554638, 32'sd-0.012212743470755471, 32'sd-0.015890946482639084, 32'sd-0.046765205937256034, 32'sd0.025779661654030568, 32'sd0.06876055602525737, 32'sd0.0027345499818602834, 32'sd0.03634019234332846, 32'sd-0.009441902412561855, 32'sd0.003431490165585811, 32'sd-0.08732751768483923, 32'sd0.053825938551014356, 32'sd-0.045170203803172215, 32'sd-0.05922069750068804, 32'sd-0.05660031362401702, 32'sd-0.05349900948501639, 32'sd-0.14257922055723493, 32'sd-0.052111575698895275, 32'sd-0.20018814856408795, 32'sd0.06636360677904996, 32'sd0.052233009059355635, 32'sd0.11009295886857427, 32'sd-0.016936774498565458, 32'sd-0.20744007136154394, 32'sd-0.12327553293009633, 32'sd-0.0042760490343507086, 32'sd-0.007771478122493507, 32'sd0.053227716366980836, 32'sd-0.034568152536082065, 32'sd-0.08070931497243039, 32'sd-0.00033035183561178674, 32'sd-0.016719289454504283, 32'sd-0.028522614406373163, 32'sd-0.07020272170895676, 32'sd-0.005934068561365593, 32'sd-0.05602011457646739, 32'sd0.06453650911073455, 32'sd0.13216668950487961, 32'sd-0.01423627987123168, 32'sd-0.07985629403586454, 32'sd-0.06368100263003494, 32'sd0.02792544045981682, 32'sd-0.15441574959659726, 32'sd-0.2185015254103824, 32'sd-0.13441211919330065, 32'sd0.012547433393175185, 32'sd-0.19969326368054346, 32'sd-0.09425123495667079, 32'sd0.014262670873501587, 32'sd-0.0846475036109855, 32'sd0.0673227203417052, 32'sd-0.07570306554572079, 32'sd0.0340211497259906, 32'sd0.11444547901660046, 32'sd0.002134064414906699, 32'sd0.12900828430904007, 32'sd0.016728705994307064, 32'sd0.03453256253376213, 32'sd0.09237686437158232, 32'sd0.01638428566458116, 32'sd0.05352085860041831, 32'sd-0.06937640501082279, 32'sd-0.06376393862704292, 32'sd0.03011403092440056, 32'sd0.10003951936541532, 32'sd0.07222660148596033, 32'sd-0.013875158269623761, 32'sd0.012030385657719286, 32'sd0.006351293242344268, 32'sd-0.0812966846462663, 32'sd-0.1616427989753775, 32'sd-0.07913664792191816, 32'sd0.002562800805228916, 32'sd0.03117084140069485, 32'sd-0.04039699664064228, 32'sd-0.058198594455973696, 32'sd0.07778060734345656, 32'sd0.07478383939562719, 32'sd0.05126416427612583, 32'sd-0.03160174964757126, 32'sd0.17512594236431206, 32'sd0.11597421784451407, 32'sd0.20786885980658926, 32'sd0.1375545934161532, 32'sd0.01634010480755878, 32'sd-0.03497933091272922, 32'sd0.10281583589899425, 32'sd0.17391022740879056, 32'sd0.09796740183742902, 32'sd-0.03356201751336491, 32'sd0.0771885980089588, 32'sd-0.11304389656248161, 32'sd-0.0002696675239729839, 32'sd0.03544619762442668, 32'sd-0.06984018199143512, 32'sd0.015490515434804283, 32'sd0.02481106188249529, 32'sd0.023302041956440558, 32'sd-0.149102918610664, 32'sd0.0056555103484677745, 32'sd0.06280952795011303, 32'sd0.0910513857534123, 32'sd-0.004835119040277275, 32'sd0.016315720916864295, 32'sd-0.025414763613783756, 32'sd0.1394972041455807, 32'sd0.24292335088409556, 32'sd0.07612927585816726, 32'sd0.001607790727476704, 32'sd0.10553417998493132, 32'sd0.0965528281082482, 32'sd0.16557586304674246, 32'sd0.07599802863231916, 32'sd0.11513278040590344, 32'sd0.151867372759669, 32'sd0.06198768634516175, 32'sd0.07984093409513765, 32'sd-0.03853833002057503, 32'sd0.07949626899385312, 32'sd0.031616688175622396, 32'sd0.021779166266558576, 32'sd-0.019520723662111772, 32'sd0.07979633557085448, 32'sd-0.007771018874330505, 32'sd-0.02508213376878027, 32'sd-0.08390737332159788, 32'sd-0.010443084999297568, 32'sd-0.04302233265076964, 32'sd0.033175827347153956, 32'sd0.050465924484883205, 32'sd0.10644413268308203, 32'sd0.17469949928184114, 32'sd0.13348324755472443, 32'sd0.19477568456501726, 32'sd0.1384714146861275, 32'sd0.032445692351197895, 32'sd-0.014029137072467238, 32'sd0.058553673489325817, 32'sd-0.03967571997257345, 32'sd0.08322461620233727, 32'sd0.04759307306470719, 32'sd0.09621432825995577, 32'sd-0.012876692712545802, 32'sd0.017530111034575392, 32'sd-0.036166275676566, 32'sd-0.012586016367183924, 32'sd-0.02359274285290996, 32'sd-0.004869424331186545, 32'sd0.07513915189603976, 32'sd0.013886211839091937, 32'sd-0.07893903033327035, 32'sd0.08772271073120791, 32'sd0.026370812260630743, 32'sd-0.0047583937562480924, 32'sd-0.17995813996205362, 32'sd0.003724035359754402, 32'sd-0.0015090770897999133, 32'sd0.15387356524329623, 32'sd0.1529511856033929, 32'sd0.12013124686575563, 32'sd0.018438385657469223, 32'sd0.12967606981434474, 32'sd0.04286276696560713, 32'sd0.029080091186700845, 32'sd0.08803468323057433, 32'sd0.07608207481947717, 32'sd-0.0032568245226171676, 32'sd0.04289123027977074, 32'sd0.10747624370237013, 32'sd0.0212600493264201, 32'sd-0.08253559080568221, 32'sd-0.16268033512338015, 32'sd-0.05390007233213065, 32'sd-0.14036027442089266, 32'sd-0.026387995617145176, 32'sd-0.02388009742732712, 32'sd-0.0030570691059717404, 32'sd0.056289446495723996, 32'sd-0.045245395971488155, 32'sd0.00984086646482958, 32'sd0.05619713753253577, 32'sd-0.055853468856663036, 32'sd-0.0848691625194346, 32'sd0.028806438805632134, 32'sd0.11883250603227485, 32'sd0.07415460253716147, 32'sd0.07014283715911057, 32'sd0.03134205346961518, 32'sd0.06866353918679546, 32'sd-0.03691513275544498, 32'sd0.1342171152056388, 32'sd0.08122208179836972, 32'sd-0.010036972288120637, 32'sd0.05217272125186896, 32'sd-0.025366283909506057, 32'sd-0.019560038321147846, 32'sd-0.14604533303976877, 32'sd-0.0066682515059047235, 32'sd-0.07840403953727387, 32'sd-0.08221678968286047, 32'sd-0.03436231515889819, 32'sd-0.009299063080961208, 32'sd-0.07825287469425814, 32'sd-0.024683980006714137, 32'sd0.06614692097929398, 32'sd0.03579560004508751, 32'sd-0.01577993777331421, 32'sd-0.004298063998010767, 32'sd0.06204292318818279, 32'sd-0.01625689430642654, 32'sd-0.09235931192171039, 32'sd-0.115073407585406, 32'sd0.06065549697402052, 32'sd-0.03966772763350507, 32'sd0.033593673908443054, 32'sd-0.05598178376934747, 32'sd-0.0026429749925271154, 32'sd0.03125066815006827, 32'sd0.020679034183340054, 32'sd0.026139392258629178, 32'sd-0.10848756786453785, 32'sd0.08764932582982905, 32'sd0.007242487595742555, 32'sd-0.10616485310795921, 32'sd-0.07779833849070437, 32'sd-0.103050064774812, 32'sd-0.09035972630733077, 32'sd-0.14331268123220547, 32'sd-0.101525014914522, 32'sd-0.0877314856862406, 32'sd0.010352051655397279, 32'sd0.04401168349297854, 32'sd-5.152814672680376e-117, 32'sd-0.0020654551271299688, 32'sd-0.07491576957212795, 32'sd-0.011411620474358085, 32'sd0.12098273903396159, 32'sd-0.06758103702735944, 32'sd-0.0375640930470198, 32'sd-0.12011438666788521, 32'sd-0.009620258471847797, 32'sd-0.06850598522527696, 32'sd0.07015952787863766, 32'sd-0.012681064417371053, 32'sd0.05558035501925038, 32'sd-0.02714503992096046, 32'sd0.036222562256472066, 32'sd-0.054456973918349666, 32'sd-0.06951184052962021, 32'sd-0.002305307555467929, 32'sd-0.012621734987825947, 32'sd-0.02135598088447405, 32'sd-0.018876132636251694, 32'sd-0.11603537956053572, 32'sd-0.08941246509362433, 32'sd-0.0835896537879344, 32'sd-0.09690258219432392, 32'sd-0.001309205908801989, 32'sd0.023558206717300578, 32'sd-0.09413419483984263, 32'sd-0.04279994975488385, 32'sd0.0366158441894041, 32'sd-0.11396799333073983, 32'sd-0.024497783269444882, 32'sd0.004561847691186883, 32'sd-0.08097632835183244, 32'sd-0.07362480682260182, 32'sd-0.035521069471030356, 32'sd-0.03074039438841904, 32'sd-0.04589513775339759, 32'sd0.11982587500213912, 32'sd0.15466010152621518, 32'sd0.087759491623372, 32'sd-0.10854474791415938, 32'sd-0.09459854750415975, 32'sd-0.10075775214096722, 32'sd-0.05974791438623886, 32'sd0.05939432750310679, 32'sd-0.0900465206851746, 32'sd-0.05713939716876162, 32'sd-0.0391071838957559, 32'sd-0.02351116379438313, 32'sd-0.20171317246192064, 32'sd-0.1795121356092076, 32'sd-0.15205364501089544, 32'sd-0.04397265060214691, 32'sd0.08049942788203747, 32'sd0.02710545457145401, 32'sd0.03855425858339551, 32'sd0.018234949415262967, 32'sd-0.07811063490566111, 32'sd-0.1365126351814797, 32'sd-0.11649433657958601, 32'sd0.07426941901938786, 32'sd-0.08387873830028532, 32'sd0.03159772828933903, 32'sd-0.05917333558059941, 32'sd0.032120075565661065, 32'sd0.11849564426249067, 32'sd0.058709381493303986, 32'sd0.03843196604945669, 32'sd-0.006717564470001962, 32'sd-0.03463075240600095, 32'sd-0.0390501964751639, 32'sd-0.02658854409311858, 32'sd0.026639224651208708, 32'sd0.028838863063500052, 32'sd-0.12877891181717496, 32'sd-0.12252283315043727, 32'sd-0.08570516278037946, 32'sd-0.17747853668001481, 32'sd-0.09689275885645669, 32'sd-0.08818212284394202, 32'sd-0.044560566590681305, 32'sd0.05806863253681589, 32'sd-0.08477374679691531, 32'sd5.429002142522299e-121, 32'sd-0.0018722442747958945, 32'sd0.08946292023772208, 32'sd-0.17315593587867836, 32'sd-0.06341469683607462, 32'sd-0.15412207133415154, 32'sd-0.02784507083219673, 32'sd-0.0742640912230705, 32'sd-0.07845101722935574, 32'sd0.005915475307336566, 32'sd0.04634235557598827, 32'sd0.035980562832378556, 32'sd-0.05808354141657051, 32'sd0.028363387748070044, 32'sd-0.0663598802533275, 32'sd0.0740457976673765, 32'sd-0.02509763987606117, 32'sd0.002551225364537776, 32'sd-0.05303704817690105, 32'sd-0.06501101172676163, 32'sd-0.14015416294668326, 32'sd-0.19888189273735377, 32'sd-0.10341727705257912, 32'sd-0.17532648451657615, 32'sd-0.11902135197720232, 32'sd0.06042951501476846, 32'sd0.0825319951261946, 32'sd0.06288579324845599, 32'sd0.08890863797881585, 32'sd-0.004062562417788922, 32'sd0.04513678518580887, 32'sd-0.011714083326724307, 32'sd-0.08408858663756573, 32'sd-0.039817228009679545, 32'sd-0.09595663990705844, 32'sd0.06907477868440809, 32'sd-0.05368177565883144, 32'sd0.10003988635055472, 32'sd-0.10157874465768527, 32'sd-0.0806593689172739, 32'sd-0.0028243389109250338, 32'sd0.008781652916247459, 32'sd-0.09072865182840469, 32'sd0.0014069522705523283, 32'sd-0.07501078978692774, 32'sd-0.036375801260839245, 32'sd-0.1026992608608654, 32'sd-0.19508631238601948, 32'sd-0.07672121220997653, 32'sd-0.10637577586561724, 32'sd-0.017545130729633852, 32'sd-0.06231660108824916, 32'sd-0.008579225668239633, 32'sd0.045136001236838155, 32'sd0.03548314853981322, 32'sd0.06905038770022069, 32'sd-0.013859001549428705, 32'sd0.05318647557446413, 32'sd0.05147826691194975, 32'sd0.0036408119274381544, 32'sd-0.09375472295180683, 32'sd-0.08587333349894728, 32'sd0.033424881978091806, 32'sd-0.015801897499300877, 32'sd0.06850598009756131, 32'sd0.0555478112413428, 32'sd0.03222196647650475, 32'sd0.018574178716319563, 32'sd0.05234647856371565, 32'sd0.02952676408529954, 32'sd0.04686591501188707, 32'sd-0.13326880729033344, 32'sd-0.2471535110990998, 32'sd-0.2559332955907199, 32'sd-0.1742732156761265, 32'sd-0.05208083112536876, 32'sd-0.1474908308005144, 32'sd-0.0880494623102296, 32'sd0.02761003678912725, 32'sd-0.10998219143769444, 32'sd-0.083911276065957, 32'sd-0.02382976204368494, 32'sd0.009356012266298884, 32'sd0.05271663694888515, 32'sd-3.810944920281064e-127, 32'sd-0.003489826828858259, 32'sd0.0010599563665058306, 32'sd-0.04729289762387922, 32'sd-0.09809688209926402, 32'sd-0.041383015909816086, 32'sd-0.06722491102196436, 32'sd-0.05428413777387804, 32'sd0.17196151724257572, 32'sd0.003855385330356534, 32'sd0.009515058984604556, 32'sd0.00492005811407597, 32'sd-0.057049991895224375, 32'sd-0.10943939173256292, 32'sd-0.07690678891939033, 32'sd-0.22743673899264508, 32'sd-0.025043394897395373, 32'sd-0.16438735504222451, 32'sd-0.07079696281857951, 32'sd-0.05275012290145134, 32'sd-0.12348168971366014, 32'sd-0.10123763983140904, 32'sd-0.01973718609602397, 32'sd0.019987589929141302, 32'sd-0.03158526950430524, 32'sd0.03144646314513201, 32'sd-0.07465466994025259, 32'sd-7.375937566492678e-121, 32'sd-1.193309632112298e-115, 32'sd1.1602353200427726e-123, 32'sd-0.00409797444480639, 32'sd-0.027991486815430268, 32'sd0.06678635467599915, 32'sd0.025473618679678307, 32'sd-0.03641561730086706, 32'sd-0.02179037929332206, 32'sd0.06015950190726592, 32'sd0.01474536444659939, 32'sd-0.009583221359470049, 32'sd0.02822874270175495, 32'sd-0.02192753709725245, 32'sd-0.019288549356268617, 32'sd0.064294495451205, 32'sd-0.06912181897094344, 32'sd0.12915949989365236, 32'sd-0.08607808926913464, 32'sd-0.15149077507209047, 32'sd-0.027528691011324116, 32'sd-0.06779818210772187, 32'sd0.048734847641988537, 32'sd0.00505016671905781, 32'sd-0.029720483058120552, 32'sd-0.04712165249930548, 32'sd-0.007677244532783203, 32'sd0.005758459469451951, 32'sd3.4247086366834956e-117, 32'sd-8.643573643478284e-127, 32'sd1.5763584624124063e-127, 32'sd0.03329817712944634, 32'sd-0.11169892580147493, 32'sd0.00785978761018324, 32'sd-0.04656185786361724, 32'sd-0.004928300374034834, 32'sd0.047820450122708975, 32'sd0.021819228168130415, 32'sd0.0034445089431520393, 32'sd-0.04948304727048186, 32'sd0.04207560034640725, 32'sd-0.11762298088996209, 32'sd-0.03679412903356917, 32'sd-0.0753634509360748, 32'sd-0.025262934186428162, 32'sd-0.05623762821812266, 32'sd-0.15325697685432843, 32'sd0.016289391662040163, 32'sd0.05015018745802741, 32'sd0.029948655124976575, 32'sd0.0005064232634699982, 32'sd-0.12578009873464752, 32'sd-0.035956374098504544, 32'sd-0.043492859883778566, 32'sd-0.021169635964213254, 32'sd-0.0006540099572525373, 32'sd5.854072826598539e-122, 32'sd1.9158547295806315e-117, 32'sd9.3305728653855e-126, 32'sd4.321810883998017e-125, 32'sd0.062078995071840386, 32'sd0.0856715318910002, 32'sd-0.046292031367605055, 32'sd-0.004735536569971476, 32'sd-0.006456541983242143, 32'sd0.011727820335935418, 32'sd-0.12179623298516835, 32'sd-0.06966836924660512, 32'sd0.18844740629464737, 32'sd-0.011815207064456603, 32'sd0.06258140630880508, 32'sd0.028271771560370116, 32'sd-0.026957806341837205, 32'sd-0.0177094172406124, 32'sd-0.07835600743803989, 32'sd0.05176971146060044, 32'sd-0.0019053500708226783, 32'sd0.044621232418518536, 32'sd-0.03966059509066625, 32'sd0.01869214265374626, 32'sd0.0294223740630484, 32'sd-0.0295632123455196, 32'sd0.004102845513941222, 32'sd-6.957937249030591e-115, 32'sd-2.1185345184511123e-126, 32'sd-1.4341567811807796e-118, 32'sd-2.8183343359704794e-118, 32'sd-1.0700811891939414e-121, 32'sd2.3336444124090884e-122, 32'sd0.017183058325099625, 32'sd0.021204692745286018, 32'sd-0.02323945779141246, 32'sd-0.02378878746823246, 32'sd-0.06258188631578532, 32'sd0.012157402259950647, 32'sd0.024416621712318495, 32'sd0.03927085377384649, 32'sd-0.045724934601506464, 32'sd0.06852871171906982, 32'sd0.047119996256500346, 32'sd0.06625949953769325, 32'sd0.012580903385469196, 32'sd0.01241782375623558, 32'sd0.055744408188217784, 32'sd-0.07020003194796197, 32'sd-0.07999717773668005, 32'sd-0.04861546149649887, 32'sd-0.016593368819599344, 32'sd-1.5178030967986902e-05, 32'sd1.2855871616539872e-118, 32'sd-8.211406329610435e-117, 32'sd1.7814033805651254e-124, 32'sd1.1651138745105461e-123},
        '{32'sd1.255850949353193e-125, 32'sd1.3292955217656762e-117, 32'sd1.516070341275775e-120, 32'sd-9.103591132903175e-118, 32'sd-5.8001719479874725e-124, 32'sd-1.0485603449437317e-122, 32'sd1.3228791711616298e-122, 32'sd-3.976918376533627e-125, 32'sd3.483047621744016e-125, 32'sd-1.7687335786452271e-124, 32'sd-4.793542963134236e-123, 32'sd1.380366787507871e-115, 32'sd-0.07232857998302149, 32'sd-0.07962002566235289, 32'sd0.022277060776497947, 32'sd-0.029832055833396164, 32'sd6.748951582143762e-124, 32'sd3.1207987316159305e-120, 32'sd-6.6833000597396675e-124, 32'sd-9.140264458853205e-125, 32'sd8.762660929767682e-123, 32'sd-4.167841119668723e-122, 32'sd-1.8946897384498585e-120, 32'sd1.6733471164699893e-126, 32'sd-3.649547119055142e-116, 32'sd5.4591980853221075e-126, 32'sd3.270080871444071e-124, 32'sd8.128795672456543e-121, 32'sd-7.894850431868351e-122, 32'sd3.340382332113984e-120, 32'sd6.893048927893795e-126, 32'sd-1.5962626610758354e-124, 32'sd0.01126275424570601, 32'sd-0.03819385395510879, 32'sd0.045711710684902915, 32'sd-0.09434908782763117, 32'sd-0.03616754693020073, 32'sd0.018410391941955456, 32'sd0.07723481612323502, 32'sd0.003876072636472987, 32'sd-0.04341848136241427, 32'sd0.029589031439721244, 32'sd-0.026911504931464308, 32'sd0.014352572817729958, 32'sd-0.013877748110597693, 32'sd0.013042089498378671, 32'sd0.01973740635824383, 32'sd0.045790775973833305, 32'sd0.05627809521018564, 32'sd0.06222100792754803, 32'sd0.04604587506839382, 32'sd0.010599868722558189, 32'sd-2.9833417672233782e-124, 32'sd4.5271099319843975e-115, 32'sd5.8820947166348335e-118, 32'sd-1.1468074739936546e-115, 32'sd3.68287114940576e-129, 32'sd5.419141918512907e-125, 32'sd0.045210349101999024, 32'sd0.047505845044285726, 32'sd0.010289688026357333, 32'sd0.0015700536856676794, 32'sd0.002786168116476882, 32'sd-0.020010326644497894, 32'sd-0.06348420839997329, 32'sd-0.0371057738985727, 32'sd0.07939389600840618, 32'sd0.08306515701752341, 32'sd-0.08021632396748278, 32'sd0.017680329836129324, 32'sd-0.06675944699107005, 32'sd0.0014112909227006068, 32'sd-0.026480069893455468, 32'sd0.1820444943204797, 32'sd0.06628580813024561, 32'sd0.1042950582199448, 32'sd-0.004708331802544059, 32'sd0.09643743294895518, 32'sd0.027473486080042547, 32'sd-0.009043987655931677, 32'sd0.06057149888772216, 32'sd0.03354189824552894, 32'sd2.1129530460251725e-123, 32'sd-1.6311845584932066e-115, 32'sd-2.4364014407626376e-124, 32'sd-1.4009406812875875e-115, 32'sd0.05571355911522724, 32'sd0.005125369471708996, 32'sd0.05130738615753838, 32'sd-0.016102373133598843, 32'sd0.05351107937854521, 32'sd0.06405292689734012, 32'sd0.0025064781160134934, 32'sd0.11966585342376747, 32'sd0.014038783858628924, 32'sd-0.1261353184598831, 32'sd-0.09135159899592525, 32'sd-0.01427575636327751, 32'sd-0.07002979461909915, 32'sd-0.10061274055922537, 32'sd-0.07979357695466509, 32'sd0.1586577779683412, 32'sd0.07788980548688838, 32'sd0.15967287606573302, 32'sd-0.029068206546794827, 32'sd-0.04254950641584571, 32'sd-0.04469397144752754, 32'sd-0.0017977010458376447, 32'sd0.005170931922616209, 32'sd-0.01832141376810388, 32'sd-0.056768165225519994, 32'sd1.6374192640853387e-120, 32'sd2.0962558673567776e-126, 32'sd0.040808912136350926, 32'sd0.07666856100387132, 32'sd-0.03589726480299879, 32'sd-0.09628925487424067, 32'sd0.0388061753806693, 32'sd-0.07244662073800201, 32'sd-0.020990871764194927, 32'sd0.03481644989602495, 32'sd0.012343054186842454, 32'sd-0.11308027678859181, 32'sd0.010061200736856441, 32'sd0.06304305066700826, 32'sd-0.017129742928351312, 32'sd-0.11290545385211379, 32'sd-0.09699681586227629, 32'sd0.020237358845823623, 32'sd0.17256591685047806, 32'sd0.11117906928319174, 32'sd0.07279008112439483, 32'sd-0.10275861602042773, 32'sd-0.16867444336610718, 32'sd-0.13920595630748217, 32'sd-0.1188807675936274, 32'sd0.03507576145486238, 32'sd0.017558265593973225, 32'sd-0.05634369853510965, 32'sd-0.02375156567884053, 32'sd6.619342694124679e-126, 32'sd-0.010136825708750305, 32'sd0.08742065022031088, 32'sd-0.06564841197220529, 32'sd0.012041699945114786, 32'sd-0.05353145547551516, 32'sd-0.12656542968156254, 32'sd-0.04522883502538962, 32'sd-0.14728090442133834, 32'sd-0.17595311909450082, 32'sd-0.15814340369025545, 32'sd-0.10129471447599686, 32'sd-0.12999016582942613, 32'sd-0.037917162734309395, 32'sd0.03794895904132373, 32'sd0.12254865230760344, 32'sd0.13592594110611278, 32'sd0.06482444168290291, 32'sd0.044596554177787344, 32'sd0.061056355506802294, 32'sd-0.008594616598818083, 32'sd-0.13548356877016157, 32'sd-0.13278868896691193, 32'sd-0.06415269355992992, 32'sd0.004647265274082422, 32'sd0.007703384427634959, 32'sd0.04676541940703706, 32'sd0.06087088985987201, 32'sd1.63787007290834e-123, 32'sd-0.010797950984570684, 32'sd0.03757578380728815, 32'sd-0.030407385524325998, 32'sd-0.051289666291669825, 32'sd-0.014109459716416053, 32'sd-0.07539949072047875, 32'sd-0.08962399589295333, 32'sd-0.05977025720023501, 32'sd-0.2583733829803902, 32'sd-0.17403336054789625, 32'sd0.01860021084554778, 32'sd-0.011002729810712349, 32'sd0.057752221934949645, 32'sd0.17752161734752986, 32'sd0.08467091366450805, 32'sd0.05766794955262119, 32'sd-0.06596135357489918, 32'sd-0.031993292212151477, 32'sd-0.018907510693833948, 32'sd-0.1365990495553782, 32'sd-0.1260534826023483, 32'sd0.00044630743342107736, 32'sd0.013283873817184428, 32'sd-0.09815951898756207, 32'sd-0.04885349801854105, 32'sd-0.009794672221036907, 32'sd-0.014865366481419527, 32'sd0.016014723314337703, 32'sd-0.006811025637921545, 32'sd-0.044751407630551764, 32'sd-0.016463048995057034, 32'sd-0.03069649786258326, 32'sd-0.05158508712259567, 32'sd-0.21349930777979664, 32'sd-0.2327904915718274, 32'sd-0.18897273906951345, 32'sd-0.16779155731091877, 32'sd-0.045069085052824, 32'sd0.14080434838238615, 32'sd0.14471550551581677, 32'sd0.1677558541311763, 32'sd0.04955231012615757, 32'sd-0.005416592814219762, 32'sd-0.0378121697100976, 32'sd-0.08399312643128799, 32'sd-0.11521281618539708, 32'sd-0.14062989209195664, 32'sd-0.12902048269894187, 32'sd-0.09428801964914295, 32'sd0.12470700142838215, 32'sd-0.08570733029588624, 32'sd-0.019089631537429645, 32'sd-0.03406780276446392, 32'sd0.10081134400286741, 32'sd0.03925245262109671, 32'sd0.00999195112210817, 32'sd-0.03884998671983982, 32'sd-0.008744627473627692, 32'sd-0.021228945600151813, 32'sd-0.1039130521066274, 32'sd-0.11039778047803707, 32'sd-0.21358321265117758, 32'sd-0.19496130219651878, 32'sd-0.14457572737578533, 32'sd-0.1778570565050166, 32'sd-0.061650933548510846, 32'sd0.07930967609692459, 32'sd0.20448334205196764, 32'sd0.055409536810087374, 32'sd-0.07738981691428141, 32'sd-0.11845989556532037, 32'sd-0.12792122215085625, 32'sd-0.07821122835261246, 32'sd-0.09424084744273788, 32'sd-0.0022076978823684554, 32'sd-0.10927273550414716, 32'sd-0.003873856312586658, 32'sd0.02090412288311217, 32'sd0.03408224600266018, 32'sd0.09744855583905407, 32'sd0.22035705263196362, 32'sd0.025242051382205626, 32'sd0.08667327404849841, 32'sd-0.010009303560054876, 32'sd-0.06845538740016271, 32'sd0.09814633668918184, 32'sd-0.04576080923256461, 32'sd-0.1421529312885252, 32'sd-0.2112230087594268, 32'sd-0.03778560260710611, 32'sd-0.15731333265654518, 32'sd0.0021961762127835362, 32'sd-0.04024070119644898, 32'sd0.043919250184053085, 32'sd0.19975239557597851, 32'sd0.12885229379604607, 32'sd0.05572449730556969, 32'sd-0.08605170291778248, 32'sd-0.1035915123671577, 32'sd0.0024945187499671065, 32'sd-0.010060182640100584, 32'sd-0.11184298835658035, 32'sd0.10375382161558189, 32'sd-0.0849360974966729, 32'sd0.005123142645272098, 32'sd0.034729867748650056, 32'sd0.06779179942295024, 32'sd0.0657709881222849, 32'sd0.03698384816294851, 32'sd0.06366762807527207, 32'sd0.0761203086593009, 32'sd-0.0666103154180006, 32'sd-0.011102392897317837, 32'sd0.09733363625319882, 32'sd0.01559616151610162, 32'sd-0.007375533004901778, 32'sd-0.0983709568225622, 32'sd-0.1488386176756785, 32'sd-0.08332444900049799, 32'sd0.07035990192641509, 32'sd-0.07845898333659411, 32'sd-0.04706852552977491, 32'sd-0.04234061175174789, 32'sd-0.016744086990585882, 32'sd-0.0036223340698009893, 32'sd0.013808402047364898, 32'sd0.01945061403205014, 32'sd-0.09658133078102404, 32'sd-0.016204768710364952, 32'sd0.056311061818763615, 32'sd0.1506560539647275, 32'sd0.06459624258345274, 32'sd0.17289523464301898, 32'sd0.02068020132148941, 32'sd0.10502781962002222, 32'sd0.05887225686113125, 32'sd0.08530220299970588, 32'sd0.07745402619804745, 32'sd-0.07584155750219777, 32'sd-0.010700451650594026, 32'sd-0.002593788267667755, 32'sd-0.0007454430418777543, 32'sd-0.05045982205421945, 32'sd-0.04136737712826952, 32'sd-0.06372882307674854, 32'sd-0.05932895754138758, 32'sd-0.03552186959451402, 32'sd-0.019994601851411904, 32'sd-0.01623345612354265, 32'sd-0.02734887233448983, 32'sd-0.0538494595238573, 32'sd-0.048900631446950525, 32'sd0.07738851753839486, 32'sd0.020647312811568126, 32'sd0.0043091393179913, 32'sd0.05545876394132952, 32'sd0.01826880027534463, 32'sd0.014761669601285835, 32'sd0.03326694588286888, 32'sd0.018358217308666255, 32'sd0.01438136375080849, 32'sd0.051832192837487696, 32'sd0.02854231787109227, 32'sd0.07198757508331582, 32'sd0.016594562568005757, 32'sd-0.02631732503146473, 32'sd0.04712368057659011, 32'sd0.05869676225254883, 32'sd0.03458937939630315, 32'sd0.04820844247718293, 32'sd-0.03693550396849189, 32'sd-0.10695538971544791, 32'sd0.002026336432459091, 32'sd0.03260270651370334, 32'sd0.05543902104194651, 32'sd-0.020940051696780752, 32'sd0.025308724423709905, 32'sd0.051312856587460105, 32'sd0.19124661268044627, 32'sd0.1101270358652603, 32'sd0.04421550538900015, 32'sd0.08828383414726301, 32'sd0.008349579385865474, 32'sd-0.05597788993601943, 32'sd0.00329761308937855, 32'sd-0.11504284366220939, 32'sd0.033527660281592694, 32'sd0.06827382900326781, 32'sd0.026335996446444573, 32'sd0.08419268506994881, 32'sd-0.012272808161813623, 32'sd-0.03517025318186486, 32'sd0.07421703397567479, 32'sd0.0353134091047037, 32'sd-0.026592360889287795, 32'sd-0.003758244514732813, 32'sd-0.031104783618881002, 32'sd-0.08476475189664427, 32'sd0.05593699999179683, 32'sd-0.0692337402882509, 32'sd-0.05690380832114098, 32'sd-0.05780672881738197, 32'sd0.004736221016314889, 32'sd0.03251826217338269, 32'sd0.16216750543063052, 32'sd-0.002513584511740523, 32'sd0.0652778697147567, 32'sd0.14915430801748059, 32'sd0.008035522641459137, 32'sd-0.004644109778771978, 32'sd-0.068362696100961, 32'sd-0.10132767860066848, 32'sd-0.04467457725344792, 32'sd-0.19897268562114326, 32'sd0.04435589533140841, 32'sd-0.10635168397182075, 32'sd-0.06550189278259871, 32'sd0.028856477179577556, 32'sd-0.07129167908191385, 32'sd-0.11337652414931497, 32'sd-0.06719924069499784, 32'sd-0.00021132114948038994, 32'sd0.03819135075850173, 32'sd0.12018978763322453, 32'sd0.013363664401503918, 32'sd-0.02950474191185538, 32'sd0.07272284000400431, 32'sd0.015483809700121316, 32'sd-0.11581052111461443, 32'sd-0.11758410480755155, 32'sd-0.014795072432318254, 32'sd0.022701048917980155, 32'sd0.14105455981955167, 32'sd0.07088435679729213, 32'sd0.07175945253967496, 32'sd0.13588022298789978, 32'sd-0.03585336208518617, 32'sd-0.1283853766225522, 32'sd-0.06371014404660545, 32'sd0.01583520128784556, 32'sd0.03825785794547487, 32'sd-0.16385611728488927, 32'sd-0.17536570798599785, 32'sd-0.09802571150966924, 32'sd0.03311025254390735, 32'sd0.1773485528357599, 32'sd-0.011161791348194405, 32'sd-0.007826080805807838, 32'sd-0.05418220605832347, 32'sd-0.0210196866185741, 32'sd0.0606951937450745, 32'sd0.05006684099267791, 32'sd0.05140219905337262, 32'sd-0.02369451681593659, 32'sd0.13521959524083688, 32'sd0.07674921897495539, 32'sd0.04824863207704593, 32'sd0.01424066934745599, 32'sd0.02953550127616241, 32'sd0.08217269426807469, 32'sd0.12460046237129072, 32'sd0.022878284541436554, 32'sd0.032392641068047914, 32'sd-0.03792050427752698, 32'sd-0.06665797791026012, 32'sd-0.06193256567251501, 32'sd0.08080928254125888, 32'sd0.09488696776993055, 32'sd-0.08466148819261991, 32'sd-0.11026662285433363, 32'sd-0.10759994575809208, 32'sd0.020639943027250834, 32'sd0.10476598060621425, 32'sd-0.021753778523693937, 32'sd-0.027785395313786633, 32'sd-0.06995083246251368, 32'sd-0.04918459351794189, 32'sd-0.01132304756777821, 32'sd0.014887994589498835, 32'sd-0.0014975962671174175, 32'sd-0.06713686521419521, 32'sd0.0003395100775303854, 32'sd0.012170560412975876, 32'sd0.039171320261866746, 32'sd-0.026120866008645077, 32'sd-0.09309415367431194, 32'sd-0.1317620017384196, 32'sd0.06792312650175787, 32'sd-0.03080386918294998, 32'sd0.10703920189305897, 32'sd-0.013832669820081621, 32'sd0.05679278569767564, 32'sd-0.05812299019138857, 32'sd0.06704702149521058, 32'sd0.04016152449231025, 32'sd0.07140996429278369, 32'sd-0.14902836018946394, 32'sd-0.14083131236310611, 32'sd-0.02565661565783635, 32'sd-0.030844396011518907, 32'sd0.01807829655092699, 32'sd-0.06991094674658692, 32'sd-0.03710163599921156, 32'sd-0.03531248882793508, 32'sd-0.020060594675968435, 32'sd0.05871574899839928, 32'sd0.008333210451454548, 32'sd-2.1086282789124877e-122, 32'sd0.08227999322620702, 32'sd0.031206465545277107, 32'sd0.0038292237854859763, 32'sd-0.01089701713117999, 32'sd0.012962537611840824, 32'sd0.0483231659660365, 32'sd-0.055731703684568513, 32'sd-0.054952616275188375, 32'sd-0.15597371891056122, 32'sd0.08604711187672254, 32'sd0.07352380124984248, 32'sd-0.0351495524134247, 32'sd-0.07819577672446576, 32'sd-0.0495064138224158, 32'sd0.1291509450561938, 32'sd0.01029399947735463, 32'sd-0.004525937551712638, 32'sd-0.18923728123143818, 32'sd-0.1103281994442357, 32'sd0.053364107757195245, 32'sd0.02180425233356013, 32'sd0.013516620596743767, 32'sd-0.10405952469649005, 32'sd-0.059135027607844046, 32'sd-0.04553248330160002, 32'sd0.13388384441935022, 32'sd-0.06146455737696224, 32'sd-0.03256042166242154, 32'sd-0.010052535553171144, 32'sd0.05356900740664371, 32'sd-0.06096852088779585, 32'sd0.010201695942991956, 32'sd-0.05335927157060693, 32'sd0.013382719407458705, 32'sd0.005824948697340206, 32'sd-0.07041589314112405, 32'sd-0.11306499771896814, 32'sd-0.10727084744972513, 32'sd-0.16183984832068243, 32'sd0.025319811003374017, 32'sd-0.05968716050095138, 32'sd0.04019646799273221, 32'sd0.1529914332815513, 32'sd0.035932890810537, 32'sd-0.15726643143591162, 32'sd-0.12168624393839508, 32'sd-0.13498917163603835, 32'sd-0.016744239960610516, 32'sd-0.027409114025799437, 32'sd0.008292922332792614, 32'sd-0.01496249054448807, 32'sd-0.03134220291881521, 32'sd0.021256189374682783, 32'sd-0.018471519710577925, 32'sd0.06765702483037121, 32'sd0.004536187888792732, 32'sd0.03570483975408389, 32'sd0.05643250001139204, 32'sd-0.016893132263743307, 32'sd-0.026296049123640877, 32'sd0.0308916897568547, 32'sd-0.0425945918021467, 32'sd-0.00541737385857189, 32'sd-0.025959013262708663, 32'sd-0.11447741981726818, 32'sd-0.029604921613723984, 32'sd-0.020286251442821944, 32'sd-0.04010681366372441, 32'sd-0.03712142106941593, 32'sd0.027222118845825455, 32'sd0.16684566772722562, 32'sd-0.05501018415210784, 32'sd-0.061442493141438966, 32'sd0.06617157832086486, 32'sd-0.09864912680812873, 32'sd0.010796464252348214, 32'sd0.03664888710888654, 32'sd-0.06584486178201886, 32'sd0.06717012877675078, 32'sd-0.011142274863675127, 32'sd-0.049294067821583826, 32'sd0.011531856722924073, 32'sd-0.02852591142914698, 32'sd2.2274378242787153e-114, 32'sd0.01664621669304176, 32'sd-0.035075467800083616, 32'sd0.032436318843987906, 32'sd-0.00486132181420674, 32'sd0.09413406275834338, 32'sd0.061212571671257265, 32'sd-0.09270477869864588, 32'sd-0.17152162629816042, 32'sd-0.06685857123355413, 32'sd0.0035999568800486287, 32'sd0.03618534566315323, 32'sd0.07516325939530571, 32'sd0.024733741408071715, 32'sd-0.043435444099580715, 32'sd0.0739821270535552, 32'sd0.14793108046020953, 32'sd0.07548452685580756, 32'sd0.13096136102046319, 32'sd0.036726426076725445, 32'sd-0.03538761533785265, 32'sd0.001730934209028873, 32'sd0.04485638357069497, 32'sd-0.03487590035877996, 32'sd0.01770685478257046, 32'sd-0.023330935624439334, 32'sd0.03797184305156216, 32'sd-0.02563202360609894, 32'sd0.08029247581043968, 32'sd-0.017413595205859177, 32'sd-0.040817596913406626, 32'sd0.09326185453570777, 32'sd-0.010824798300405373, 32'sd-0.09854109377345102, 32'sd-0.08206803257331127, 32'sd-0.03637535661537311, 32'sd-0.014655614466607255, 32'sd0.11302453399527625, 32'sd-0.020047366960308562, 32'sd0.08416691877060557, 32'sd0.08101168562111143, 32'sd0.10101779982567725, 32'sd0.0389035960264207, 32'sd0.09941675724116834, 32'sd0.03186159251779789, 32'sd0.1081477379170005, 32'sd-0.019209413878483433, 32'sd-0.049019341019144944, 32'sd0.0028955815257564834, 32'sd-0.022703031631396503, 32'sd-0.003685487335169763, 32'sd0.08365138511020467, 32'sd0.055997820848925, 32'sd0.03524652025859079, 32'sd0.016652837166573158, 32'sd-0.014742303273135327, 32'sd0.06355229432034147, 32'sd0.07068798347487132, 32'sd-0.047603723019748516, 32'sd0.11600947747509635, 32'sd0.007760176273397126, 32'sd-0.1718923529303087, 32'sd-0.2020360425374525, 32'sd-0.09412447521389165, 32'sd-0.04781431053806811, 32'sd-0.005794789747161439, 32'sd0.058504466170485124, 32'sd-0.03719658200634397, 32'sd0.08713878415049466, 32'sd0.058217763180616056, 32'sd0.01484704162967213, 32'sd-0.00990258074127896, 32'sd0.08191387197430257, 32'sd0.12565845431213563, 32'sd0.12651424876061168, 32'sd0.012979882221982198, 32'sd-0.05689729903523747, 32'sd0.024537529558292692, 32'sd0.04645142517791879, 32'sd0.08057429481313749, 32'sd-0.06420015139534398, 32'sd-0.06787712826045235, 32'sd0.043795867811126724, 32'sd0.00494934810800969, 32'sd5.036452226025631e-122, 32'sd0.04253422135228812, 32'sd-0.0352745341653891, 32'sd0.09469547136569137, 32'sd0.05531359677220245, 32'sd-0.0516026393160283, 32'sd-0.10683033673308731, 32'sd-0.13898839471454327, 32'sd0.04416137560459766, 32'sd-0.06259957937199054, 32'sd0.009114666758929746, 32'sd-0.03427691021697292, 32'sd0.042057425103109024, 32'sd0.12201295077992447, 32'sd0.05460994211263826, 32'sd-0.03467115911118169, 32'sd0.10534801243372655, 32'sd0.05711378860938303, 32'sd-0.015421403673003885, 32'sd-0.07591908661305687, 32'sd0.017345279927164548, 32'sd0.038339314365787316, 32'sd0.0378319011558997, 32'sd0.04463161014400577, 32'sd-0.07557460165187814, 32'sd0.06213110566431524, 32'sd0.09743374875303708, 32'sd-7.426625809076086e-123, 32'sd-7.155706624390175e-115, 32'sd-1.2164431860623495e-126, 32'sd-0.026760222666789145, 32'sd0.034306159264237406, 32'sd0.031723205164343474, 32'sd-0.04243621109075651, 32'sd-0.0830879603412248, 32'sd-0.23747259086305764, 32'sd-0.20209714384825087, 32'sd-0.11158524151344357, 32'sd0.03750157680135473, 32'sd0.03934685525726004, 32'sd0.026820397971794408, 32'sd-0.112623214700468, 32'sd-0.0365596451051559, 32'sd0.0073237620341468105, 32'sd0.12330182908953394, 32'sd-0.0492119679266187, 32'sd0.018162317442687044, 32'sd0.021543928062683217, 32'sd0.06948544280091569, 32'sd-0.01887553126085222, 32'sd-0.0028863193771580184, 32'sd-0.04411661526701764, 32'sd-0.020689673145182292, 32'sd0.03162451212223599, 32'sd0.03049064962044999, 32'sd-3.7779033001916634e-129, 32'sd2.550008736060644e-120, 32'sd2.900877038382324e-121, 32'sd-0.037453243560827514, 32'sd0.07266482421769806, 32'sd-0.035186773649098786, 32'sd-0.044028236210202014, 32'sd-0.13569596670058975, 32'sd-0.17651777921246714, 32'sd-0.1282062864716087, 32'sd-0.13156426322022086, 32'sd-0.05664993209648783, 32'sd-0.02654255863040355, 32'sd0.031375412237003034, 32'sd0.0072901532220722345, 32'sd-0.04614528436871834, 32'sd0.030347583203849737, 32'sd0.035249560380720156, 32'sd0.11547060544007455, 32'sd-0.01583753660565239, 32'sd-0.040884232300602195, 32'sd0.13918370979930111, 32'sd0.06742255743284405, 32'sd-0.0353276257104823, 32'sd-0.005454036068164161, 32'sd0.023074678842237416, 32'sd-0.01647842386819271, 32'sd0.01660727998265818, 32'sd-1.519625101825427e-116, 32'sd-3.3004116075824185e-123, 32'sd-7.906121326121648e-119, 32'sd-4.121555097472519e-122, 32'sd0.04914318795223621, 32'sd-0.012686454670199252, 32'sd-0.031043205070462328, 32'sd-0.059402001324252676, 32'sd0.061313073156287104, 32'sd0.002008660864169246, 32'sd-0.025013881184243036, 32'sd0.03601412097795019, 32'sd0.030754919038061188, 32'sd0.04232498640545779, 32'sd0.06635150481654345, 32'sd0.014262306984793933, 32'sd0.06977463257347101, 32'sd0.0369250687049142, 32'sd0.07236616865581648, 32'sd-0.0019627484155774946, 32'sd0.002206988615511408, 32'sd0.07049089433353722, 32'sd-0.06712563175257993, 32'sd-0.06625079862826358, 32'sd0.028894609061343078, 32'sd-0.034566963743195976, 32'sd0.04117120100783764, 32'sd-2.410303913708073e-125, 32'sd-1.636934939916947e-121, 32'sd5.334549917441324e-125, 32'sd-3.509821922508295e-125, 32'sd2.794537781190898e-115, 32'sd1.4087267932225283e-118, 32'sd0.028499241924351833, 32'sd0.06478571644445684, 32'sd-0.00025141964760625694, 32'sd0.0382625990839242, 32'sd-0.06844121070370954, 32'sd0.03684151847831829, 32'sd0.02643332590829202, 32'sd-0.04751769053057411, 32'sd-0.00041453276324217753, 32'sd0.04381690625868697, 32'sd-0.05354832921045313, 32'sd0.07063370728232192, 32'sd0.017551459703318045, 32'sd-0.031130381379203, 32'sd0.07214821267791693, 32'sd-0.008933289470408343, 32'sd-0.011797451672606141, 32'sd-0.009261353409161958, 32'sd0.0746587320590264, 32'sd0.02317136755279219, 32'sd-5.091536475522746e-125, 32'sd1.2349129925031592e-122, 32'sd-7.966287655637294e-120, 32'sd5.43075320991649e-123},
        '{32'sd-1.4362439448737e-123, 32'sd-5.979866110232433e-122, 32'sd5.774511921778884e-122, 32'sd-2.9465955559368767e-120, 32'sd1.442405365764318e-123, 32'sd-9.049471560730453e-125, 32'sd-8.766003915818958e-125, 32'sd7.337161783346994e-124, 32'sd3.309975906240234e-121, 32'sd5.40566046681218e-118, 32'sd5.7221224332483097e-126, 32'sd3.325012902866895e-122, 32'sd0.098788408615114, 32'sd0.08731293916238812, 32'sd0.09655661692337977, 32'sd0.11628270483725578, 32'sd-3.4847566390337536e-118, 32'sd3.371169909239952e-120, 32'sd3.3156413544134746e-122, 32'sd-2.103828682812613e-119, 32'sd-7.347893682387712e-116, 32'sd-2.0913724889528662e-124, 32'sd9.372427558894502e-125, 32'sd-3.4283170900677288e-124, 32'sd-1.5936495476911152e-125, 32'sd-9.844434258571911e-122, 32'sd1.585867599237723e-115, 32'sd-1.1993032366870867e-120, 32'sd3.601555494212801e-114, 32'sd3.3416726876798344e-121, 32'sd-6.25497198428939e-127, 32'sd5.282739558163197e-118, 32'sd0.03500534648746947, 32'sd0.10601957382990748, 32'sd0.062775549495331, 32'sd0.033073985376647186, 32'sd0.06890263681215118, 32'sd-0.030621292319249423, 32'sd0.13350303083598003, 32'sd0.138931124476061, 32'sd0.11782790745440412, 32'sd0.06537322862085398, 32'sd-0.0017444894132496959, 32'sd-0.04863195476732411, 32'sd0.003970897071768139, 32'sd-0.09024958438886878, 32'sd-0.04330627284755704, 32'sd-0.008614942899782764, 32'sd-0.053306241400541805, 32'sd-0.010526681876549298, 32'sd-0.0036160210682776037, 32'sd0.001761411766988788, 32'sd-3.16181394940844e-123, 32'sd2.4711734449947374e-120, 32'sd-1.819238976404624e-116, 32'sd1.882662739009015e-126, 32'sd-9.716925676198103e-121, 32'sd2.0571171688408924e-123, 32'sd-0.0019995067529523167, 32'sd-0.013098642237226992, 32'sd-0.025338841748598098, 32'sd0.06835826043003301, 32'sd0.07729635081113256, 32'sd0.12514264969095443, 32'sd0.059088882154994214, 32'sd0.05844675160772383, 32'sd-0.01487819209135659, 32'sd0.003236349981000761, 32'sd0.013214544611754604, 32'sd-0.016210572801650305, 32'sd-0.001374889641634123, 32'sd0.011662067920142061, 32'sd-0.03437431461554476, 32'sd-0.06160857891638832, 32'sd0.028728837421178086, 32'sd0.04700717717068374, 32'sd-0.018744657174342396, 32'sd0.09634519069632, 32'sd0.15594154479895062, 32'sd0.0465033021254365, 32'sd0.02660162461337601, 32'sd-0.0180867082907954, 32'sd-1.6834516772289277e-126, 32'sd-2.0805414543238858e-117, 32'sd2.699614042984016e-124, 32'sd6.632825822038807e-125, 32'sd-0.04059897876192609, 32'sd-0.018964109036822566, 32'sd0.03009738780376641, 32'sd0.06705018729134363, 32'sd0.06966670473493217, 32'sd0.006847298453805779, 32'sd0.08665269218407369, 32'sd0.002098968208050947, 32'sd-0.1027931684580069, 32'sd0.00032604664801596383, 32'sd-0.028967631768250852, 32'sd-0.08140166697783784, 32'sd-0.02735994646462963, 32'sd0.006227548007644621, 32'sd-0.08334646891007248, 32'sd0.0395465972960118, 32'sd0.04234560553272561, 32'sd0.01101355831550609, 32'sd0.0016820202159655918, 32'sd0.10478067771504952, 32'sd-0.029308712158843467, 32'sd0.13806098340100517, 32'sd-0.020026009590721372, 32'sd-0.0056977081307750125, 32'sd-0.13930957574771774, 32'sd-1.0161666435561545e-119, 32'sd1.7164158311462355e-126, 32'sd0.07226674628594405, 32'sd0.05465794803330392, 32'sd-0.02745000663200996, 32'sd-0.09159774961856403, 32'sd-0.11072388469171258, 32'sd0.07085626755189346, 32'sd0.006213309309057944, 32'sd-0.09834447741566793, 32'sd0.02539169688567019, 32'sd-0.024679893176803656, 32'sd-0.007327352584893396, 32'sd-0.002110198913508615, 32'sd0.12843751966948577, 32'sd0.07815782446159797, 32'sd0.06451385609930689, 32'sd-0.04077059053162514, 32'sd0.07451388249420697, 32'sd0.09308322652778106, 32'sd0.10281431707613761, 32'sd0.08818861134609646, 32'sd0.16862783348189433, 32'sd0.07399064499337435, 32'sd0.00982731921321211, 32'sd-0.08378028472064816, 32'sd-0.026112251051853642, 32'sd-0.08465354327413727, 32'sd0.07170229720591616, 32'sd-7.296225696153213e-125, 32'sd0.03794337217857394, 32'sd-0.03798442614787594, 32'sd0.06618841366136331, 32'sd-0.0160917323051601, 32'sd-0.01796682196269921, 32'sd0.025963660307252515, 32'sd-0.06778234696482004, 32'sd0.05870941014020211, 32'sd0.07343412946565293, 32'sd0.12013255240497613, 32'sd-0.015547416788159022, 32'sd-0.10913041488164066, 32'sd-0.14980565832697368, 32'sd-0.07612152877893454, 32'sd-0.08150529668293172, 32'sd-0.03442924897895039, 32'sd-0.0112589629084712, 32'sd-0.05896383026396862, 32'sd0.038519132522783564, 32'sd0.07666978075791003, 32'sd0.07362709840802446, 32'sd0.20302155214605533, 32'sd0.06512732252836095, 32'sd0.02425488545983943, 32'sd0.058580451988209076, 32'sd-0.14946840601436362, 32'sd0.019512717721179122, 32'sd2.2095963907728817e-119, 32'sd0.0007238035146764866, 32'sd-0.05661545105763424, 32'sd-0.00689575362378045, 32'sd-0.01428007704593311, 32'sd-0.053817556287071355, 32'sd-0.0446595688413834, 32'sd-0.024073122197004252, 32'sd0.036052711379769425, 32'sd0.06839653451670444, 32'sd0.0003356533572591839, 32'sd-0.04980745503151826, 32'sd-0.0971919407998709, 32'sd-0.012107758643496128, 32'sd-0.11208398821986865, 32'sd-0.06923141899664498, 32'sd-0.15249358991418513, 32'sd0.048191198379899235, 32'sd-0.021744178514922666, 32'sd-0.030446328228348894, 32'sd0.07515088562544638, 32'sd-0.02523813011890348, 32'sd0.0459266737452133, 32'sd0.03230007514175762, 32'sd0.14073573047723956, 32'sd-0.0438427638014818, 32'sd-0.028584889267248306, 32'sd-0.057316762481731856, 32'sd0.028666973245171687, 32'sd0.015374324735403688, 32'sd-0.023565857432208376, 32'sd-2.022220307912008e-07, 32'sd-0.005034341484967653, 32'sd-0.1378067390853748, 32'sd-0.13594584358852765, 32'sd-0.14572764698285873, 32'sd0.0387973405584054, 32'sd0.07728721952574892, 32'sd-0.08799446156548531, 32'sd-0.18376101363958908, 32'sd-0.17929648053562938, 32'sd-0.07302340247578325, 32'sd0.0544699026522904, 32'sd0.054591368968068446, 32'sd-0.04161087857564418, 32'sd0.030381752139112764, 32'sd-0.08354920966364464, 32'sd0.054027210774760984, 32'sd0.03206519897515158, 32'sd-0.01227943988470107, 32'sd0.00935512676549486, 32'sd0.04864676744381377, 32'sd0.019470624544431877, 32'sd0.02337600257284887, 32'sd0.043304506457621045, 32'sd-0.03366520687772756, 32'sd0.05773179943969408, 32'sd0.0026426813125645485, 32'sd-0.06257149055380822, 32'sd0.055784822707280385, 32'sd-0.07084422398114135, 32'sd-0.012484082060791078, 32'sd-0.043139602865176103, 32'sd-0.02317963803629651, 32'sd-0.05517562693510013, 32'sd-0.02430332260115033, 32'sd-0.06575025615885673, 32'sd0.010360621131300375, 32'sd-0.17800269279916753, 32'sd-0.039921149953516435, 32'sd0.15346914504371156, 32'sd-0.02514756724030429, 32'sd-0.13630098498568435, 32'sd-0.1060675738485061, 32'sd0.000847231366394505, 32'sd0.0006174860377950979, 32'sd-0.0012601855262283895, 32'sd0.02353939208946022, 32'sd0.03362674290832454, 32'sd0.11074825507302467, 32'sd0.03416409525045184, 32'sd-0.05405526363683692, 32'sd-0.014063174159573257, 32'sd-0.057903947284261716, 32'sd0.10767366545616167, 32'sd-0.037807336727070366, 32'sd0.017936421639628917, 32'sd0.10607175815723413, 32'sd-0.05568039718213289, 32'sd-0.017013525430951155, 32'sd0.03524544118095438, 32'sd0.0671488159157333, 32'sd-0.01259043057789639, 32'sd0.09243478472268249, 32'sd0.04779129911798601, 32'sd-0.00705324272999073, 32'sd-0.12715813193199446, 32'sd-0.0939880992776348, 32'sd-0.06269653119958879, 32'sd0.03841002407373042, 32'sd0.01967869330892254, 32'sd-0.05808188097972364, 32'sd-0.08288190688699992, 32'sd0.10890802262043212, 32'sd0.020060065741731872, 32'sd0.05805929040703057, 32'sd0.07930254765732915, 32'sd0.12986256997871287, 32'sd-0.04104202278216301, 32'sd0.018430193618364316, 32'sd-0.06077363220336098, 32'sd-0.056055727884913184, 32'sd-0.00647854145342395, 32'sd0.06205200734119324, 32'sd-0.025212493833419905, 32'sd-0.0632641506497732, 32'sd0.016941999601023227, 32'sd0.06407381807586236, 32'sd-0.04080524447104973, 32'sd0.14864718944199873, 32'sd0.10094414474995228, 32'sd0.11717638125901952, 32'sd0.06364342294387429, 32'sd0.06607272446777265, 32'sd-0.12884458214761976, 32'sd-0.026214978719240917, 32'sd-0.09294304041896854, 32'sd0.03116173860176135, 32'sd-0.10771236453855572, 32'sd-0.11110456299569424, 32'sd-0.0034740624752574545, 32'sd-0.08973463163669357, 32'sd-0.012807844583375829, 32'sd-0.07641865838665825, 32'sd-0.027321202448182032, 32'sd-0.02296817676610217, 32'sd0.024133026076285164, 32'sd-0.094539192415373, 32'sd-0.004899379178027973, 32'sd-0.016019534043366656, 32'sd0.06715798028073422, 32'sd0.010536581111489684, 32'sd-0.05768859017842773, 32'sd-0.018353459296938237, 32'sd0.03643490865329645, 32'sd0.08737550622646297, 32'sd0.07292207565784707, 32'sd0.07324431969834166, 32'sd0.15717032432532724, 32'sd0.19030369132307728, 32'sd0.15629891500914989, 32'sd0.08639264041941823, 32'sd0.05121951220906836, 32'sd-0.0854194836637106, 32'sd0.01000534287501546, 32'sd0.035050678329265963, 32'sd-0.11803547426855106, 32'sd-0.10549947231979467, 32'sd-0.07666205020008768, 32'sd-0.10623850339499405, 32'sd-0.03690442595627962, 32'sd0.04771818758971951, 32'sd-0.03210494400008879, 32'sd-0.049795745038238304, 32'sd-0.010289979044751879, 32'sd-0.0327072818078204, 32'sd0.1055137161305967, 32'sd0.029314760419863913, 32'sd0.041934239423838955, 32'sd0.03192220790404812, 32'sd0.019999529846296396, 32'sd0.08734408455842371, 32'sd0.0389580806290333, 32'sd0.07294841659640254, 32'sd-0.0677655031334135, 32'sd0.0991686111839047, 32'sd0.07725016832430308, 32'sd0.1596216040627011, 32'sd0.16424739849516581, 32'sd0.07378833133583154, 32'sd0.07902575294089065, 32'sd-0.12990616834450647, 32'sd-0.01037553055610446, 32'sd0.010123624685189936, 32'sd0.02780808223262088, 32'sd-0.04035908958225758, 32'sd-0.15586139990039177, 32'sd-0.016498739365280086, 32'sd0.012243032873466638, 32'sd-0.028690064255327597, 32'sd-0.13635014664462405, 32'sd-0.06671429317567805, 32'sd0.06113518493955635, 32'sd-0.01432676049902306, 32'sd-0.012622406024743066, 32'sd0.07982336910539352, 32'sd0.05929491828108797, 32'sd0.01567631406926902, 32'sd0.04186270312879244, 32'sd0.07066956875298236, 32'sd0.028798946283724626, 32'sd0.04874434478587629, 32'sd-0.06590639756608374, 32'sd0.029245027211837082, 32'sd0.10167104055122542, 32'sd0.12954237036223887, 32'sd0.05336656393223988, 32'sd0.00010774253235618421, 32'sd0.04670801102658889, 32'sd-0.12229008779384969, 32'sd0.03289357736926065, 32'sd0.11958161920013115, 32'sd-0.06673497344326287, 32'sd-0.06918490222764062, 32'sd0.04752285136600431, 32'sd-0.11604531681862615, 32'sd-0.020878402835935363, 32'sd-0.13798303174572873, 32'sd-0.005172532682783595, 32'sd0.0480216404477468, 32'sd-0.12993467650693147, 32'sd0.0784730988819294, 32'sd0.04909286637321878, 32'sd-0.04863004896263039, 32'sd-0.03290207342121938, 32'sd0.10455841784274963, 32'sd-0.047541967464799696, 32'sd-0.018585716114169152, 32'sd-0.07695799079452491, 32'sd0.05361188953966723, 32'sd0.003900144525059329, 32'sd0.051728374166669984, 32'sd-0.025956290242765474, 32'sd0.05688522027214881, 32'sd0.000503571495823858, 32'sd0.14414990112769466, 32'sd0.005305613214135698, 32'sd-0.023224647283447346, 32'sd0.035563565255898676, 32'sd-0.11069976403011755, 32'sd-0.0465105893548577, 32'sd-0.09900375569035394, 32'sd-0.03866119495693474, 32'sd-0.1055141759359519, 32'sd-0.02899714181143552, 32'sd0.011707378949642886, 32'sd-0.028473330553368356, 32'sd-0.057174551538031505, 32'sd-0.047571359063170136, 32'sd-0.022977164741329343, 32'sd0.06273680781390187, 32'sd-0.06225467144524899, 32'sd0.037725037276514696, 32'sd0.023604334566505514, 32'sd0.05549400532709097, 32'sd-0.14483884502324518, 32'sd-0.00692384078985663, 32'sd0.009452188616010325, 32'sd0.0810408861095822, 32'sd0.11886425190321481, 32'sd0.07124383309746733, 32'sd0.010043530361110041, 32'sd-0.00496868491202296, 32'sd0.10113819424052393, 32'sd0.06423825154076131, 32'sd-0.04419867512638217, 32'sd0.057244674549441675, 32'sd-0.09924177809409199, 32'sd-0.03783441638922592, 32'sd-0.14374274148098948, 32'sd-0.03462215459010329, 32'sd0.001663961209808616, 32'sd0.008092081014561115, 32'sd-0.0755199496744658, 32'sd-0.09959156844607586, 32'sd-0.09091897454831026, 32'sd-0.02609114390675058, 32'sd0.006230466352152729, 32'sd-0.06650260762193584, 32'sd-0.02209838304113627, 32'sd0.010636000048865259, 32'sd0.006503410929823337, 32'sd0.0015313630915073646, 32'sd-0.09041966322375537, 32'sd-0.0814086694496851, 32'sd-0.060664471904371756, 32'sd-0.04675393505493699, 32'sd-0.01661726926599455, 32'sd0.07964485090362906, 32'sd0.07944297393834514, 32'sd0.025933780982070172, 32'sd0.0935025958963231, 32'sd-0.027941434915011106, 32'sd-0.04796181314171475, 32'sd0.01744028300547159, 32'sd0.0002610783833770491, 32'sd0.033507271967100474, 32'sd0.0767026912854498, 32'sd-0.026200109564317915, 32'sd0.03706654259866093, 32'sd0.01317036002595105, 32'sd0.012996157932754543, 32'sd-0.003928300404519906, 32'sd0.052637786403983304, 32'sd0.057065449027285955, 32'sd0.06583140915065623, 32'sd-0.026563610784692812, 32'sd-0.00857373039312142, 32'sd1.8742288989830503e-117, 32'sd0.054472703355460714, 32'sd-0.08253847551550975, 32'sd0.014614129689805638, 32'sd-0.03904477508550668, 32'sd-0.10964343150706277, 32'sd0.07085234332215064, 32'sd0.05561061343168282, 32'sd0.07952134343964563, 32'sd-0.0654377369214182, 32'sd0.03550604756926376, 32'sd-0.04713663173972852, 32'sd-0.002412450461314253, 32'sd0.0032090753495909994, 32'sd0.08023680509826447, 32'sd-0.010186348693553652, 32'sd0.04207419674035823, 32'sd0.06999789184639564, 32'sd0.09000831092762998, 32'sd-0.004059494676714518, 32'sd0.08115288081356123, 32'sd-0.02073567264317342, 32'sd-0.016029241886805295, 32'sd-0.05345371140482924, 32'sd-0.019351468270220797, 32'sd-0.0317065777098944, 32'sd-0.05094582517706829, 32'sd0.10402935811720129, 32'sd-0.022680834908173103, 32'sd-0.030597277267975807, 32'sd-0.0059296025477270625, 32'sd-0.08229577204611692, 32'sd-0.025270147633295388, 32'sd-0.054971125171383, 32'sd-0.01774989469592704, 32'sd0.13776418222020298, 32'sd0.09772385085201477, 32'sd0.10269143699865137, 32'sd0.05136456490593744, 32'sd-0.1131574823315669, 32'sd0.08257521283882865, 32'sd0.010981680696308527, 32'sd0.12580103676884716, 32'sd0.1897799335216766, 32'sd0.03575519224754963, 32'sd-0.06711335958726654, 32'sd0.04119617270854536, 32'sd0.07598750931519883, 32'sd-0.004255248297848773, 32'sd-0.08352589511806607, 32'sd0.015524526458888098, 32'sd-0.03937521084139359, 32'sd-0.01888873893280604, 32'sd0.039736898914202574, 32'sd0.019317283534500903, 32'sd-0.023176440515255595, 32'sd-0.0038813292147202192, 32'sd0.014614783394939074, 32'sd-0.06023597391562143, 32'sd0.03975407659301143, 32'sd-0.10844989989620639, 32'sd-0.12944248711622555, 32'sd0.03588062587667785, 32'sd0.03169399805911659, 32'sd0.061113027789021716, 32'sd0.026080939389066957, 32'sd0.05012047581868761, 32'sd-0.07943974770776004, 32'sd-0.02213960302283391, 32'sd0.16467230451957457, 32'sd0.07660356325393934, 32'sd0.08051040746319438, 32'sd0.003397669362029805, 32'sd-0.001166890918167123, 32'sd-0.07112662838012582, 32'sd-0.05979917689922078, 32'sd-0.010318117972485963, 32'sd0.025764365864896253, 32'sd0.055459583681630266, 32'sd0.017872044233383563, 32'sd-0.07152486829786911, 32'sd-0.02206556851589967, 32'sd0.009508235112262547, 32'sd-0.027154170711943586, 32'sd2.2392463126579515e-125, 32'sd0.006229762928361548, 32'sd-0.08183567696621348, 32'sd-0.023543696303741694, 32'sd-0.09499273544373399, 32'sd-0.09518307485113205, 32'sd-0.04991515958566266, 32'sd-0.007235584632118268, 32'sd-0.028071216232955835, 32'sd0.0016732985311511104, 32'sd-0.07605521066521875, 32'sd-0.0516844637076738, 32'sd0.07054013648343073, 32'sd-0.005499093953905222, 32'sd0.10675605684986537, 32'sd0.12232692273599911, 32'sd-0.06777422269979858, 32'sd-0.041854628614944295, 32'sd-0.03870016355417009, 32'sd-0.024079493699529237, 32'sd-0.033666863257833454, 32'sd0.04749041654688628, 32'sd0.0645888351569114, 32'sd-0.07381376433447509, 32'sd0.011831230179387137, 32'sd0.011530197427873059, 32'sd0.1348876704918782, 32'sd0.14562496875567266, 32'sd-0.030896654358201353, 32'sd-0.03490859600255308, 32'sd0.03750357906401603, 32'sd-0.08445521015066856, 32'sd-0.04549238904571466, 32'sd-0.11833273430868982, 32'sd-0.03247198411288936, 32'sd-0.074861320803268, 32'sd-0.046606488057303504, 32'sd-0.027032917012121904, 32'sd-0.049114852218189786, 32'sd0.035499548949720044, 32'sd0.1038264098522709, 32'sd0.07626328546723327, 32'sd0.025240469511327253, 32'sd0.02556726268245864, 32'sd0.06050449488991754, 32'sd0.06246395606365116, 32'sd-0.07478847156547942, 32'sd0.01609294990621234, 32'sd0.0924511928605613, 32'sd0.06114397903642946, 32'sd-0.03250474731723245, 32'sd0.06456400269107637, 32'sd-0.08961833631980438, 32'sd0.06515711957080358, 32'sd-0.012197623117658684, 32'sd-0.018769561096120845, 32'sd0.03416236206241035, 32'sd0.00036457752300917995, 32'sd-0.06997978888540793, 32'sd-0.06006793368497329, 32'sd-0.03826701484160145, 32'sd-0.0701187173129962, 32'sd-0.007261106395013602, 32'sd-0.11244048008745851, 32'sd-0.07079627322984045, 32'sd-0.08103851134609022, 32'sd-0.07282325278509943, 32'sd-0.026703233523994306, 32'sd0.10093646169796897, 32'sd0.16950218954881835, 32'sd0.0038627657469950654, 32'sd0.11756354692528187, 32'sd0.15487734558020816, 32'sd0.10296986792583211, 32'sd0.10833709474940785, 32'sd0.12702436511553075, 32'sd0.005361989044296274, 32'sd0.07178562186454533, 32'sd0.028771015855549795, 32'sd-0.12492142392454587, 32'sd-0.13001398092829047, 32'sd-0.10521491266421208, 32'sd0.0795562213989709, 32'sd0.007138412089637623, 32'sd2.0509139411994528e-116, 32'sd-0.01733653058108829, 32'sd-0.05150579149298103, 32'sd0.022871032612430568, 32'sd0.05441625910158467, 32'sd0.012479372714087897, 32'sd0.00830854997097071, 32'sd0.05558611036785788, 32'sd-0.019597712434196796, 32'sd-0.1082305304349962, 32'sd0.014735832059712765, 32'sd-0.04860270110493148, 32'sd0.04147590084986642, 32'sd-0.03204797863908445, 32'sd0.10655634099418232, 32'sd-0.07528427179866523, 32'sd0.03893897418871488, 32'sd0.061239836900128124, 32'sd0.13292240985862658, 32'sd0.0791101373402588, 32'sd-0.022428489260218953, 32'sd0.006756128301953761, 32'sd-0.06681083070977431, 32'sd-0.06863457446895656, 32'sd-0.002353218097968066, 32'sd0.04063414568016676, 32'sd-0.061254182623300346, 32'sd1.1807036635351341e-122, 32'sd-4.705001502320802e-128, 32'sd-7.403401466455116e-115, 32'sd-0.034531943719710134, 32'sd-0.024676860151997815, 32'sd0.08240383177265422, 32'sd0.045813090849252745, 32'sd0.03436518727147148, 32'sd0.039857013768643826, 32'sd0.05773520399133882, 32'sd0.014168180653234398, 32'sd-0.011139103113540487, 32'sd-0.12393062590359545, 32'sd-0.14850851095541143, 32'sd-0.15286901878527068, 32'sd-0.059735894054721024, 32'sd-0.007661000845830679, 32'sd0.02641712903434719, 32'sd0.026263538879188225, 32'sd-0.004658206885214278, 32'sd0.0020656270273653396, 32'sd-0.07385943136850834, 32'sd-0.10157460832882895, 32'sd-0.11508052957639012, 32'sd-0.08154080397642222, 32'sd-0.018415374344124432, 32'sd0.03851667179963029, 32'sd-0.021314858054846845, 32'sd-8.218968721381019e-119, 32'sd2.6893983399871524e-124, 32'sd-1.2891596022408039e-114, 32'sd0.07414381906156614, 32'sd0.03417727052677119, 32'sd-0.0419986687337303, 32'sd-0.04825510669026919, 32'sd0.04270151439719492, 32'sd0.03641398786815383, 32'sd-0.09021886679674382, 32'sd-0.018885605962096486, 32'sd-0.08081293710583837, 32'sd-0.07721029830742653, 32'sd-0.12166491448172714, 32'sd-0.1055475413501157, 32'sd-0.046172397612013236, 32'sd-0.0365213436790288, 32'sd-0.033942497873447525, 32'sd0.08709827214728891, 32'sd0.08317108917417179, 32'sd-0.0897468545523859, 32'sd-0.06118657062932832, 32'sd-0.05770120226669377, 32'sd-0.02114959885860928, 32'sd-0.005347170590268288, 32'sd0.00567515872451677, 32'sd0.03966652269681222, 32'sd0.0348725428864473, 32'sd2.0179143883519875e-117, 32'sd1.2210183542979712e-118, 32'sd-9.344366368399406e-126, 32'sd-9.63431451110366e-121, 32'sd-0.019198037368235714, 32'sd0.014916936718464571, 32'sd-0.04422677973986827, 32'sd0.006270945003006459, 32'sd-0.08834832620124727, 32'sd-0.14690742655479766, 32'sd-0.06905766423802286, 32'sd-0.02795888465473741, 32'sd0.0948987276292197, 32'sd0.03822595015483175, 32'sd0.103385215743889, 32'sd0.03577367824827839, 32'sd0.05008282628941957, 32'sd-0.1095837949627735, 32'sd-0.024356753655787145, 32'sd-0.08331401679034582, 32'sd-0.10442904255592729, 32'sd-0.09279444071983665, 32'sd-0.04387630697048158, 32'sd0.042071725144832664, 32'sd0.04714177601959415, 32'sd-0.012819209273255321, 32'sd0.027783260971224532, 32'sd-6.700529372433096e-120, 32'sd1.1049633205883313e-122, 32'sd-5.660584072784467e-128, 32'sd3.7602778812127334e-119, 32'sd-6.203920663395737e-124, 32'sd-7.315216177633078e-118, 32'sd0.045507716757534795, 32'sd-0.03234871427702333, 32'sd0.018245767187086245, 32'sd0.02102884725133883, 32'sd-0.042733903897606146, 32'sd0.018874725235081873, 32'sd0.01740431174815096, 32'sd-0.0008872996535088841, 32'sd-0.023792372051676405, 32'sd-0.00854865449440204, 32'sd0.032154951769878246, 32'sd0.03400252697791557, 32'sd0.0266827723281266, 32'sd-0.026691643939311862, 32'sd0.05234977304126184, 32'sd-0.02379506145177125, 32'sd-0.023785585140979917, 32'sd0.11319233197958255, 32'sd0.03627178293680116, 32'sd0.052317854409113636, 32'sd-1.8063422591917789e-127, 32'sd-2.2414543225225054e-122, 32'sd4.624514906332157e-118, 32'sd3.331642126967644e-124},
        '{32'sd1.2876094990985924e-125, 32'sd-3.188566101654033e-116, 32'sd9.852227415056136e-119, 32'sd-8.34997907526865e-117, 32'sd-1.3904042335226426e-125, 32'sd-7.681330438465663e-124, 32'sd-5.22852475833364e-124, 32'sd2.837965663627899e-126, 32'sd2.1658876760387967e-118, 32'sd2.7133778620021413e-124, 32'sd-5.381515087348417e-126, 32'sd1.3083754942099625e-124, 32'sd0.05309714422943896, 32'sd-0.05531019064166472, 32'sd-0.026980271121253032, 32'sd0.013195018343868225, 32'sd4.881183911023187e-118, 32'sd-1.6716163666763962e-123, 32'sd2.035271730468814e-127, 32'sd-2.2757192853953215e-119, 32'sd6.244288168306144e-126, 32'sd-1.287788329195353e-118, 32'sd2.3390092401670617e-124, 32'sd3.060219095825229e-122, 32'sd-9.841729916485285e-124, 32'sd-1.3803926444630006e-123, 32'sd-2.000512602646986e-124, 32'sd-8.548912242100531e-123, 32'sd9.765414893976291e-123, 32'sd1.549629939737286e-123, 32'sd-3.76600864736435e-119, 32'sd1.1618840826535508e-115, 32'sd0.0945564950306643, 32'sd-0.04560018748030133, 32'sd-0.038885245181670705, 32'sd-0.0012520967294090486, 32'sd0.0017208073949934145, 32'sd-0.05887670741765971, 32'sd0.03940114739776879, 32'sd0.03743887638798031, 32'sd0.1253229820326349, 32'sd-0.03175700031816393, 32'sd0.05979386189366935, 32'sd-0.13328004665015852, 32'sd-0.023728028326181094, 32'sd-0.004301157993395136, 32'sd0.005574895623916399, 32'sd-0.017065506488648154, 32'sd0.07900784635018329, 32'sd0.035155326206232844, 32'sd-0.019164323290415106, 32'sd-0.021417452190076038, 32'sd8.530844481046986e-117, 32'sd-6.256547141717728e-117, 32'sd3.3426993418928963e-118, 32'sd-1.1957293363275187e-126, 32'sd-2.0948740915311843e-117, 32'sd-3.2406313455345993e-116, 32'sd-0.01839420588402075, 32'sd-0.01990234060761615, 32'sd-0.008984985604372211, 32'sd-0.03096906885094392, 32'sd0.014515609353205717, 32'sd-0.002514384292702829, 32'sd-0.10599010979678501, 32'sd-0.1343614568552941, 32'sd-0.004149612380527326, 32'sd0.08301352523603445, 32'sd-0.019305739475978027, 32'sd-0.025308529587312372, 32'sd-0.014286695200963958, 32'sd-0.040707219532329926, 32'sd0.03685436962124313, 32'sd0.050361660138943956, 32'sd0.08061999029255267, 32'sd0.0093394268652438, 32'sd0.06571764974785516, 32'sd0.10402131706890197, 32'sd0.1061786940239496, 32'sd0.04844064358998567, 32'sd-0.05019018466723032, 32'sd0.007070923163808264, 32'sd-1.0185295253706684e-119, 32'sd8.438262209858026e-115, 32'sd1.3539446422661507e-125, 32'sd-7.356858599205174e-124, 32'sd-0.004460512965010198, 32'sd-0.03602992666648018, 32'sd-0.09818133836289207, 32'sd-0.013519018413519362, 32'sd0.010927448893176376, 32'sd-0.10302382115170987, 32'sd-0.11714191452238905, 32'sd-0.012288145234112018, 32'sd-0.026205504383988953, 32'sd-0.001960466046616366, 32'sd-0.18243318661413818, 32'sd-0.16131170471836256, 32'sd0.006400769677523201, 32'sd-0.09446457421204502, 32'sd-0.16213588332454862, 32'sd0.09609124503001229, 32'sd-0.02858638570928344, 32'sd-0.021600967004372328, 32'sd-0.09876612366607271, 32'sd-0.06821641214358928, 32'sd0.07314451897767861, 32'sd-0.07645283232559795, 32'sd0.03074059557089735, 32'sd0.03614701333470749, 32'sd-0.005243504018209946, 32'sd3.121434347461754e-116, 32'sd7.628652292121937e-116, 32'sd-0.017038688299532822, 32'sd-0.03313875838442063, 32'sd0.07266053903321651, 32'sd-0.09825839726070598, 32'sd-0.07930205620247377, 32'sd-0.058572458072833386, 32'sd-0.07323809649387264, 32'sd-0.10478801883227157, 32'sd0.017141455937784017, 32'sd0.02335085022420571, 32'sd-0.05506324374275234, 32'sd-0.05410725580383092, 32'sd-0.01162519320458115, 32'sd-0.059714879503972924, 32'sd-0.06676485351998764, 32'sd-0.05038077464306684, 32'sd0.021951474220801997, 32'sd0.11628421663770257, 32'sd0.05412178319172684, 32'sd0.031074292507988682, 32'sd0.023593120026896373, 32'sd-0.017143412227778876, 32'sd-0.05829251533152614, 32'sd0.00031360378323852815, 32'sd0.047148372846712854, 32'sd0.005094757020937303, 32'sd0.028626106242540167, 32'sd9.583467024478346e-118, 32'sd0.03354111533412688, 32'sd-0.017465908202508956, 32'sd0.04080558274133458, 32'sd-0.026671450700555006, 32'sd-0.06623156286009374, 32'sd-0.21764246951727095, 32'sd-0.10775321576860349, 32'sd-0.049975184547336786, 32'sd0.05871108741587826, 32'sd0.13339124050936693, 32'sd-0.006357423755433182, 32'sd-0.03061486578259231, 32'sd0.008414520236724479, 32'sd-0.05294218675307735, 32'sd-0.11494643601559712, 32'sd-0.05962476820365565, 32'sd0.10543281582236455, 32'sd0.046396716082751664, 32'sd0.004390031844667288, 32'sd0.051046548108824925, 32'sd0.07304521413584218, 32'sd-0.11481658617265243, 32'sd-0.1136295415370557, 32'sd-0.0911400785041899, 32'sd0.004612923415352185, 32'sd0.04334397246240577, 32'sd-0.05976100967830674, 32'sd-2.1846958084217318e-116, 32'sd-0.014488666662223315, 32'sd-0.02794176191455135, 32'sd-0.03444952258441978, 32'sd0.08859586120493768, 32'sd0.03204366976596691, 32'sd-0.29669096822597796, 32'sd-0.11193632716976011, 32'sd-0.04933849596791701, 32'sd0.10603941557552078, 32'sd0.0032914410533993565, 32'sd0.010062411942262466, 32'sd0.04453502374835769, 32'sd-0.00984971346192895, 32'sd-0.05943704261824067, 32'sd-0.11363254196556212, 32'sd-0.014773967851617152, 32'sd0.0015914446040407521, 32'sd0.01721451812692937, 32'sd0.025371245211957383, 32'sd0.11628510176529468, 32'sd-0.04869185582127208, 32'sd0.021645056033488954, 32'sd-0.06308181197850472, 32'sd-0.08755767761431152, 32'sd-0.03331478637105753, 32'sd-0.08806130789324855, 32'sd0.0889121436515139, 32'sd-0.04957982561326041, 32'sd-0.03027360348276914, 32'sd-0.13261319830791618, 32'sd-0.07155483646485479, 32'sd-0.09535974788299506, 32'sd-0.18494641817057228, 32'sd-0.22693987519777506, 32'sd-0.1426996495325985, 32'sd0.08433921086718454, 32'sd0.05712665260823823, 32'sd0.0901680187793636, 32'sd0.1124268368396922, 32'sd0.03232237128019466, 32'sd-0.04626315618103587, 32'sd-0.018322508227788397, 32'sd0.07408374678657581, 32'sd0.09190318655187485, 32'sd0.08953859832368292, 32'sd0.07329173352836924, 32'sd-0.00878340790415694, 32'sd0.07527059206393329, 32'sd-0.050772171003181966, 32'sd-0.07216257222276118, 32'sd-0.08393403914118104, 32'sd0.04237348845208087, 32'sd-0.08337374123112266, 32'sd0.03269315442042416, 32'sd-0.06396268076548253, 32'sd-0.009053884858995711, 32'sd-0.011204109869672605, 32'sd0.029770181295581708, 32'sd0.02813666994935278, 32'sd-0.044592777802069314, 32'sd-0.2165701260942703, 32'sd-0.27440177368904844, 32'sd-0.11062748399849061, 32'sd0.06125762008166191, 32'sd0.03440020181012648, 32'sd-0.0672452093709319, 32'sd0.15234434833045196, 32'sd-0.01970893100435648, 32'sd0.009796391252362563, 32'sd-0.04968777542924785, 32'sd-0.05107619669610668, 32'sd0.03053332062575938, 32'sd0.042967121054636404, 32'sd-0.027035384148377375, 32'sd-0.22189759969882744, 32'sd-0.1222574186899597, 32'sd-0.15034505591563546, 32'sd-0.1388231994461838, 32'sd-0.08467667381672206, 32'sd0.08539812972205067, 32'sd-0.1366358059387604, 32'sd-0.028028520071195474, 32'sd0.0044516827898631916, 32'sd-0.035567407510180435, 32'sd-0.0949117550540238, 32'sd0.02877325583663374, 32'sd-0.0076666446916864904, 32'sd-0.06913481390865373, 32'sd-0.21336580011531997, 32'sd-0.18228968511119217, 32'sd-0.032695611334075524, 32'sd0.00998172592175217, 32'sd-0.017745786419171475, 32'sd-0.03381454660776707, 32'sd0.11424580874899204, 32'sd0.02815864391361378, 32'sd0.009236811927831049, 32'sd-0.17660352999921228, 32'sd-0.07475158259782043, 32'sd0.11795838080406851, 32'sd-0.11570581455950515, 32'sd-0.2230063763850402, 32'sd-0.19201709148100787, 32'sd-0.1170320339302877, 32'sd-0.1088465585781874, 32'sd-0.1578214242241179, 32'sd-0.055892595742480386, 32'sd-0.05799705764726956, 32'sd0.038046085824146154, 32'sd0.04398742404404094, 32'sd0.0193696101576564, 32'sd-0.06411802364141907, 32'sd0.00860113451136867, 32'sd-0.06472435787459721, 32'sd-0.03855800421118972, 32'sd-0.05600064208970772, 32'sd-0.14096925037157465, 32'sd-0.33318757307910113, 32'sd-0.10807083003478596, 32'sd0.04440965382833778, 32'sd0.10804039458268538, 32'sd-0.018571435152066974, 32'sd0.08873507080741495, 32'sd0.027589599411001104, 32'sd-0.028324009187979005, 32'sd-0.1991473617022306, 32'sd0.045990160965447696, 32'sd-0.05567860957879294, 32'sd-0.15290590297867404, 32'sd-0.1423880062309681, 32'sd-0.20272454028887316, 32'sd-0.04808754695478446, 32'sd-0.06584246442077647, 32'sd-0.07053298546581264, 32'sd-0.06030880969057543, 32'sd0.059054487593658646, 32'sd-0.017771610777282155, 32'sd0.058203000584538096, 32'sd-0.06999514935980063, 32'sd-0.04252067698408261, 32'sd-0.028527468181300815, 32'sd0.007406462257464999, 32'sd-0.06789161020525639, 32'sd-0.07669218057366696, 32'sd-0.05856894961968876, 32'sd-0.18063519979040815, 32'sd-0.09199797284659539, 32'sd0.08730158683567252, 32'sd0.13303926195891197, 32'sd0.04640601730066236, 32'sd0.028862636668659982, 32'sd0.12629294328679458, 32'sd0.01946019708700172, 32'sd-0.16040515193718688, 32'sd-0.14889022202207217, 32'sd0.06902220198929265, 32'sd0.022624534832706517, 32'sd0.008291639144375371, 32'sd0.04194691953191932, 32'sd-0.06288373373135242, 32'sd-0.04954181923917989, 32'sd-0.11494854020286188, 32'sd0.034250521993404705, 32'sd-0.045999159785378364, 32'sd-0.07539924529782872, 32'sd0.055831619426939594, 32'sd-0.1079877678298261, 32'sd-0.037670229395701096, 32'sd0.020149429833208343, 32'sd-0.09046544000141761, 32'sd-0.005776356590911327, 32'sd-0.021992771960520734, 32'sd-0.08497960393291651, 32'sd-0.14539595283307843, 32'sd-0.036045620047528135, 32'sd-0.035602597309894034, 32'sd-0.0016263992743025283, 32'sd0.08691006775905273, 32'sd0.17378769783247808, 32'sd0.20988721478624048, 32'sd-0.07065363209020878, 32'sd-0.14809713942734595, 32'sd-0.0074131569454243896, 32'sd-0.1521437784103121, 32'sd-0.01566341364356247, 32'sd-0.05502474803400727, 32'sd-0.10173322002487264, 32'sd-0.015482644427055785, 32'sd-0.002572635722748099, 32'sd0.019902940640012023, 32'sd-0.025489494371785215, 32'sd-0.022682486028193748, 32'sd-0.00015850571932589128, 32'sd0.024649693850405923, 32'sd-0.04137071565585678, 32'sd-0.044550636646625126, 32'sd0.0007820906261153565, 32'sd-0.014611713260058733, 32'sd-0.06637877420845625, 32'sd0.08065256254632129, 32'sd-0.05139566309864585, 32'sd-0.18864009837876522, 32'sd-0.08745453294599875, 32'sd-0.08912078408185603, 32'sd-0.04344901204361207, 32'sd0.11106091782229756, 32'sd0.012915456340434561, 32'sd0.10469337181994068, 32'sd-0.05779339462446262, 32'sd-0.16519240049862005, 32'sd-0.11384767116951408, 32'sd-0.14544255465343986, 32'sd-0.07715114089554465, 32'sd-0.07051714703314634, 32'sd0.002609376259101867, 32'sd0.0704776460830279, 32'sd0.04362973849750262, 32'sd0.022283127918450146, 32'sd-0.16436368510905397, 32'sd-0.131334801271916, 32'sd-0.24620449201926736, 32'sd-0.06145905320652373, 32'sd-0.046509773951283445, 32'sd0.04404896121843103, 32'sd-0.02643489261306782, 32'sd0.012085450283803279, 32'sd-0.07986902424585339, 32'sd0.00040117508510562354, 32'sd0.029509916822391763, 32'sd-0.14154356609296936, 32'sd-0.07487865303192812, 32'sd-0.07861105340878909, 32'sd0.05364132926590592, 32'sd0.07356225071222654, 32'sd-0.010981206754185074, 32'sd0.08557018431102759, 32'sd0.05606736483568154, 32'sd-0.038622492033946194, 32'sd-0.11545860303770694, 32'sd-0.02631561320698032, 32'sd-0.07093419876265546, 32'sd0.0008964602840854728, 32'sd0.005897476225682711, 32'sd0.061652684677829125, 32'sd0.04144276460766692, 32'sd-0.03953444000425607, 32'sd-0.05749043557435539, 32'sd0.01952006929191441, 32'sd-0.1291970651223378, 32'sd-0.03837656945780732, 32'sd0.010341443582210022, 32'sd0.04182862545953308, 32'sd0.0031807781733751484, 32'sd-0.12935110719003406, 32'sd-0.053367575388594046, 32'sd-0.027473845183245988, 32'sd0.03853732625521212, 32'sd-0.14482162710341567, 32'sd-0.0844535014422664, 32'sd-0.10373848327629386, 32'sd0.08615091831873282, 32'sd0.08552074664304486, 32'sd0.15248329671221528, 32'sd0.06452768563710273, 32'sd-0.051780995095789484, 32'sd-0.11449369512952656, 32'sd-0.06661108346467047, 32'sd-0.12973469113008718, 32'sd-0.04009363288479974, 32'sd-0.017997561343734446, 32'sd-0.02888113470373696, 32'sd0.05703346515024395, 32'sd0.05662706353037414, 32'sd-0.10196726554015018, 32'sd0.0060380482331493296, 32'sd-0.0899635136157131, 32'sd-0.11127811066055367, 32'sd-0.0891038576852381, 32'sd0.01697645248381286, 32'sd0.04306101855457712, 32'sd-0.011749646393799803, 32'sd-0.08522135532068373, 32'sd0.042092220517999025, 32'sd-0.028814056726974506, 32'sd0.08423063091574087, 32'sd-0.04354733761025428, 32'sd-0.03138598388323831, 32'sd-0.009455557097603666, 32'sd0.030580041453239747, 32'sd0.08140125542992635, 32'sd0.11878616724177514, 32'sd-0.02605166493575558, 32'sd0.007161967016589435, 32'sd-0.07709872695620835, 32'sd-0.11861726587568618, 32'sd-0.11103544294410948, 32'sd-0.03823236842997731, 32'sd0.1410073504149063, 32'sd0.06487045907960232, 32'sd0.03247593034898524, 32'sd0.12779183652668952, 32'sd-0.11911401662552643, 32'sd0.007064067023766975, 32'sd-0.06816006540469648, 32'sd-0.10297913603211972, 32'sd-0.11878443774295092, 32'sd-0.07504175723969578, 32'sd1.4939883821742185e-123, 32'sd-0.052701332737006265, 32'sd0.041557281079732965, 32'sd-0.12768911875535152, 32'sd0.03158652772676735, 32'sd0.04010075692021235, 32'sd0.06404500859757051, 32'sd0.06641651586006368, 32'sd0.06403534133968247, 32'sd-0.04304986910032688, 32'sd0.06332138774892265, 32'sd0.08986683301845659, 32'sd0.03338775343830571, 32'sd-0.0066571805842194865, 32'sd0.0027009702002141756, 32'sd-0.1441886141182463, 32'sd-0.003686635355573306, 32'sd0.1667487305412836, 32'sd0.14658968387774723, 32'sd0.07551328402731511, 32'sd0.10010537830907434, 32'sd0.09396473343598134, 32'sd-0.03405851506267349, 32'sd-0.1374135202275056, 32'sd-0.03254113681153985, 32'sd-0.1012807951060287, 32'sd-0.03669513386591401, 32'sd-0.07569624250090483, 32'sd-0.006212515234144969, 32'sd-0.01812736401144965, 32'sd-0.03962878419694948, 32'sd0.015770620306634446, 32'sd0.03699514280485536, 32'sd0.08046906320308149, 32'sd0.04441191754881619, 32'sd0.025488007605489773, 32'sd0.12245133514939802, 32'sd-0.007422194442917415, 32'sd0.016002774007314986, 32'sd0.010905624041831975, 32'sd-0.04246047125820337, 32'sd4.232268547239858e-05, 32'sd0.009513297843897463, 32'sd0.10200137413609787, 32'sd0.010111373753757539, 32'sd0.12202951457703548, 32'sd0.0505469607928114, 32'sd0.0569252012641281, 32'sd0.07173703377812533, 32'sd-0.0301937378512044, 32'sd-0.12884509578506695, 32'sd-0.16942339987604457, 32'sd-0.0808465589747231, 32'sd-0.14222448971524168, 32'sd0.06977094263729998, 32'sd-0.022750431570680196, 32'sd-0.00019034185012856584, 32'sd-0.033322008078477565, 32'sd0.06069950621601711, 32'sd0.0940417502046999, 32'sd0.014780809756441584, 32'sd0.021880445417044175, 32'sd0.13210015359222319, 32'sd0.06795554541944814, 32'sd0.09499814152997253, 32'sd0.003652721892865639, 32'sd-0.026225367122018266, 32'sd0.010506045498260067, 32'sd-0.04927056751569848, 32'sd-0.018118594872917938, 32'sd-0.038130051859286106, 32'sd0.1382359017479481, 32'sd0.1335512661464958, 32'sd0.01702131363082135, 32'sd0.014220949452398619, 32'sd0.10617545838741374, 32'sd0.1164867030478873, 32'sd-0.032738614094373925, 32'sd-0.11219547278990907, 32'sd-0.08859868756970316, 32'sd-0.002488057301464197, 32'sd-0.1482654008297202, 32'sd-0.058613012011924884, 32'sd-0.02556973625839405, 32'sd-6.305505082362219e-118, 32'sd0.005217165044392624, 32'sd0.07396785176755999, 32'sd-0.029509744707773945, 32'sd0.010416359928769325, 32'sd-0.09113360562704606, 32'sd0.06312636516064629, 32'sd-0.045295835788994605, 32'sd0.004555626168091302, 32'sd0.016081100223743823, 32'sd-0.029944770641599287, 32'sd-0.06444136775063916, 32'sd-0.23151265184745826, 32'sd-0.1381323049320601, 32'sd-0.05818576045148905, 32'sd0.11843563064910592, 32'sd0.0823103951527102, 32'sd0.16946244457510812, 32'sd0.13395420146952897, 32'sd0.1330232279332569, 32'sd-0.007839157525068374, 32'sd-0.022921219491542338, 32'sd0.08224617424904923, 32'sd-0.14981714273145916, 32'sd-0.07919797310011666, 32'sd-0.04724499470244385, 32'sd0.007265764435867425, 32'sd0.02506764655319669, 32'sd0.019026273973654584, 32'sd-0.08872443490183157, 32'sd-0.03636140721037463, 32'sd0.017433037986796403, 32'sd-0.012642975230097126, 32'sd-0.034323028751692915, 32'sd-0.04984074296668387, 32'sd-0.14353598258899114, 32'sd-0.04687737621385207, 32'sd-0.06890002800197177, 32'sd-0.07849956418559602, 32'sd-0.06540267048214121, 32'sd-0.10644330939528217, 32'sd-0.18514584715298016, 32'sd0.07263926378990221, 32'sd0.032743944288113114, 32'sd0.07507287908566948, 32'sd0.08777984305282552, 32'sd0.08544495320045987, 32'sd0.04295566263119038, 32'sd0.14374150761328747, 32'sd-0.00204479980618944, 32'sd0.07041361374055348, 32'sd-0.16840015033706188, 32'sd-0.05213372331298088, 32'sd-0.02598728435223915, 32'sd0.004914341732862224, 32'sd-0.04345643107455931, 32'sd-0.020649938274436785, 32'sd-0.015300247234979875, 32'sd0.020745489387731197, 32'sd-0.03746005001492879, 32'sd0.053536709885982844, 32'sd0.031084943630405627, 32'sd-0.011003872829257993, 32'sd-0.12930432558505092, 32'sd-0.026468716131923708, 32'sd-0.08108185942526697, 32'sd0.0275414261057279, 32'sd-0.0812396345061743, 32'sd-0.13617227714882757, 32'sd-0.15772169946534936, 32'sd0.06664037217526356, 32'sd-0.06335106966916437, 32'sd0.13479756860339792, 32'sd0.146585580641731, 32'sd0.11938969044689546, 32'sd0.009690662907681344, 32'sd0.059823577513551905, 32'sd-0.02389663288540753, 32'sd0.012472087393186155, 32'sd-0.048120747079778786, 32'sd0.014272800969927248, 32'sd-0.06201278845646037, 32'sd0.05102342367321694, 32'sd-0.03976794563219833, 32'sd2.763584803138982e-122, 32'sd0.010449706010387878, 32'sd0.007708497781371732, 32'sd0.027047296488761197, 32'sd0.014973906620283367, 32'sd0.07023166972757361, 32'sd0.012051005864219928, 32'sd-0.07419582726319829, 32'sd0.0027276993352572817, 32'sd-0.121047916805311, 32'sd-0.11352477392604313, 32'sd-0.03114486084141565, 32'sd-0.02355720183726784, 32'sd-0.047865765760797624, 32'sd0.0005674542116092914, 32'sd0.032242484281153415, 32'sd0.11727664500227344, 32'sd0.13960299397901763, 32'sd0.06950210052082106, 32'sd0.061065524667807056, 32'sd0.028037838174474305, 32'sd-0.06420227757140262, 32'sd-0.1011142397595631, 32'sd-0.02569210711473653, 32'sd-0.03887662010765488, 32'sd-0.0033768178943003116, 32'sd0.005927362165419101, 32'sd3.485250083067307e-115, 32'sd-3.623180255292886e-123, 32'sd-4.0499331015806465e-119, 32'sd-0.07332765733367079, 32'sd0.014282497522317842, 32'sd0.05317061160655598, 32'sd-0.08510163013649429, 32'sd-0.12618937511431869, 32'sd-0.0827533052241464, 32'sd-0.09009789961037905, 32'sd-0.07776535478788744, 32'sd-0.022990781169211674, 32'sd-0.06806151649157573, 32'sd-0.10738105622676963, 32'sd0.07037159631912068, 32'sd0.010359603970967479, 32'sd0.0524183714191264, 32'sd0.11889427927738358, 32'sd0.12478709748699843, 32'sd0.03512724438231269, 32'sd0.07509011499727077, 32'sd-0.05270650768171884, 32'sd-0.15367379443150428, 32'sd-0.013749337693975613, 32'sd-0.016490758486485072, 32'sd0.02482170988292657, 32'sd-0.01248879312143794, 32'sd0.013197134459957299, 32'sd-2.977802579297816e-119, 32'sd-1.5287345596361071e-115, 32'sd-4.0387776807655147e-115, 32'sd-0.051088053553885106, 32'sd0.04191981538560272, 32'sd-0.020782981398124453, 32'sd0.020276809112042146, 32'sd0.05270866768031628, 32'sd-0.06600362805278276, 32'sd-0.06342931504906997, 32'sd0.11849254763834283, 32'sd0.008171941229847659, 32'sd0.0034752265533505794, 32'sd-0.03475430478082574, 32'sd0.002833899262290936, 32'sd0.022481353447735913, 32'sd0.12268788605288036, 32'sd0.21194715057892383, 32'sd0.07619108863996622, 32'sd0.031006696371048192, 32'sd-0.10810320263224983, 32'sd-0.01591891428749596, 32'sd0.037523573292838196, 32'sd0.04294948688108925, 32'sd-0.009680565109923567, 32'sd-0.0006030117809591617, 32'sd0.01693027714427027, 32'sd-0.029841468891787765, 32'sd-9.09315589969163e-120, 32'sd-1.3967612990515953e-115, 32'sd-7.94065979736283e-126, 32'sd5.915458116300997e-125, 32'sd0.008833632549427553, 32'sd-0.052239822765769134, 32'sd0.05587753700418194, 32'sd-0.04019800945181907, 32'sd-0.03378868542051434, 32'sd-0.009410030942915516, 32'sd0.014340569212369701, 32'sd-0.16717887783353294, 32'sd0.03640137479568732, 32'sd-0.017876437034566865, 32'sd0.008226079691470836, 32'sd-0.03959618728918927, 32'sd0.04013994967363968, 32'sd0.04343569143202467, 32'sd-0.12055579293097506, 32'sd-0.10617187904122248, 32'sd0.056031185411477676, 32'sd0.02742354472367467, 32'sd0.015428353778031688, 32'sd-0.023827153141076057, 32'sd0.0551437108357668, 32'sd0.07944441346435739, 32'sd-0.0325630219529955, 32'sd-1.7191415698552917e-124, 32'sd-2.1153110223132922e-117, 32'sd-5.146152353721481e-116, 32'sd9.560444640817624e-119, 32'sd-3.5722096439340115e-116, 32'sd1.5976469768401038e-127, 32'sd-0.01846082017595039, 32'sd0.0601754661857026, 32'sd0.05868308970799557, 32'sd0.04859190368576722, 32'sd-0.0004929689086773329, 32'sd0.0034082777752694627, 32'sd0.035960315068877695, 32'sd-0.07198102444449891, 32'sd0.006385369326128942, 32'sd-0.03457330733616617, 32'sd-0.019940559310044466, 32'sd0.11031882521207938, 32'sd-0.07598120735448545, 32'sd0.03762503466136913, 32'sd0.03565498915569396, 32'sd0.02263707186820634, 32'sd-0.09327960699165347, 32'sd-0.001957291539769532, 32'sd-0.01804384472954346, 32'sd-0.008821568299879137, 32'sd1.942577014913977e-114, 32'sd-3.482573427356277e-124, 32'sd3.2931759583398983e-122, 32'sd-6.412739568863544e-117},
        '{32'sd7.138501373986991e-116, 32'sd3.837734569519557e-122, 32'sd1.6098785513059131e-125, 32'sd-1.3174523302605917e-118, 32'sd3.701318381935605e-122, 32'sd1.707626160865914e-126, 32'sd1.8049416289955916e-119, 32'sd-1.9738648655502875e-114, 32'sd3.936804307366972e-119, 32'sd1.2195144757896913e-125, 32'sd-8.252889521511515e-125, 32'sd-1.3162988074280062e-122, 32'sd0.03218991897049938, 32'sd0.13631495064202148, 32'sd0.06707897922781718, 32'sd0.10085246497782789, 32'sd2.6395893172485394e-124, 32'sd1.112011620693792e-121, 32'sd-7.806689096572031e-125, 32'sd-1.5006693331893555e-126, 32'sd-6.115587951430202e-120, 32'sd1.2006461400359483e-123, 32'sd3.555734837585929e-116, 32'sd-1.0375541482792193e-115, 32'sd-2.8346839512457843e-118, 32'sd-3.2862528923565606e-114, 32'sd5.5491696417090815e-121, 32'sd1.444480611461718e-122, 32'sd-1.9428590632385676e-114, 32'sd-1.494897866492916e-124, 32'sd-1.0488644679304397e-120, 32'sd-2.7769330877372147e-123, 32'sd0.027149040616254862, 32'sd0.11646703839391921, 32'sd0.0795894855576865, 32'sd0.10357883123576779, 32'sd0.05916619406166681, 32'sd0.1075113046554639, 32'sd0.12553517282072266, 32'sd0.0589318444510614, 32'sd0.020975763226452875, 32'sd-0.026026372113861208, 32'sd-0.09313494316909002, 32'sd0.05428102377104427, 32'sd0.13466775099603623, 32'sd0.1316919515344549, 32'sd0.08894656888290453, 32'sd0.03605158880148624, 32'sd-0.011513644921985096, 32'sd-0.012381442998864726, 32'sd0.08589396952335916, 32'sd0.04006032222463899, 32'sd-4.546944245807245e-126, 32'sd5.844273400666575e-124, 32'sd-1.9348075195318287e-124, 32'sd1.1187338211662645e-115, 32'sd-1.2932862534329132e-125, 32'sd1.1356859375122835e-123, 32'sd0.06841679222959367, 32'sd-0.02420356763472678, 32'sd-0.001418101096996707, 32'sd0.08780965257402065, 32'sd0.026615352401532868, 32'sd-0.025238999258084965, 32'sd0.060525913631106466, 32'sd0.08328390982207658, 32'sd0.034661469665012955, 32'sd-0.03269405570837829, 32'sd-0.06791943819865516, 32'sd-0.042898930135339845, 32'sd0.021317267892250063, 32'sd0.04496798953106999, 32'sd0.04994451135033937, 32'sd0.05879186315754359, 32'sd0.020275365272529558, 32'sd0.2264037398213571, 32'sd0.17997358569894656, 32'sd0.07277602640961106, 32'sd-0.00538457759120818, 32'sd0.146511626130886, 32'sd0.006115936439912275, 32'sd0.08457048301606883, 32'sd-2.921656693745396e-125, 32'sd2.45188926014243e-126, 32'sd-1.3237703711245271e-125, 32'sd9.343985776869991e-123, 32'sd-0.020945694003374097, 32'sd0.03336294408973794, 32'sd-0.008113451056974202, 32'sd-0.005006807205035531, 32'sd-0.03981591410827414, 32'sd-0.1250431359218275, 32'sd-0.04556087186431076, 32'sd0.0738489337949658, 32'sd0.005865336211214502, 32'sd0.0688478549929626, 32'sd-0.01604307375125709, 32'sd0.07883241309371154, 32'sd0.0005086937877656044, 32'sd-0.05967180865018827, 32'sd-0.045785240205458315, 32'sd0.015209565034928483, 32'sd0.0664350124476987, 32'sd0.06031622925769206, 32'sd0.04153364579682099, 32'sd0.0054036522633600865, 32'sd-0.04091853795301959, 32'sd-0.1621823289923645, 32'sd-0.06583180194557255, 32'sd-0.06984882829081257, 32'sd0.0511920683980931, 32'sd3.57209682438384e-114, 32'sd3.9080381357882526e-116, 32'sd0.05195797951908102, 32'sd0.03109665037048798, 32'sd-0.0003571172943889219, 32'sd-0.022451277968799123, 32'sd-0.03744073403138433, 32'sd-0.14123778472668302, 32'sd-0.11483248713505632, 32'sd-0.09670753555999584, 32'sd-0.06741273201057128, 32'sd-0.053825869857105475, 32'sd0.06294184850067214, 32'sd0.03392983795132466, 32'sd-0.017489634234454158, 32'sd-0.0709290516745213, 32'sd-0.06653718325540828, 32'sd-0.07879284077665845, 32'sd-0.06908188814677829, 32'sd-0.04356858499263641, 32'sd-0.011142189429771356, 32'sd-0.11281159196608376, 32'sd-0.02949915544903118, 32'sd-0.06907009335448688, 32'sd0.028222821241544672, 32'sd0.01071876422231499, 32'sd0.06072230909408265, 32'sd0.0818862523541891, 32'sd0.0475088977660176, 32'sd2.6020505490948823e-126, 32'sd0.051817574250369, 32'sd-0.044516160021828795, 32'sd-0.006659363453985718, 32'sd-0.09641705878297688, 32'sd-0.08730436583307531, 32'sd-0.028979981872945756, 32'sd-0.14847825683993685, 32'sd-0.10270814255939832, 32'sd-0.11172486326790768, 32'sd0.015954186949937266, 32'sd0.027346041205791774, 32'sd-0.012168607332258533, 32'sd0.018174308406606266, 32'sd0.028818423757022628, 32'sd0.0046899756074239, 32'sd-0.01829387725957533, 32'sd0.03740852606971915, 32'sd-0.0025036591724702673, 32'sd0.07327510761492753, 32'sd0.11023829098718553, 32'sd0.12463133356385761, 32'sd0.039596086834509034, 32'sd-0.01738731042323498, 32'sd0.12449563303346088, 32'sd0.12473619443442353, 32'sd0.1320233357837461, 32'sd-0.06508425026382357, 32'sd-5.406080248580773e-118, 32'sd0.03266425639763329, 32'sd-0.051532525427556757, 32'sd-0.027267190634651602, 32'sd-0.13065614192956426, 32'sd-0.059489775666888144, 32'sd-0.0757144126993444, 32'sd0.006875691926891667, 32'sd-0.12707408407961068, 32'sd-0.1744439513146849, 32'sd-0.009009800369923174, 32'sd0.10310999393796182, 32'sd0.007354787186986946, 32'sd-0.016775540267915633, 32'sd0.039875615676864345, 32'sd-0.017683626119836336, 32'sd0.07392600637068704, 32'sd0.10039055623975993, 32'sd0.10890438402411111, 32'sd0.08305345167840289, 32'sd0.10307648869901938, 32'sd0.02289606114155606, 32'sd0.0005253963841150985, 32'sd-0.010534009639853546, 32'sd-0.00791463088610067, 32'sd-0.03910198696506865, 32'sd0.04775983433740066, 32'sd-0.014676941770320789, 32'sd0.10135690923214931, 32'sd-0.06569365367703298, 32'sd-0.01351449493449778, 32'sd0.02262159794538734, 32'sd-0.09636775387942179, 32'sd-0.0439306590834708, 32'sd0.08884807450874123, 32'sd-0.08580681533477985, 32'sd-0.042785181365561704, 32'sd-0.018286805062335584, 32'sd0.05385734489848973, 32'sd0.07409108675265516, 32'sd-0.13517796150123643, 32'sd-0.11308456906289867, 32'sd-0.012861836026252719, 32'sd-0.09526657420025851, 32'sd-0.10388623569157743, 32'sd0.011675258750859186, 32'sd-0.05234747010655555, 32'sd0.14277317713111845, 32'sd0.062423236290482506, 32'sd0.05499311946968554, 32'sd0.17261973262112054, 32'sd-0.027636663620069515, 32'sd-0.024418782690051512, 32'sd0.013839893261997437, 32'sd-0.07086057427747622, 32'sd-0.016809880536847264, 32'sd-0.0011960861096669145, 32'sd0.02345350092815103, 32'sd0.08055734547647006, 32'sd-0.0637404861034762, 32'sd-0.11241308895133949, 32'sd0.01686514583093239, 32'sd-0.0238412918683424, 32'sd-0.034470599203241296, 32'sd-0.08731253623099886, 32'sd-0.06040539471281117, 32'sd0.07875345780160628, 32'sd0.11080350796651345, 32'sd-0.07776602085122582, 32'sd-0.11340257371250587, 32'sd-0.05948509840886741, 32'sd-0.12531420842910515, 32'sd-0.011057696476556625, 32'sd-0.005201765401978335, 32'sd-0.042482919139447246, 32'sd0.06462320501430208, 32'sd0.18694991901026287, 32'sd0.051318616805891504, 32'sd0.08162371750352815, 32'sd0.06808828823378815, 32'sd-0.04088028311232848, 32'sd0.03596466001415947, 32'sd-0.04504337147782993, 32'sd-0.012395527609949475, 32'sd0.04469020209005146, 32'sd-0.020033867799168163, 32'sd-0.03588765490862301, 32'sd0.16745093458823557, 32'sd0.21068736923078044, 32'sd0.1404654472158475, 32'sd0.09744748542038857, 32'sd0.0025660033141539675, 32'sd-0.005380339897903096, 32'sd0.003892758575142353, 32'sd-0.015776735735636576, 32'sd0.06081057720434717, 32'sd-0.10642866101097359, 32'sd-0.09650764611012141, 32'sd-0.0251454660295399, 32'sd-0.21512457823538045, 32'sd-0.24394367578473894, 32'sd-0.18706515812737828, 32'sd0.04862544044838026, 32'sd0.0665638886317877, 32'sd0.11989754785120242, 32'sd0.081463549110011, 32'sd0.10933652505580681, 32'sd0.05968943449651609, 32'sd-0.015097604324649534, 32'sd0.09255571567931449, 32'sd0.03350167365778436, 32'sd-0.050209905272130456, 32'sd-0.012422878498546914, 32'sd0.004354848312411322, 32'sd0.06496474327951192, 32'sd0.0026592421928039603, 32'sd0.06545494109407295, 32'sd0.12446249198617626, 32'sd-0.009925212001159346, 32'sd-0.02167510310167645, 32'sd0.030369600930239143, 32'sd0.11170555190999666, 32'sd0.13458794310133265, 32'sd0.17412418646664898, 32'sd0.07038674904831042, 32'sd0.02815117850444865, 32'sd-0.0633578214342412, 32'sd-0.06184570179842176, 32'sd-0.08433387437166935, 32'sd-0.12361164398361238, 32'sd-0.011379373418144444, 32'sd-0.005641118236614081, 32'sd0.08104298886810307, 32'sd0.01010058785542322, 32'sd0.13545569462893328, 32'sd0.08970177797847359, 32'sd-0.06608247780318344, 32'sd-0.038587326483130006, 32'sd-0.07501278807208342, 32'sd0.0016709741289594685, 32'sd0.030231443574244045, 32'sd0.10327081698973686, 32'sd0.09440105342799246, 32'sd0.03885701977553122, 32'sd0.07349179627671046, 32'sd0.002640214318556338, 32'sd-0.07862778518698643, 32'sd0.09825548695934519, 32'sd-0.030769503271745456, 32'sd0.11412103433232826, 32'sd0.09491418118714055, 32'sd0.004516410163919322, 32'sd0.030846776757096874, 32'sd0.11267674604626622, 32'sd0.06282671439188758, 32'sd-0.07200640974466113, 32'sd-0.12412554580346542, 32'sd-0.15080930862674838, 32'sd-0.07773638570871684, 32'sd0.010777295931159904, 32'sd0.04195975629128039, 32'sd0.03767222937342305, 32'sd0.16069299152780964, 32'sd0.07765080256252398, 32'sd0.04352946839498225, 32'sd0.08907222533081231, 32'sd0.06569011635299417, 32'sd0.0607282205557595, 32'sd0.06940551607878132, 32'sd0.048949265899343744, 32'sd-0.017220308192866726, 32'sd-0.007924301781496071, 32'sd0.02078541312014835, 32'sd-0.08060929818107697, 32'sd0.05809009918025741, 32'sd0.14025117308553434, 32'sd0.060195364293704326, 32'sd0.12357635686381507, 32'sd0.06338039905861755, 32'sd0.05451736410274231, 32'sd-0.009149799523180121, 32'sd-0.09899313495123134, 32'sd-0.16906417869536586, 32'sd-0.07110348907137425, 32'sd-0.15228259356556467, 32'sd-0.17836597576939436, 32'sd-0.1144360007192792, 32'sd-0.1010293347825241, 32'sd0.020800780372166344, 32'sd-0.0530084916805408, 32'sd0.022284814285882568, 32'sd0.07864110943227112, 32'sd0.007197060521224553, 32'sd-0.02293042630526741, 32'sd0.014189143543505206, 32'sd0.1327540616359948, 32'sd0.059960747687751656, 32'sd-0.004712811365081824, 32'sd-0.08293401285432868, 32'sd-0.13417993647253407, 32'sd0.02455914075821497, 32'sd0.017609404494557997, 32'sd0.07916713894621291, 32'sd0.048079564195742275, 32'sd-0.015110767045982187, 32'sd-0.042788227071620215, 32'sd-0.0404129726407363, 32'sd-0.06667596664949858, 32'sd-0.1330172057927784, 32'sd-0.03050610891579629, 32'sd-0.10369874106390375, 32'sd-0.166627466039233, 32'sd-0.013213196921526879, 32'sd-0.08601893504269534, 32'sd-0.13299306050667886, 32'sd-0.06040705756957847, 32'sd0.017146151554923262, 32'sd-0.0035146124182325942, 32'sd-0.05097279685299033, 32'sd-0.026082684539184428, 32'sd0.12988517221846013, 32'sd0.05028880939456192, 32'sd0.11851466331663885, 32'sd0.17207141915736052, 32'sd0.07085404538542515, 32'sd-0.05407418047136931, 32'sd-0.012810325252739153, 32'sd-0.14833672047741614, 32'sd-0.02838196881286896, 32'sd0.04797056185826179, 32'sd-0.07178011701905432, 32'sd-0.016547908943828914, 32'sd0.0038297072608852656, 32'sd-0.12537178544479027, 32'sd-0.08538179612024485, 32'sd-0.156101818693293, 32'sd-0.1092516236997744, 32'sd-0.12806544596439323, 32'sd-0.04752715357939157, 32'sd-0.1712735381852906, 32'sd-0.15143921783464118, 32'sd0.10171845531353559, 32'sd0.05400365079036827, 32'sd-0.02299459135734753, 32'sd0.10278679461197898, 32'sd-0.02308587167853679, 32'sd-0.005001743055074054, 32'sd0.04414410881352568, 32'sd-0.011616607560515694, 32'sd0.045947300771291985, 32'sd-0.06521919763413928, 32'sd0.1731290249687433, 32'sd0.06255953164479867, 32'sd0.03185310939710549, 32'sd-0.02050659754078115, 32'sd-0.023454431010412648, 32'sd0.045308199798349484, 32'sd-0.0227010271904844, 32'sd-0.007105597962721783, 32'sd-0.043944237105022925, 32'sd-0.011111614397954044, 32'sd0.019292000071548108, 32'sd-0.10024363796293517, 32'sd-0.01657517478440267, 32'sd-0.12256666700964307, 32'sd-0.03777249870495235, 32'sd-0.05384407385814424, 32'sd-0.07112962055743974, 32'sd-0.054489262433407265, 32'sd0.09505306581013963, 32'sd0.06869481493745008, 32'sd0.12288400501652877, 32'sd0.005320627886195044, 32'sd-0.00888883529523982, 32'sd-0.053632984549259834, 32'sd-0.008406398319946055, 32'sd-0.0033487815415445396, 32'sd-0.08574928649243341, 32'sd0.027608050091979145, 32'sd0.04722969825087414, 32'sd0.06019302076172298, 32'sd-0.07068198456072855, 32'sd-0.013605176031741216, 32'sd0.045253494004397585, 32'sd-0.03760461359346278, 32'sd0.10273788497628639, 32'sd0.08114403027959267, 32'sd0.11562697837956543, 32'sd-0.001610458170654582, 32'sd0.014357067388428678, 32'sd0.027817438646321017, 32'sd0.020425468277402895, 32'sd-0.10083056193683486, 32'sd0.0030744394823675613, 32'sd-0.0599117306645955, 32'sd-0.032658846732111925, 32'sd-0.05143880627210255, 32'sd0.1600482411871749, 32'sd0.009442281581315262, 32'sd0.053855447872120106, 32'sd0.09813286709119502, 32'sd0.011992224095571135, 32'sd-0.04348557442600051, 32'sd-0.028172257900265618, 32'sd-0.03704680517960436, 32'sd0.07227417107961355, 32'sd0.07562676959439138, 32'sd0.10436978151068552, 32'sd7.998194883926426e-123, 32'sd0.0528640873932095, 32'sd-0.07416088330819266, 32'sd-0.031166893093313858, 32'sd0.1259835824578126, 32'sd0.12642854925029057, 32'sd-0.0005962641209960346, 32'sd0.12396296175448202, 32'sd0.011495541900840175, 32'sd0.10982120014805313, 32'sd-0.05994961283342024, 32'sd-0.0825966894129165, 32'sd-0.08409968338904385, 32'sd-0.0051430265425295935, 32'sd0.049964938978353024, 32'sd-0.02106168431764133, 32'sd-0.010123559302817813, 32'sd0.0776298677163685, 32'sd0.08391033017458192, 32'sd-0.09471501216379742, 32'sd0.06470826783257627, 32'sd-0.05897682909835366, 32'sd-0.03648157680214019, 32'sd0.03218218906704209, 32'sd0.06859570408471416, 32'sd0.07922662360120938, 32'sd-0.038811841777710354, 32'sd0.005215938910787416, 32'sd-0.01966855281435698, 32'sd0.05376513659733018, 32'sd0.041826028640672676, 32'sd-0.09367313636329616, 32'sd0.0919929420741016, 32'sd0.10976643088395845, 32'sd-0.022449577179147903, 32'sd0.08454592037966294, 32'sd0.0662526041469355, 32'sd0.014436240041368436, 32'sd-0.17774727967092274, 32'sd-0.12962845818836619, 32'sd-0.18403128086281034, 32'sd-0.061985569791190534, 32'sd0.013792632139975032, 32'sd-0.054003275935672425, 32'sd-0.11778257396200985, 32'sd-0.008680635077791484, 32'sd0.04811145969701385, 32'sd-0.14452194058047946, 32'sd0.035582131952049345, 32'sd0.019701223041508207, 32'sd-0.06508470882551848, 32'sd0.05775498091033001, 32'sd0.009119325096754767, 32'sd-0.018700511175892484, 32'sd-0.01925515502239202, 32'sd0.11038837479006229, 32'sd0.05241476372607315, 32'sd-0.06768323497728869, 32'sd0.0259415737700264, 32'sd-0.07190194066472047, 32'sd0.12041789115936795, 32'sd0.10850198277157828, 32'sd0.002575360887557016, 32'sd0.03186672019896165, 32'sd0.11891257271407106, 32'sd0.11497198132623968, 32'sd-0.09591641723582423, 32'sd-0.12553567444082606, 32'sd-0.008920962072133186, 32'sd-0.05878007770775063, 32'sd-0.08803629985603156, 32'sd-0.050849834665855284, 32'sd-0.015125410398034328, 32'sd-0.01777849379008178, 32'sd-0.08139592500172949, 32'sd-0.03779440155323495, 32'sd-0.0835079837983238, 32'sd-0.008927540307613018, 32'sd-0.0717001606034561, 32'sd-0.004868377072664232, 32'sd-0.04514594202261929, 32'sd-0.011710653830865602, 32'sd-0.08543898127165006, 32'sd-0.035432946676774414, 32'sd-5.5284805348077e-119, 32'sd-0.017184354395489813, 32'sd0.019295052410880933, 32'sd0.030281886104148826, 32'sd0.1098835595357062, 32'sd0.14068124440621085, 32'sd0.10641651306823173, 32'sd0.16254305913640632, 32'sd0.05966843044465242, 32'sd-0.04410249223740903, 32'sd-0.03433942725436674, 32'sd0.024670062032394826, 32'sd-0.09390676602186335, 32'sd-0.07872432844237892, 32'sd-0.11645421325737611, 32'sd-0.17015700886109517, 32'sd-0.15684590907049764, 32'sd-0.1440811756068904, 32'sd-0.10030544047225945, 32'sd0.008086963816313367, 32'sd-0.030629890753232244, 32'sd-0.06463778660962557, 32'sd-0.04612797819230738, 32'sd-0.06065480172194163, 32'sd-0.04660377997322649, 32'sd-0.08370108520575821, 32'sd-0.08742124792550479, 32'sd0.05731898586055989, 32'sd0.06280318855167216, 32'sd0.022425884625978297, 32'sd-0.0048188597479801075, 32'sd0.02050839819824324, 32'sd0.03213519720581363, 32'sd0.09479458812145543, 32'sd0.12771661141569676, 32'sd0.1283912592010945, 32'sd0.10292361591680738, 32'sd0.0034686632767002685, 32'sd-0.03502127389441882, 32'sd0.02746698010390724, 32'sd-0.06111860771255619, 32'sd-0.06668834696519098, 32'sd-0.0673902783724807, 32'sd0.001351374842887698, 32'sd-0.06142294708529598, 32'sd0.03548116088400715, 32'sd-0.06927897799761006, 32'sd-0.06277110180772251, 32'sd-0.03200017859043782, 32'sd0.013541717715949054, 32'sd0.041824729036090975, 32'sd-0.03178000035149743, 32'sd0.00018605439028741632, 32'sd-0.039304813801719504, 32'sd0.050527853304738746, 32'sd0.06993393187170627, 32'sd0.07789196511209776, 32'sd0.018538398361575063, 32'sd-0.010783484832631775, 32'sd0.10458245745585579, 32'sd-0.010176344673125172, 32'sd0.020630624867613516, 32'sd0.2020220656029877, 32'sd0.11581043607924604, 32'sd0.015975866149220832, 32'sd-0.05892588935370551, 32'sd-0.015216329161312318, 32'sd0.03208856970945215, 32'sd0.05513274260097463, 32'sd-0.09547461044582047, 32'sd-0.06425269980889932, 32'sd-0.008773701208563679, 32'sd0.03295793029639384, 32'sd-0.03254472416332129, 32'sd-0.08812935980761394, 32'sd-0.02053541718463582, 32'sd-0.029135769694719732, 32'sd0.024994605436556832, 32'sd-0.06140404958117898, 32'sd-0.14229229947208302, 32'sd-0.03662485821657461, 32'sd-0.010349716934162973, 32'sd0.039109919572400856, 32'sd0.1210399650613784, 32'sd2.2322157576978884e-116, 32'sd0.053254130928980986, 32'sd0.10729473221921998, 32'sd0.10968832510475102, 32'sd0.014952307831851275, 32'sd-0.035163362424212294, 32'sd0.09601571654052174, 32'sd0.11744889362299579, 32'sd0.1426125186427435, 32'sd-0.03071329340092734, 32'sd0.05453963092826204, 32'sd-0.04270069704148646, 32'sd-0.08688644110958091, 32'sd-0.0408342408200215, 32'sd-0.05912612770620047, 32'sd0.0031621288571911624, 32'sd0.005372484872157747, 32'sd0.06311982143707127, 32'sd0.013870040356190499, 32'sd0.008352894600800752, 32'sd0.03124709540426026, 32'sd-0.09398160915276305, 32'sd-0.003338386399644544, 32'sd-0.04070484685981442, 32'sd0.035408851934066524, 32'sd-0.015012709220582942, 32'sd-0.006947917613818706, 32'sd1.5504676600262873e-116, 32'sd3.061200783103999e-119, 32'sd-8.703133531619133e-126, 32'sd0.022742942356731344, 32'sd0.07355038357050037, 32'sd0.13928216158896273, 32'sd0.013874859788990786, 32'sd0.024930846595168768, 32'sd0.11306774919149218, 32'sd0.14514749883228842, 32'sd0.03212325018679751, 32'sd0.07222170580102359, 32'sd0.004891453386211958, 32'sd0.038834230785004316, 32'sd0.02138399574871688, 32'sd-0.12823990505656305, 32'sd-0.07465788218970014, 32'sd-0.09789693851472688, 32'sd-0.03984901808969797, 32'sd0.03671165762478973, 32'sd0.03509811384824873, 32'sd0.0315375839378805, 32'sd0.03471188629234819, 32'sd-0.014099951081627952, 32'sd0.03277138141849422, 32'sd-0.0616544363503345, 32'sd0.06378528827131222, 32'sd0.04403146640438778, 32'sd-1.1360058769437797e-119, 32'sd8.15638012522093e-120, 32'sd-7.351813559129631e-116, 32'sd-0.07046731877537338, 32'sd-0.011526341543540227, 32'sd-0.027311952694632026, 32'sd-0.1067106802921164, 32'sd-0.10651566627237825, 32'sd-0.034547687304185705, 32'sd0.050560149029189955, 32'sd0.08394683684853774, 32'sd0.08125653782526993, 32'sd-0.04095613103013761, 32'sd0.026280461670083303, 32'sd0.0491827175531972, 32'sd0.08158211809077032, 32'sd-0.025580445193097517, 32'sd0.0656314207882558, 32'sd-0.07378126356807219, 32'sd-0.042712249023183976, 32'sd0.12530123128018372, 32'sd0.04376951025042488, 32'sd0.08686681936335694, 32'sd-0.07312314031466613, 32'sd0.051985010674397036, 32'sd-0.016346077188574473, 32'sd0.05713516938902734, 32'sd0.10394659674494329, 32'sd7.12998110833296e-117, 32'sd8.594042299983845e-120, 32'sd2.979963337357181e-116, 32'sd2.9851181784648234e-122, 32'sd0.09324501898135085, 32'sd0.021760000459542798, 32'sd-0.10513730606776135, 32'sd-0.04200668825890999, 32'sd-0.058924638507487165, 32'sd-0.02054332373552049, 32'sd0.03505766581044389, 32'sd0.06316666626468545, 32'sd0.0024664906937951468, 32'sd0.07200591029231475, 32'sd-0.07464512647802246, 32'sd-0.019752086213659877, 32'sd-0.04501985322873238, 32'sd0.1216543526971981, 32'sd0.017173742928513862, 32'sd0.0787750629557812, 32'sd0.0893558132332784, 32'sd0.00035099175399729173, 32'sd-0.03304646345739769, 32'sd0.14417276845849564, 32'sd0.08576288878884843, 32'sd-0.02345216098439962, 32'sd0.10490909410869152, 32'sd6.567722238412016e-125, 32'sd-1.4550174962541212e-115, 32'sd-1.6188202114270916e-115, 32'sd-1.5590073570072602e-124, 32'sd1.5880089104102946e-115, 32'sd-1.1379004393496487e-118, 32'sd0.10187602321869278, 32'sd0.05921501927088091, 32'sd0.027978612925147195, 32'sd0.07829118337344783, 32'sd0.00233777175976271, 32'sd-0.008857300030579074, 32'sd0.09903870663679593, 32'sd-0.014538579467757351, 32'sd0.08249015818845679, 32'sd0.04678053838394345, 32'sd0.11628642013001454, 32'sd0.08402307768317298, 32'sd0.01452428704356251, 32'sd0.039401254427512605, 32'sd0.04967460389290843, 32'sd-0.06308002404780234, 32'sd0.01105421727854916, 32'sd0.012808856231956288, 32'sd0.05920566635060326, 32'sd0.09117771433518199, 32'sd-6.953659191220768e-124, 32'sd-2.6418142378160334e-120, 32'sd1.8171685704097452e-123, 32'sd2.65884854218433e-118},
        '{32'sd3.247985268729037e-127, 32'sd3.6914323716422527e-121, 32'sd-1.074922773528862e-124, 32'sd2.3032614206298987e-119, 32'sd5.045820067576413e-126, 32'sd-1.0695477329299472e-126, 32'sd-8.199210892890103e-119, 32'sd-3.511279148130579e-119, 32'sd1.3451542971744494e-120, 32'sd-1.1149989495258666e-114, 32'sd3.546838000962273e-116, 32'sd1.454152016579461e-122, 32'sd-0.005865248950561107, 32'sd-0.015514086501169888, 32'sd-0.017650823732644493, 32'sd-0.0003481728104924093, 32'sd3.494187805718951e-122, 32'sd1.199750675709981e-124, 32'sd1.087798274584882e-118, 32'sd5.3958707139940045e-126, 32'sd1.7175374207941153e-125, 32'sd-4.9206295203212756e-120, 32'sd6.893645487137205e-126, 32'sd1.808808265009036e-123, 32'sd-4.788696567028699e-118, 32'sd5.707019116130591e-127, 32'sd5.509786882437783e-117, 32'sd6.703893486981318e-121, 32'sd-5.180484619262813e-124, 32'sd6.544151130688874e-121, 32'sd-1.8808466124153162e-121, 32'sd1.7256854933590516e-123, 32'sd0.04323302856689574, 32'sd-0.05410479494107593, 32'sd-0.01183985855328643, 32'sd0.030800979842390535, 32'sd0.004969416748962012, 32'sd0.0035591702227867252, 32'sd0.10713831305854213, 32'sd-0.0640460222846808, 32'sd0.0045055550849385385, 32'sd-0.06569304365997072, 32'sd0.0076497566239011015, 32'sd0.007939114738772587, 32'sd0.05403695277077278, 32'sd0.06987765279318184, 32'sd0.06875707315778504, 32'sd-0.04378968894798896, 32'sd0.08724716541497518, 32'sd0.04195113247733533, 32'sd0.10366017379446842, 32'sd0.009507251257781275, 32'sd-4.01483814618275e-120, 32'sd3.943376249860756e-119, 32'sd1.1692617146613262e-122, 32'sd1.778125030062406e-124, 32'sd-3.4596522862495823e-128, 32'sd3.9335656871248064e-115, 32'sd0.06902792736646615, 32'sd0.09586904760302067, 32'sd0.026963407584592976, 32'sd-0.03485641528130304, 32'sd0.017281088069344634, 32'sd-0.04291963198750286, 32'sd-0.014964770644355545, 32'sd-0.04193232925069809, 32'sd0.059722457483996905, 32'sd0.006623170276512349, 32'sd-0.0645330947252073, 32'sd-0.020514447024931593, 32'sd-0.013270521111714801, 32'sd0.09017022430297206, 32'sd0.11069798162504299, 32'sd-0.014526657472025185, 32'sd0.12354917796809103, 32'sd0.21718226737314913, 32'sd0.07756353184000021, 32'sd-0.01712731246102889, 32'sd0.02446546866645794, 32'sd0.09317698814101877, 32'sd-9.354206895585697e-05, 32'sd0.04886658839959218, 32'sd3.2260309514631506e-114, 32'sd8.648430784406425e-120, 32'sd5.1365441307149965e-124, 32'sd-5.5947788088186454e-124, 32'sd0.03328709995342782, 32'sd0.028919979262287242, 32'sd0.02443566376485184, 32'sd-0.0917728738686244, 32'sd-0.08675983609061946, 32'sd-0.020163727953348268, 32'sd-0.05977914413661207, 32'sd0.0736564502494791, 32'sd0.034914883972302024, 32'sd-0.05820697437713929, 32'sd0.04800833243041323, 32'sd0.14245245375048105, 32'sd0.11635803518127764, 32'sd0.08741469651354175, 32'sd0.012505275543750166, 32'sd-0.06848497069404647, 32'sd-0.0077175601479093974, 32'sd-0.026487938307324422, 32'sd-0.08898209383495954, 32'sd-0.031163250820722486, 32'sd0.06520413083891481, 32'sd0.012213483840001984, 32'sd0.059399913192439556, 32'sd0.06818823187022266, 32'sd0.0141000385559706, 32'sd-9.982407094812087e-121, 32'sd2.290165821025725e-116, 32'sd0.010076793276559585, 32'sd0.04076694024201106, 32'sd-0.07957889216959335, 32'sd0.02336029403015119, 32'sd-0.00010232266043551787, 32'sd0.055366462642285535, 32'sd-0.07392794772475614, 32'sd-0.029742887497333302, 32'sd-0.05075942111663692, 32'sd-0.05696725344492039, 32'sd0.07095317959202249, 32'sd0.02637640624652884, 32'sd-0.06332022245930158, 32'sd0.12319312022796715, 32'sd0.17249022505794193, 32'sd-0.047738190821021674, 32'sd-0.022828177789100294, 32'sd-0.06512680432133748, 32'sd-0.041658635890849394, 32'sd-0.04824868259925947, 32'sd0.13020530382656756, 32'sd0.01713505209863687, 32'sd0.11518437769883458, 32'sd-0.04083529079042388, 32'sd0.09804597446077283, 32'sd0.011765945285312199, 32'sd0.042825016202971286, 32'sd-1.4566723977363527e-122, 32'sd0.018667417237626337, 32'sd-0.040184917936725, 32'sd0.011843109710592343, 32'sd-0.023260014233535, 32'sd0.016110197714930274, 32'sd-0.0033146662257103965, 32'sd-0.047792582388392665, 32'sd0.08908060735163528, 32'sd-0.08304154073533554, 32'sd0.0350989576204475, 32'sd0.06463914415382924, 32'sd0.05344408505313756, 32'sd0.09118174933801143, 32'sd-0.011400739212752366, 32'sd0.14053355474058127, 32'sd0.03982240313886924, 32'sd0.05605481934279561, 32'sd0.10599526509291969, 32'sd-0.010571898500452708, 32'sd0.11193735991798054, 32'sd0.040852094502183287, 32'sd0.0336738817703216, 32'sd0.11137591797783092, 32'sd0.09520469773073056, 32'sd0.039293203688053134, 32'sd0.018407516786853585, 32'sd0.048117688907861854, 32'sd5.515962668343717e-124, 32'sd-0.025260632890639654, 32'sd-0.00671654011392812, 32'sd0.06070238138378489, 32'sd0.05053450444252864, 32'sd0.016769087581792602, 32'sd-0.051890569448507534, 32'sd-0.03354198650127286, 32'sd0.13442487228282973, 32'sd0.03386510918019, 32'sd-0.045430327694041865, 32'sd0.11687754141005317, 32'sd0.1262840823097794, 32'sd0.2029183782117394, 32'sd0.08548872831665771, 32'sd0.1887700084312201, 32'sd0.1673790260359044, 32'sd0.13220437974593954, 32'sd0.07595642226505565, 32'sd0.0031348276523765354, 32'sd-0.049692033038475004, 32'sd0.0035887559757736254, 32'sd-0.0017557647616416076, 32'sd-0.1137692367150568, 32'sd-0.08391112534505653, 32'sd-0.07303168387615186, 32'sd-0.041141653352236095, 32'sd0.06354772882425307, 32'sd0.0892082692511578, 32'sd0.059510327216622194, 32'sd0.09042362218382236, 32'sd0.05522205031083057, 32'sd-0.004869056473896865, 32'sd-0.032932441146066055, 32'sd0.014905681782309044, 32'sd-0.007206700684928913, 32'sd0.11967909800817877, 32'sd0.059206240562760006, 32'sd0.06945297348814945, 32'sd0.0920949757546659, 32'sd0.18764656856906525, 32'sd0.15747459254908075, 32'sd0.13784911237225486, 32'sd-0.006010504798294118, 32'sd0.01318243760495122, 32'sd-0.14670552715592272, 32'sd-0.07127095381117991, 32'sd-0.04202713838239608, 32'sd-0.08161949599580487, 32'sd-0.04268481274657694, 32'sd-0.025927287809094333, 32'sd-0.14605950993283232, 32'sd-0.0794282956668106, 32'sd0.07777505906214123, 32'sd-0.07594660136581532, 32'sd0.0018184344971950463, 32'sd0.07553637516570123, 32'sd0.07907096296761884, 32'sd0.016723648930464796, 32'sd-0.06587903341800998, 32'sd-0.15479304843770506, 32'sd0.04347237881605445, 32'sd-0.05173931966830771, 32'sd0.06776999536715726, 32'sd0.10755776394459567, 32'sd0.005261428490605341, 32'sd0.11900024055629665, 32'sd0.1810539129546299, 32'sd0.11257316743509234, 32'sd-0.031240275052537764, 32'sd0.02142879513536706, 32'sd-0.20317176721341937, 32'sd-0.3053668603435115, 32'sd-0.2401717589288569, 32'sd-0.20857350840448485, 32'sd-0.21873759515393315, 32'sd-0.1636702895735138, 32'sd-0.0795779464466483, 32'sd-0.07439287547566203, 32'sd-0.15577332292089188, 32'sd-0.09366758995141336, 32'sd-0.0892265800390938, 32'sd-0.014721604895116727, 32'sd-0.03680613904644329, 32'sd-0.023028449991043577, 32'sd0.11684799292704834, 32'sd0.08351788097450126, 32'sd-0.08485338511562616, 32'sd0.009034411854953463, 32'sd-0.011705349092694555, 32'sd0.1149721050463809, 32'sd-0.011136939745338716, 32'sd0.10717069721947506, 32'sd0.013000267113395693, 32'sd0.08312513410045042, 32'sd0.11038384638379674, 32'sd-0.12286069904495606, 32'sd-0.18496015048189962, 32'sd-0.08325942430785256, 32'sd-0.1391911136823621, 32'sd-0.1933758677164494, 32'sd-0.11373971094514278, 32'sd-0.23685893626330773, 32'sd-0.2906569430900688, 32'sd-0.2635887338610556, 32'sd-0.2303200822792057, 32'sd-0.17859462662323478, 32'sd-0.1902825588684198, 32'sd-0.11388004990760578, 32'sd-0.02057535716349519, 32'sd-0.016637439785566577, 32'sd0.005618880408212001, 32'sd0.0052336027859567836, 32'sd-0.01641276099247288, 32'sd0.08243832748685241, 32'sd-0.07497365165961736, 32'sd-0.08084241035051919, 32'sd0.071130816478013, 32'sd0.08053183647962803, 32'sd0.008569204599770074, 32'sd-0.05621561047716184, 32'sd0.004685488554363382, 32'sd-0.014362542821526998, 32'sd-0.025338549654327747, 32'sd-0.20355181997836472, 32'sd0.002344128438548325, 32'sd0.06345700791084129, 32'sd0.019540835926269366, 32'sd0.08220852474411432, 32'sd0.034443625108611355, 32'sd0.07149904383952096, 32'sd-0.05629525264836227, 32'sd-0.10277981950096549, 32'sd-0.12181808146192535, 32'sd-0.011979590962398872, 32'sd-0.07361594712505103, 32'sd-0.047656571914011514, 32'sd-0.034691612572253394, 32'sd-0.026902970561695865, 32'sd0.021346903679223615, 32'sd0.050451661399224405, 32'sd-0.018347695143791094, 32'sd-0.0840822797713245, 32'sd-0.0369628796902968, 32'sd-0.09306735666467264, 32'sd-0.02614023371233177, 32'sd0.07545005740379869, 32'sd0.06020028486177278, 32'sd-0.003219156538006543, 32'sd-0.06198699762554786, 32'sd0.06819554015359978, 32'sd0.030363590909317395, 32'sd-0.023327885394602812, 32'sd0.238052677858473, 32'sd0.14576249429746874, 32'sd0.25862946818394417, 32'sd0.32868533684505274, 32'sd0.3056551112245316, 32'sd0.12581407842625375, 32'sd0.01317589288859308, 32'sd0.03768899570893078, 32'sd0.07672453780601661, 32'sd-0.044991541291602516, 32'sd0.006693430918200958, 32'sd-0.016819301505334044, 32'sd-0.18876513336386708, 32'sd-0.00623339365990107, 32'sd-0.020168904653442062, 32'sd0.023516553998203592, 32'sd0.020784566185567725, 32'sd0.04072139834178754, 32'sd-0.012382462920317095, 32'sd0.05785426514137394, 32'sd0.001954881572244423, 32'sd0.003478530420011754, 32'sd0.08281910846063298, 32'sd0.11435557576705681, 32'sd0.07159328619849195, 32'sd-0.010108495542374236, 32'sd0.041972987347580454, 32'sd-0.01367548729773796, 32'sd0.11139988721574869, 32'sd0.05362494157961989, 32'sd0.18080308932835396, 32'sd0.10127370401190133, 32'sd0.06802928085784422, 32'sd0.11917456409011927, 32'sd0.13846153189832133, 32'sd0.17434341748170534, 32'sd0.07481811444711167, 32'sd0.051602654234576203, 32'sd0.12487681132376278, 32'sd-0.05587175498746599, 32'sd-0.2893734076461048, 32'sd-0.12339449277370049, 32'sd-0.02804384161388449, 32'sd0.041203286441458375, 32'sd0.055923514551651614, 32'sd0.055677147728103296, 32'sd0.0125444720019918, 32'sd-0.013534567077375824, 32'sd0.06785238801511034, 32'sd0.04849398378381003, 32'sd0.060913740212621775, 32'sd0.0008593728780641536, 32'sd0.04290933242032683, 32'sd0.027833868384079793, 32'sd-0.09915051890296309, 32'sd-0.037034801078365494, 32'sd-0.14017135571170522, 32'sd-0.14329093665411283, 32'sd-0.00823495128635018, 32'sd0.08558784174925277, 32'sd-0.0533943163684135, 32'sd-0.007931013291076405, 32'sd0.04986463641984759, 32'sd0.13495865460976747, 32'sd0.05906635538391956, 32'sd0.05906782740646996, 32'sd0.14428453814069533, 32'sd-0.013846923648552055, 32'sd-0.08956268867569198, 32'sd0.006697341369855098, 32'sd-0.0313025785223708, 32'sd0.05432004510232408, 32'sd0.026877224466095195, 32'sd0.03904167457999209, 32'sd-0.10196605637281897, 32'sd-0.05330884992749417, 32'sd-0.08701092197920354, 32'sd0.06930435188574731, 32'sd0.014775316253896633, 32'sd0.027504106008132138, 32'sd-0.06250258354624065, 32'sd0.06067572025192506, 32'sd0.06950531819134585, 32'sd0.05210321678494775, 32'sd-0.00900090920758821, 32'sd-0.11050691018111648, 32'sd-0.17578165358707953, 32'sd-0.04462078637840881, 32'sd-0.06447487981118444, 32'sd0.10918991916526351, 32'sd0.07112434894972593, 32'sd0.0031074102482089795, 32'sd0.04446572439275408, 32'sd0.03645894077316198, 32'sd0.17030061268023008, 32'sd0.08037818445912945, 32'sd-0.0033982239425966476, 32'sd0.048518581849909856, 32'sd0.0205559905176386, 32'sd0.09340966125633116, 32'sd-0.07501048446465582, 32'sd-0.022096587462271593, 32'sd-0.14189193273348175, 32'sd-0.14032254565684585, 32'sd-0.10767192679430801, 32'sd0.006522489172103994, 32'sd-0.06153039547608966, 32'sd-0.02850456287897264, 32'sd-0.06549842765519602, 32'sd-0.006826531021173961, 32'sd-0.0726043791757197, 32'sd-0.055399384151855136, 32'sd-0.13957470500506497, 32'sd-0.2114749768159351, 32'sd-0.1130909326933623, 32'sd-0.03500316376924762, 32'sd-0.01285482778279199, 32'sd0.011750839860538891, 32'sd-0.010782458960834948, 32'sd0.06060641791885187, 32'sd0.005837290670361499, 32'sd-0.002728041472740801, 32'sd0.009156242129871244, 32'sd-0.02559971769753087, 32'sd-0.08069707698004842, 32'sd0.003564411101485976, 32'sd-0.013227342642247467, 32'sd0.009748139909133842, 32'sd-0.042766901024509765, 32'sd-0.1101473783829114, 32'sd-0.012727304719751954, 32'sd-0.020405164893704454, 32'sd-0.03315101694125965, 32'sd-0.0249826583887646, 32'sd-0.1496209521694162, 32'sd-0.1534448651723158, 32'sd-0.14037845956018466, 32'sd-0.08435989332752786, 32'sd-0.14599177373605632, 32'sd-0.15398821177463842, 32'sd-0.10064819628647927, 32'sd-0.1370056714668157, 32'sd-0.022205293608748258, 32'sd-0.06453583709522179, 32'sd0.0038426372608848895, 32'sd-0.06204784442333711, 32'sd0.08912437587964145, 32'sd0.07385985105622776, 32'sd0.15766773207350904, 32'sd-0.04754400305594708, 32'sd0.023220966078422237, 32'sd0.045510736748002246, 32'sd-0.08047825760138795, 32'sd-0.04929310359513904, 32'sd-0.06302087654814993, 32'sd2.168318359915932e-127, 32'sd0.04996793633724627, 32'sd0.014944764523572407, 32'sd0.06675345172637481, 32'sd-0.11241665858176252, 32'sd-0.017409190530618446, 32'sd0.08418546859139199, 32'sd-0.04758131134756351, 32'sd0.020330284478411807, 32'sd-0.061722397866916065, 32'sd-0.13384201545161142, 32'sd-0.07717410349940464, 32'sd-0.1604032666356235, 32'sd-0.1979775352668633, 32'sd0.009599071010435816, 32'sd-0.04491517370358393, 32'sd0.024911389989759378, 32'sd-0.034584392348779636, 32'sd0.0664991183893725, 32'sd0.005850198912376765, 32'sd-0.03227934025529516, 32'sd-0.01001038710214276, 32'sd0.03292790390621983, 32'sd-0.04672027970590638, 32'sd0.07000017203849648, 32'sd0.0521736590425244, 32'sd0.04578455978116438, 32'sd0.020438206984331537, 32'sd-0.030214028175985994, 32'sd0.020627280335589398, 32'sd-0.032696042204442444, 32'sd0.062201061189276305, 32'sd0.07689520398763708, 32'sd0.10120591199905687, 32'sd-0.06619478133956745, 32'sd-0.09218365058221123, 32'sd-0.027709521637827104, 32'sd-0.09848388244056756, 32'sd-0.012811110727919057, 32'sd-0.06212548110837123, 32'sd0.01064641448245806, 32'sd-0.07330153001698321, 32'sd0.00513458497955736, 32'sd0.08416033999900963, 32'sd0.05542754559625737, 32'sd0.07859439688136084, 32'sd0.027879159255858328, 32'sd0.004234468869300029, 32'sd0.003039599266908363, 32'sd-0.07480741172689186, 32'sd-0.10335420845479719, 32'sd-0.0063010795085758665, 32'sd0.017803883931653674, 32'sd-0.027766043472114577, 32'sd-0.022982386541531483, 32'sd-0.05073740555873555, 32'sd0.05551731596644111, 32'sd-0.004457544946815467, 32'sd-0.03139683505532578, 32'sd-0.0008134522696376088, 32'sd0.0067546712673711455, 32'sd0.049375188573116464, 32'sd-0.04066118246594654, 32'sd-0.04093213238114958, 32'sd-0.11087802641673059, 32'sd-0.03217516770982717, 32'sd-0.14258023324559047, 32'sd-0.04033231006748574, 32'sd-0.005741414574764575, 32'sd-0.041913341669236756, 32'sd0.05117773282105243, 32'sd0.01813042636258364, 32'sd-0.02017780729087864, 32'sd-0.031063550065971172, 32'sd-0.10286251605942026, 32'sd0.003140078145535594, 32'sd-0.1224937091310838, 32'sd-0.038105377818908305, 32'sd-0.07191607597686399, 32'sd0.036916743943207445, 32'sd0.06875036449694878, 32'sd0.004922667197689234, 32'sd-0.012957097461520127, 32'sd-0.014823282425522884, 32'sd3.8413128804289985e-119, 32'sd0.019718975295208618, 32'sd-0.0852162428899587, 32'sd0.08420538818833904, 32'sd0.08288184244912422, 32'sd0.03308823257594208, 32'sd0.0032891903342377343, 32'sd0.015996335186944818, 32'sd0.024071094856353583, 32'sd0.03015857786126302, 32'sd0.06022060280065678, 32'sd0.04870926106052068, 32'sd0.028637583488052874, 32'sd-0.047025011455936266, 32'sd0.00513256352531539, 32'sd-0.01996997457632623, 32'sd-0.012137122767002346, 32'sd0.034761362277816545, 32'sd-0.08739134328996254, 32'sd-0.009235285491182415, 32'sd-0.06468235329543015, 32'sd0.002925301904600948, 32'sd-0.05319318400645056, 32'sd0.032982916339994034, 32'sd0.095752215171576, 32'sd0.010394916081866696, 32'sd-0.01931216375528383, 32'sd0.041333340394008385, 32'sd0.06748331730119193, 32'sd-0.0005756436049966811, 32'sd0.0797849244868397, 32'sd-0.07470894608942001, 32'sd-0.03742602139143781, 32'sd-0.014008177754000161, 32'sd0.09307193211989795, 32'sd0.0228315394655904, 32'sd0.07104344101949164, 32'sd0.02097636231510379, 32'sd0.06955463779041444, 32'sd0.03287433858965178, 32'sd0.03506934447683871, 32'sd-0.05516373660285118, 32'sd0.05390687636934014, 32'sd0.05240077705166826, 32'sd-0.09747916735392632, 32'sd0.010318648162928578, 32'sd-0.021577484551032148, 32'sd-0.08257053767186344, 32'sd0.06179984787213135, 32'sd0.09439668547353747, 32'sd-0.053973594406211786, 32'sd0.008171297500212041, 32'sd0.09883210316290933, 32'sd0.03884998942668375, 32'sd0.015582636753093418, 32'sd0.034713221767968726, 32'sd0.11524039083601212, 32'sd0.08320920337811621, 32'sd0.023981440740363576, 32'sd0.022258829262592365, 32'sd0.02359403851170643, 32'sd-0.11313160008881105, 32'sd-0.06641727186340497, 32'sd-0.010249976311395183, 32'sd0.061144292078107704, 32'sd0.07191653862556491, 32'sd0.12573669422747027, 32'sd0.03602896048157391, 32'sd0.06170594664695515, 32'sd0.0137614302043273, 32'sd0.06074699987670697, 32'sd0.021755762613405817, 32'sd-0.00834450943423199, 32'sd-0.027042043629012875, 32'sd-0.03495486846864575, 32'sd-0.13985150037020994, 32'sd-0.04442237273872595, 32'sd-0.02981713142989836, 32'sd0.02994443703382221, 32'sd0.11106353434465548, 32'sd0.04440692386923721, 32'sd0.014680133338030426, 32'sd0.01905417307644985, 32'sd0.030214189909080792, 32'sd5.483224967765635e-125, 32'sd-0.0041972658825023415, 32'sd-0.019587204765259013, 32'sd-0.024640754496661133, 32'sd0.02784492284989413, 32'sd0.07148738122499919, 32'sd-0.08785588737823709, 32'sd0.005946129779977168, 32'sd0.13155513472601188, 32'sd0.10609662202337458, 32'sd0.014110160017523188, 32'sd0.016114116970365164, 32'sd0.019831090024827306, 32'sd0.06490939886141547, 32'sd0.0008240950810135482, 32'sd0.01537259033160235, 32'sd-0.00708345932409552, 32'sd0.026113883387146035, 32'sd0.001857491911814357, 32'sd-0.05324051412714026, 32'sd0.0830681754139914, 32'sd-0.02540569636455127, 32'sd0.0288101885377538, 32'sd0.007302131051038568, 32'sd0.05642850038440631, 32'sd-0.009231020541855685, 32'sd0.006713754534601341, 32'sd1.2424887366088065e-119, 32'sd-2.1705844693574493e-127, 32'sd-5.092155840899708e-128, 32'sd-0.05832231355860186, 32'sd0.03219503807480334, 32'sd-0.0578371837047274, 32'sd0.040817181225951266, 32'sd0.028939548681983444, 32'sd0.09381671878826355, 32'sd0.18043765106974374, 32'sd0.06389023312106333, 32'sd0.1250649614516596, 32'sd0.014041101337494562, 32'sd-0.07884197191760751, 32'sd-0.15605118419282243, 32'sd-0.10162487982913077, 32'sd0.02294963815048664, 32'sd0.10064224828210794, 32'sd-0.0018862436201243084, 32'sd-0.05039811214187117, 32'sd0.0617181073294601, 32'sd-0.007798954808132957, 32'sd0.007305818854459687, 32'sd-0.05295744189131359, 32'sd0.04422230855807431, 32'sd0.0724789538085959, 32'sd-0.0552288104364386, 32'sd-0.07947324732273926, 32'sd3.704009044888068e-122, 32'sd5.8454748983164453e-126, 32'sd3.257303026695523e-120, 32'sd0.03793104921140834, 32'sd0.05802340844339805, 32'sd-0.08733945458116761, 32'sd-0.028873546920643266, 32'sd0.16093139298959205, 32'sd0.08601455067818381, 32'sd0.07681549631089128, 32'sd0.1182416391271627, 32'sd0.0034042542130703554, 32'sd0.02530454371427909, 32'sd0.0899594440574459, 32'sd-0.029857372969789908, 32'sd0.035418421178500886, 32'sd0.16254901399269503, 32'sd0.17353829765839215, 32'sd-0.03210442353525767, 32'sd-0.093604976856507, 32'sd0.10867144857703355, 32'sd-0.05195736818622815, 32'sd-0.06626686348219257, 32'sd-0.14871817757306965, 32'sd-0.05094464362426459, 32'sd-0.12070812890522159, 32'sd0.04842247477287512, 32'sd0.017941694469683, 32'sd-4.407841213226942e-123, 32'sd-7.289883020179721e-115, 32'sd3.6279280585723162e-127, 32'sd-9.897268550151934e-122, 32'sd0.09224681719890246, 32'sd-0.020179563773501292, 32'sd0.05602430049622017, 32'sd0.002342537386324631, 32'sd0.03881532762078993, 32'sd-0.04214752333715126, 32'sd-0.08498229448766152, 32'sd0.010459761791789798, 32'sd0.07990756562579206, 32'sd0.030752252694684238, 32'sd0.055157786968385636, 32'sd0.10614838438419352, 32'sd0.05985667087503883, 32'sd0.014266347307320404, 32'sd0.05658418206567116, 32'sd-0.021502707513456214, 32'sd-0.01488523156855688, 32'sd0.008937000636525336, 32'sd-0.08540919942893375, 32'sd-0.0033515051490272756, 32'sd-0.01354031777433618, 32'sd0.019844952737531334, 32'sd-0.0044016840969210574, 32'sd2.895228995406996e-116, 32'sd5.251566415158716e-120, 32'sd-7.112717783693987e-117, 32'sd-1.2877234837478977e-122, 32'sd2.4044727758534566e-125, 32'sd-5.000256871547999e-117, 32'sd0.015782722128184542, 32'sd-0.05289214612220204, 32'sd0.09086993503414108, 32'sd0.08234949718275815, 32'sd0.06135398316940037, 32'sd0.05736702070407493, 32'sd-0.01456213474612158, 32'sd-0.037646648000337984, 32'sd-0.00301920927433417, 32'sd-0.01622979765131497, 32'sd0.07709004568487053, 32'sd0.020491612436522748, 32'sd-0.06351217832670923, 32'sd0.0795746958820386, 32'sd-0.08272629778488266, 32'sd-0.07249171260641867, 32'sd0.042014115946202454, 32'sd-0.019040112867168366, 32'sd0.008779341817378931, 32'sd0.031109894188776074, 32'sd4.776557682539499e-121, 32'sd3.43404684796205e-116, 32'sd-3.3446255183742814e-116, 32'sd-1.1394794800817427e-119},
        '{32'sd8.748008223739207e-124, 32'sd-2.8079360326332937e-117, 32'sd1.9210605468125362e-121, 32'sd-7.05312464953414e-120, 32'sd1.7584034475737835e-123, 32'sd-9.878644655590028e-120, 32'sd-2.1707914498915982e-127, 32'sd6.260992677664203e-123, 32'sd3.7873529685293836e-125, 32'sd1.829691392330581e-116, 32'sd3.8315149060685714e-125, 32'sd6.264888384150886e-126, 32'sd-0.011744328742805718, 32'sd-0.0703799970465918, 32'sd0.03164310269958952, 32'sd0.005682725685513417, 32'sd-6.160168571956839e-120, 32'sd1.0833876868834525e-115, 32'sd-7.199823569130936e-116, 32'sd4.7845130424845405e-124, 32'sd-6.473674455214453e-124, 32'sd3.6200949798601746e-116, 32'sd-6.325547253663619e-125, 32'sd1.488196418468401e-123, 32'sd-1.5135860069146044e-115, 32'sd1.0585478741899681e-119, 32'sd5.763349404138356e-119, 32'sd-1.3725847976845743e-117, 32'sd-1.036758109811673e-120, 32'sd1.0137662473957157e-124, 32'sd-1.6792009568607872e-120, 32'sd-1.8447687496662145e-118, 32'sd-0.020400779495143073, 32'sd-0.05191224274187703, 32'sd-0.030699127176718514, 32'sd-0.054983930444465354, 32'sd-0.034575395114638224, 32'sd-0.07783848942949569, 32'sd-0.06462275831040616, 32'sd-0.046401712042245476, 32'sd-0.05807254455951472, 32'sd0.03493694125269363, 32'sd-0.0591195599428587, 32'sd-0.0853511264692117, 32'sd-0.06495830426566182, 32'sd-0.08817431680077777, 32'sd-0.006303053735371768, 32'sd-0.03548156892690289, 32'sd0.06577279579013671, 32'sd0.003967684691028534, 32'sd-0.06002062100611767, 32'sd0.022774059645940568, 32'sd-2.817725830497902e-123, 32'sd1.4935176676662318e-125, 32'sd4.749752882870109e-126, 32'sd5.308353840865636e-130, 32'sd7.766717614218622e-122, 32'sd1.0311774180015847e-122, 32'sd-0.05002016329245407, 32'sd-0.00562695343767513, 32'sd-0.045662191991823545, 32'sd-0.063460254474897, 32'sd0.02222117440944168, 32'sd-0.017396810622625717, 32'sd-0.058749850477027785, 32'sd0.03887718427629602, 32'sd-0.03370739139312868, 32'sd-0.1751514465741297, 32'sd0.12914539011329126, 32'sd0.03329233850461232, 32'sd-0.03616619690154473, 32'sd-0.08135430104304855, 32'sd-0.01170956949590198, 32'sd-0.013405163796392922, 32'sd0.02900732506585938, 32'sd-0.0884324386515004, 32'sd-0.009338178222609893, 32'sd-0.07013063474206123, 32'sd-0.08677895585893738, 32'sd-0.04493517343061816, 32'sd-0.01279121122217239, 32'sd-0.05189124790219894, 32'sd-7.564843011466903e-115, 32'sd-1.5475572126969563e-115, 32'sd1.0013595385052045e-120, 32'sd-7.993048773460486e-115, 32'sd0.010297992825294755, 32'sd-0.027326927197492152, 32'sd-0.05094137105960801, 32'sd-0.03852126473613429, 32'sd0.059119463183233356, 32'sd-0.054347168142084186, 32'sd-0.08479369932201239, 32'sd-0.055329945543494734, 32'sd-0.03448739146384227, 32'sd-0.1404006141508856, 32'sd-0.12089906606383317, 32'sd-0.12321421618464405, 32'sd-0.06941712417834599, 32'sd-0.02162157424917463, 32'sd-0.02351556019380223, 32'sd-0.09700098976831555, 32'sd0.024055300484411037, 32'sd-0.0367624675127251, 32'sd0.048709473999036156, 32'sd0.04171442095171707, 32'sd-0.05518849338057749, 32'sd-0.008691063207662367, 32'sd-0.02119215914056907, 32'sd0.011295522295344187, 32'sd-0.023817064922308628, 32'sd-8.851540248987952e-127, 32'sd-6.807934703738958e-128, 32'sd-0.02274031371389962, 32'sd-0.0330277754526587, 32'sd-0.054872984429469245, 32'sd-0.04742748159737397, 32'sd0.027910702860560476, 32'sd-0.001322246799983232, 32'sd0.016721015508602926, 32'sd-0.10309480315241802, 32'sd-0.12558098031306, 32'sd-0.10942921530561268, 32'sd-0.13355696480523832, 32'sd-0.02193070777538875, 32'sd-0.15752892502981486, 32'sd-0.11123571360042239, 32'sd-0.22863873079333633, 32'sd-0.21379617148613025, 32'sd-0.07802358334100709, 32'sd-0.04523587858546595, 32'sd-0.022780491469242548, 32'sd0.062310721878505664, 32'sd0.11703379320094076, 32'sd0.0679823915541807, 32'sd-0.033500590586741014, 32'sd-0.014282886506402817, 32'sd-0.06346955960748885, 32'sd-0.08210013415034194, 32'sd0.08317354710477874, 32'sd-2.129537740437681e-124, 32'sd0.00960086203213532, 32'sd-0.06122502738858546, 32'sd-0.07222940524407095, 32'sd-0.1330957082918713, 32'sd0.010063692275226346, 32'sd0.022484181566221915, 32'sd0.08151278001334918, 32'sd0.133223912574772, 32'sd-0.018982617684182985, 32'sd0.09229834975272179, 32'sd0.020876001595657837, 32'sd0.13441155727535614, 32'sd-0.004777588378001599, 32'sd-0.030485444500699198, 32'sd0.008400296797623177, 32'sd-0.04934791542216597, 32'sd0.08157928989115272, 32'sd-0.14274966299900413, 32'sd-0.22619838447556945, 32'sd-0.06198174078606969, 32'sd0.12537017854961727, 32'sd0.15029923936082848, 32'sd-0.028723213077201562, 32'sd-0.0765599348511117, 32'sd-0.09075311169449668, 32'sd0.04128416438473628, 32'sd0.029788243581753273, 32'sd2.3964013179203108e-124, 32'sd-0.049782014412208746, 32'sd0.016887140463369126, 32'sd0.05184531853985717, 32'sd0.02903830266652283, 32'sd-0.00825423662323967, 32'sd-0.06156685142134353, 32'sd0.07830422031986185, 32'sd0.01752573357249246, 32'sd0.07242433032061074, 32'sd0.15286234675475457, 32'sd0.0763903983971907, 32'sd0.06643918400747438, 32'sd0.09738641732293807, 32'sd-0.015087274126227826, 32'sd-0.02821197967209466, 32'sd0.1258823834462471, 32'sd0.1542288018397528, 32'sd0.03253462282349489, 32'sd-0.09534162944167099, 32'sd-0.029686210188640556, 32'sd0.09665225621780207, 32'sd0.16351965448167013, 32'sd0.14086454857879127, 32'sd0.045643497259768184, 32'sd0.06327008730407498, 32'sd0.06886262945167317, 32'sd-0.14434594027907627, 32'sd0.012134969907594656, 32'sd-0.03421395313852324, 32'sd0.09792904112935544, 32'sd-0.010682670659525466, 32'sd-0.07887164735816844, 32'sd-0.18657554054193332, 32'sd-0.10431745834450529, 32'sd0.028457758279277143, 32'sd-0.04042194267592685, 32'sd0.002233289811688152, 32'sd0.026285105001032393, 32'sd0.1515267992522011, 32'sd0.10335019400050864, 32'sd0.08012499372256922, 32'sd-0.08027426912532937, 32'sd-0.17231855504947052, 32'sd-0.001413757374829378, 32'sd0.022812916549724203, 32'sd0.0028520019298203885, 32'sd-0.08246988984472688, 32'sd-0.026396724969917615, 32'sd0.10134530282685837, 32'sd0.10280640069678704, 32'sd0.1181415295805715, 32'sd0.058496666213358285, 32'sd-0.10952999883124469, 32'sd0.03455280543060083, 32'sd-0.0598402260727281, 32'sd-0.05253645015569425, 32'sd-0.04038402278053454, 32'sd0.0865535749342022, 32'sd0.008998450608365955, 32'sd0.005641582289239153, 32'sd-0.01765201299619883, 32'sd0.02859941832432917, 32'sd-0.021921613484530138, 32'sd0.08551313072323406, 32'sd0.003534711113575489, 32'sd0.0637175749836128, 32'sd0.14600384825996032, 32'sd0.14556252920220009, 32'sd-0.10425065932483832, 32'sd-0.08702450432490257, 32'sd-0.0468872340257712, 32'sd-0.016750611132236255, 32'sd-0.05093198855212485, 32'sd-0.001389017539135778, 32'sd-0.005800611804372319, 32'sd0.06126012598064938, 32'sd0.03106928131558628, 32'sd0.07649358357594215, 32'sd0.1483939037338227, 32'sd-0.029202993327457984, 32'sd-0.0793431099614492, 32'sd-0.13486172255391599, 32'sd0.012522314943074401, 32'sd0.06675607223368185, 32'sd0.09292127823076199, 32'sd-0.04550045809270106, 32'sd0.0503141946589362, 32'sd0.11358131996543272, 32'sd-0.03473628029386177, 32'sd0.03586770751194704, 32'sd0.0509987095022515, 32'sd-0.01519863047998484, 32'sd0.04792244894076006, 32'sd0.05258429286931265, 32'sd0.06519939743878062, 32'sd0.1397931323316711, 32'sd-0.055343328298030306, 32'sd-0.051651373787926926, 32'sd-0.12091338345090118, 32'sd-0.08542083768959392, 32'sd0.04583757543752195, 32'sd0.07242834348539547, 32'sd0.05799372414150725, 32'sd0.13395950887019736, 32'sd0.03785007841779704, 32'sd-0.02892302264379315, 32'sd0.005000756121521103, 32'sd-0.03984992743065581, 32'sd0.02516822877042611, 32'sd0.013539845615398808, 32'sd0.026172447108197914, 32'sd-0.03470487075692981, 32'sd0.02675669506476539, 32'sd0.019145834921375313, 32'sd-0.00363722478092153, 32'sd0.15552929125191597, 32'sd0.014617859513997711, 32'sd0.0014993647445010777, 32'sd-0.06616435789924231, 32'sd0.06693633640945156, 32'sd0.08529153000538825, 32'sd0.07052019402243953, 32'sd0.16584806330333698, 32'sd-0.016329701646604782, 32'sd0.0532767059487347, 32'sd-0.03245626187712762, 32'sd0.013361093749766333, 32'sd0.017478801444969848, 32'sd-0.04776808388220477, 32'sd0.0961529161110454, 32'sd0.07820894107245546, 32'sd0.04885612830681787, 32'sd0.036758520082751336, 32'sd0.06898380809310573, 32'sd0.03006500064847785, 32'sd0.015945042165708346, 32'sd0.0979661320952071, 32'sd0.043616019309132545, 32'sd0.026946709343972246, 32'sd-0.038942726765985584, 32'sd-0.011533371913300327, 32'sd0.07863797061139888, 32'sd0.05553008121201335, 32'sd0.05507099576431989, 32'sd0.04544371528187983, 32'sd-0.013032321019496203, 32'sd0.1666108092987173, 32'sd0.21331469044985993, 32'sd0.09650929151964979, 32'sd0.03540132217738647, 32'sd0.16086305962069652, 32'sd0.2035188262150177, 32'sd0.0581747207162883, 32'sd0.0006704524330484348, 32'sd0.17530392849990498, 32'sd0.022099696217845112, 32'sd-0.01230180594495175, 32'sd-0.030769670701784, 32'sd0.09493164806051697, 32'sd0.14757128510452533, 32'sd0.07858034094042547, 32'sd-0.02457910876579094, 32'sd-0.009946381159945292, 32'sd0.012542376765152657, 32'sd0.0022264210989787407, 32'sd0.05554354082529615, 32'sd0.04582687331307202, 32'sd0.002389840565032536, 32'sd0.02474217195829703, 32'sd-0.009687221776836338, 32'sd-0.04480099622717455, 32'sd-0.03593493751684573, 32'sd-0.05636417965383627, 32'sd-0.07711065318629517, 32'sd0.15623496291091188, 32'sd0.1365647851007088, 32'sd0.03463186821558425, 32'sd0.16839238283414615, 32'sd0.16034328191722585, 32'sd0.11629845478282962, 32'sd0.08699287426213237, 32'sd-0.1240555817258376, 32'sd0.07766797753727897, 32'sd-0.06005903749103513, 32'sd-0.03294193549219383, 32'sd0.009843012088687717, 32'sd-0.013163085012826323, 32'sd-0.050065617747742285, 32'sd0.008493108150796881, 32'sd-0.012912459050023382, 32'sd-0.0630835186509442, 32'sd-0.008084983454767486, 32'sd0.001294069663999453, 32'sd-0.0725436589519243, 32'sd-0.0830175743237698, 32'sd-0.038008270893661364, 32'sd-0.06255839253769467, 32'sd-0.04004691706759884, 32'sd0.006209388882290046, 32'sd-0.018053055463410964, 32'sd-0.0031942352941138, 32'sd0.12406831619377294, 32'sd0.14443128348450238, 32'sd0.03158250866581553, 32'sd-0.03419142824114664, 32'sd-0.09394230889418272, 32'sd-0.058150389997109524, 32'sd-0.029132432774425933, 32'sd-0.01342050201638821, 32'sd-0.12348392370100968, 32'sd0.05769485377136076, 32'sd-0.04593168718584724, 32'sd-0.06503352082955663, 32'sd0.041846188850046984, 32'sd-0.0363748439299924, 32'sd-0.1259077801531241, 32'sd-0.030045018616713434, 32'sd-0.07370061176190665, 32'sd0.0005303560656985413, 32'sd0.1579688885384883, 32'sd0.10808864192977807, 32'sd0.04563386754966446, 32'sd-0.04067805910771588, 32'sd-0.05438678211408918, 32'sd0.015894892559495624, 32'sd-0.046641366905739265, 32'sd0.011940900740925752, 32'sd0.09711576791735904, 32'sd0.017040912708452968, 32'sd0.11968432141413551, 32'sd0.0759036679050619, 32'sd0.08215424309708105, 32'sd0.01640957580151992, 32'sd-0.08331377029237612, 32'sd-0.11130423624341768, 32'sd0.06935823934944309, 32'sd-0.050592521023937166, 32'sd-0.1174275842796826, 32'sd-0.05381077215263116, 32'sd-0.1583182825061434, 32'sd0.03613613032278617, 32'sd-0.015919960130774197, 32'sd0.002815205180479902, 32'sd-0.13295999133840516, 32'sd-0.1169516110842689, 32'sd-0.07042374338957127, 32'sd-0.08765149992783265, 32'sd0.0005070119617221475, 32'sd0.01687134043643013, 32'sd-0.12143515681649288, 32'sd0.018482507349679995, 32'sd0.056034932362389024, 32'sd0.004013892504129525, 32'sd-0.1038374626703594, 32'sd-0.04701281592871866, 32'sd-0.006913972633475034, 32'sd-0.0245504151724294, 32'sd0.09996397871555493, 32'sd0.05472509045192093, 32'sd-0.06551728562783564, 32'sd-0.0988174902158186, 32'sd0.01503596574197761, 32'sd-0.1130311930823872, 32'sd-0.1295414423425082, 32'sd-0.11873572974555313, 32'sd-0.07965600934136774, 32'sd0.07360538918496502, 32'sd-0.0953925975908852, 32'sd-0.07373742538358699, 32'sd-0.02583703366059227, 32'sd0.01323369242235245, 32'sd-0.09462171495767946, 32'sd-0.01355335338882577, 32'sd-0.01493976421450183, 32'sd-0.0452942025147671, 32'sd-0.04548919254076315, 32'sd-0.04884396946920324, 32'sd0.005415573573474129, 32'sd0.05236555812147857, 32'sd0.011740626112953744, 32'sd-0.03749161991212064, 32'sd-0.06922898710554914, 32'sd-0.09484726373018935, 32'sd-0.045607966807749464, 32'sd0.0015006692923603996, 32'sd-0.09566719881367185, 32'sd-0.048026921460653904, 32'sd0.044577075095431344, 32'sd-0.13590941795459172, 32'sd-0.010697613477694481, 32'sd-0.16477638946297293, 32'sd-0.14126501333491076, 32'sd-0.0817391090741185, 32'sd0.009940027394074583, 32'sd0.08704967428729177, 32'sd-0.015353618463988056, 32'sd0.058103689439880105, 32'sd-0.0003047900438992875, 32'sd-0.017205686369029843, 32'sd-0.06055358841932417, 32'sd0.02659380130336039, 32'sd0.09296505386200721, 32'sd0.07208340543145536, 32'sd-0.019594435336867364, 32'sd0.069345091702421, 32'sd-0.006987706745149889, 32'sd-0.03690840479783401, 32'sd1.9659877653041425e-127, 32'sd-0.004548092206938254, 32'sd0.0028720736641489088, 32'sd-0.1337495495416301, 32'sd-0.09788098383596887, 32'sd-0.10616670639437874, 32'sd-0.1393274387544227, 32'sd-0.08077790214315415, 32'sd-0.01281494652534764, 32'sd-0.10928288035078484, 32'sd-0.0052610057147514655, 32'sd-0.0488991160779302, 32'sd-0.1516099699363095, 32'sd-0.07156151862219202, 32'sd-0.1284609435008227, 32'sd0.04091926087990493, 32'sd-0.030315551938760645, 32'sd-0.03273017552415684, 32'sd-0.033817295265942196, 32'sd-0.08420615097432844, 32'sd0.021690266126236386, 32'sd0.09535927321657697, 32'sd0.05588947360671833, 32'sd-0.04719929511477025, 32'sd0.02497465444897638, 32'sd0.057012554903180586, 32'sd0.10106624835852682, 32'sd-0.003116179889015833, 32'sd-0.04392030062426682, 32'sd-0.009136780294727954, 32'sd0.00873617206486116, 32'sd0.036115246118236376, 32'sd0.009179884581936368, 32'sd-0.20780096775339693, 32'sd-0.12862209720410775, 32'sd-0.15587733032528256, 32'sd-0.06577823375962065, 32'sd-0.15167719252664374, 32'sd-0.006677589174839448, 32'sd-0.16062038579827917, 32'sd-0.06669623091071665, 32'sd0.06740768931848226, 32'sd0.002828495870468813, 32'sd0.02156856372619118, 32'sd-0.00106825066687806, 32'sd-0.06300152045637711, 32'sd-0.13431002688285523, 32'sd-0.15893671586417177, 32'sd-0.04616291296256732, 32'sd0.07595277795394506, 32'sd0.03731877688889809, 32'sd-0.026180584709213445, 32'sd-0.14182395224716243, 32'sd-0.12913410846420145, 32'sd-0.02198661008306447, 32'sd-0.045709110272548634, 32'sd-0.04810185108759253, 32'sd0.007916162039753104, 32'sd0.03872078665601812, 32'sd-0.07328256444007894, 32'sd0.028493236001781632, 32'sd-0.11745415904742672, 32'sd-0.1405812322676576, 32'sd-0.196520383495347, 32'sd-0.11160194280538402, 32'sd-0.09963459527766944, 32'sd-0.16904275458137608, 32'sd-0.1736761824221448, 32'sd0.11475471241061207, 32'sd0.06284611111896551, 32'sd0.09125569434802142, 32'sd-0.05759722693905584, 32'sd-0.10794340686191299, 32'sd-0.11877918592776135, 32'sd-0.13851789228563807, 32'sd-0.20452738689854946, 32'sd-0.11815105934863339, 32'sd-0.0015626481270130993, 32'sd0.0010032515856840763, 32'sd0.0781059122096948, 32'sd-0.07934595314892554, 32'sd-0.06313099400978989, 32'sd0.059589992210897204, 32'sd-0.08718386677450465, 32'sd2.967406665203171e-119, 32'sd0.02458268936811627, 32'sd0.028433942011546656, 32'sd-0.06756085726872431, 32'sd-0.14730592574803106, 32'sd-0.1752539815535723, 32'sd-0.17425191554424532, 32'sd-0.10661427376256885, 32'sd0.0014831421622672207, 32'sd0.05159753385100606, 32'sd-0.10630888045321839, 32'sd0.007603567261446141, 32'sd0.1398765939514584, 32'sd0.057438527297982434, 32'sd-0.08793506723785918, 32'sd-0.14400465539601734, 32'sd-0.17291243538716924, 32'sd-0.16200638698587905, 32'sd-0.14663674232084928, 32'sd-0.11282495974803178, 32'sd-0.045001804390139954, 32'sd-0.026323600350267293, 32'sd-0.06718262985616713, 32'sd0.07346801897258294, 32'sd-0.03925855924578085, 32'sd-0.009424029074720163, 32'sd0.000787551619609148, 32'sd-0.007830875619409686, 32'sd7.227922565328556e-05, 32'sd-0.014632825939830871, 32'sd-0.06886411751393143, 32'sd-0.1202671473651993, 32'sd-0.030484031716352934, 32'sd-0.13181077316551637, 32'sd-0.0795895122933064, 32'sd-0.12714778603105675, 32'sd-0.03669601527119172, 32'sd-0.06324451946226485, 32'sd-0.10819061771603167, 32'sd0.015510086381530275, 32'sd0.06628380802899422, 32'sd-0.0364140793511822, 32'sd-0.036034974493698156, 32'sd-0.07354995891589565, 32'sd-0.04420380563702615, 32'sd-0.07383879195856458, 32'sd-0.16439426673256943, 32'sd-0.12003738541146461, 32'sd0.023959820758710688, 32'sd0.11333696659942269, 32'sd0.08754871995411058, 32'sd0.0033973574601132445, 32'sd0.003934769594951661, 32'sd-0.009247409644874936, 32'sd-0.045712867061708864, 32'sd-0.016946848404335208, 32'sd-0.007619773833977713, 32'sd-0.13484780866089952, 32'sd0.06659618910636696, 32'sd-0.05506690131138344, 32'sd-0.025941483679790493, 32'sd-0.147536062388333, 32'sd0.014177935227498257, 32'sd0.07901904727934433, 32'sd-0.07219937689432261, 32'sd0.0023242931170164216, 32'sd0.06764341263781713, 32'sd-0.010028941548438065, 32'sd-0.008765019792845946, 32'sd-0.02362640568560287, 32'sd-0.049293923310791216, 32'sd-0.005383099326134235, 32'sd-0.11508254254322987, 32'sd-0.0946388900415177, 32'sd-0.09712540277815201, 32'sd-0.1244964043683929, 32'sd0.0033052791829176016, 32'sd0.005137524585213167, 32'sd-0.10158343262538472, 32'sd-0.04170508017229814, 32'sd-0.04093838509407448, 32'sd0.007322767098311248, 32'sd-0.05301201819942226, 32'sd-0.009129191413213477, 32'sd-6.9221661661415705e-124, 32'sd-0.01991447149204545, 32'sd0.05662703626049178, 32'sd0.105167490476695, 32'sd0.0957031173634162, 32'sd-0.10775533481797608, 32'sd0.08402601203660055, 32'sd0.09123535693454989, 32'sd0.07237835000891117, 32'sd0.07233848730339767, 32'sd-0.07760121203937917, 32'sd0.07733530568728494, 32'sd-0.013207886502041206, 32'sd-0.025789154143385062, 32'sd0.04325109477564805, 32'sd-0.09201502553457638, 32'sd0.006503654217918332, 32'sd-0.055668950221750606, 32'sd-0.18596650785030677, 32'sd-0.21958545006701422, 32'sd-0.013130189896251036, 32'sd0.06920481414050231, 32'sd-0.04150192602714028, 32'sd-0.07313014051419206, 32'sd-0.08671783948529083, 32'sd0.03948367488236692, 32'sd-0.019288757753897563, 32'sd-3.1502811625502007e-115, 32'sd2.3379530323899034e-114, 32'sd1.2705248289765665e-123, 32'sd-0.08261190023852587, 32'sd-0.032159108738879234, 32'sd-0.06929825568534603, 32'sd-0.0669189232118872, 32'sd0.012808337891594353, 32'sd-0.011705775240909962, 32'sd0.08900654375950519, 32'sd-0.04124579060296086, 32'sd0.08234743071963445, 32'sd0.13725477551270707, 32'sd-0.03960419383977788, 32'sd0.07114589024828319, 32'sd0.041024434080648715, 32'sd0.09681249515691773, 32'sd-0.02574030873791403, 32'sd0.016558407314610356, 32'sd-0.08879727237947103, 32'sd-0.22980893721966128, 32'sd-0.07057511110994542, 32'sd-0.0875494543111285, 32'sd0.13066547747792004, 32'sd-0.003016869849015159, 32'sd0.028756049272748874, 32'sd-0.02836902117722268, 32'sd-0.021474009116415577, 32'sd-3.8194745687017823e-119, 32'sd6.894317811143145e-120, 32'sd9.143337964666186e-122, 32'sd-0.044909896252016517, 32'sd0.04069733524018705, 32'sd0.016584534581565984, 32'sd0.006120690095755119, 32'sd-0.06505790418573573, 32'sd0.07621095584891198, 32'sd-0.021367359614455537, 32'sd0.010747478951718115, 32'sd-0.0053710640722325394, 32'sd-0.030662433414792627, 32'sd-0.08558636063915842, 32'sd-0.044748127816055465, 32'sd0.037929282975120666, 32'sd0.018691168507194288, 32'sd0.055685963162963925, 32'sd0.042999147578938336, 32'sd-0.05624542266557761, 32'sd-0.1870130351340089, 32'sd-0.14622896283096395, 32'sd-0.09449804286558887, 32'sd0.05871562102973682, 32'sd-0.0012655429516770702, 32'sd-0.02308131427484717, 32'sd-0.04620590801860652, 32'sd-0.039608314823574325, 32'sd-1.035961251038214e-122, 32'sd-3.6449850116871125e-116, 32'sd1.7242422996844246e-124, 32'sd3.676541562985067e-116, 32'sd0.0037066373344124214, 32'sd-0.054270363072331546, 32'sd-0.06341353364248986, 32'sd0.00534927570788701, 32'sd-0.08741920790739732, 32'sd0.07607314821326037, 32'sd-0.00926589892883979, 32'sd0.07880864463379865, 32'sd-0.028287811964686473, 32'sd0.03644810831926061, 32'sd0.06246708489198457, 32'sd0.021684884005439498, 32'sd-0.12171265074005129, 32'sd-0.03587640855336909, 32'sd0.11998736404303803, 32'sd0.05943850122960139, 32'sd-0.07048264645875012, 32'sd0.06034574343354767, 32'sd0.014567939619801783, 32'sd0.030021282688291875, 32'sd0.03836023028362496, 32'sd-0.12522789193756365, 32'sd0.05029998913254073, 32'sd1.5397942779680282e-115, 32'sd-8.850805980494868e-125, 32'sd-8.474730425524649e-119, 32'sd-1.7786959267339968e-122, 32'sd-1.10992906257638e-121, 32'sd1.2714388297104875e-118, 32'sd-0.0415268175078861, 32'sd-0.030512615098299303, 32'sd0.009929728878382811, 32'sd0.015065865973139058, 32'sd-0.05121794019247089, 32'sd0.047690182405807094, 32'sd-0.027409363764362118, 32'sd-0.05874678067548809, 32'sd0.010263612484085765, 32'sd-0.07988599122473947, 32'sd0.07069614677177809, 32'sd-0.001365951311027112, 32'sd0.008633642195107922, 32'sd0.107021563665267, 32'sd0.015737960943044693, 32'sd-0.03569008579941381, 32'sd-0.043039459971543736, 32'sd0.012832059863559264, 32'sd0.07626102403744855, 32'sd0.09545263585226765, 32'sd-7.400773831241279e-120, 32'sd6.886134445184346e-126, 32'sd-2.0453238084816413e-126, 32'sd3.688974092996422e-122},
        '{32'sd-2.1456737599943905e-127, 32'sd2.55213963328791e-116, 32'sd-2.0534842604460585e-117, 32'sd-4.816947534776885e-125, 32'sd4.663821934811415e-124, 32'sd3.6313959407396705e-126, 32'sd-5.2735455774301015e-118, 32'sd-8.38975096046311e-117, 32'sd-8.339629486752964e-116, 32'sd-8.51755213306088e-119, 32'sd7.561585389635008e-115, 32'sd9.707847978059516e-125, 32'sd0.08100933007451094, 32'sd0.09281021876371245, 32'sd-0.019735485223744693, 32'sd-0.0017843526178701627, 32'sd-2.6930212738619976e-124, 32'sd1.1517352183055476e-119, 32'sd-4.577867635397192e-118, 32'sd5.940310354509888e-124, 32'sd2.5605690905695212e-117, 32'sd3.6902834256918506e-118, 32'sd-1.0127008857919451e-124, 32'sd5.0614314431137335e-115, 32'sd-8.914799483609868e-123, 32'sd3.8744913096884876e-125, 32'sd2.1623561170300724e-116, 32'sd-3.1837510721238244e-125, 32'sd-4.520393631520032e-123, 32'sd1.0863526230024448e-118, 32'sd1.2111053777214646e-125, 32'sd2.1285111559487245e-120, 32'sd-0.02005432212202672, 32'sd0.0005478983450561729, 32'sd-0.010046639437016803, 32'sd0.02716837407688283, 32'sd0.014461912231460977, 32'sd-0.0051453013576492415, 32'sd-0.026723245376659405, 32'sd0.1090687020935724, 32'sd-0.02093162277370378, 32'sd-0.03605403960933961, 32'sd0.04311731840334342, 32'sd-0.07415646500881534, 32'sd-0.11240178444863572, 32'sd0.0015719542438699546, 32'sd-0.04018311822873689, 32'sd0.02960926853614165, 32'sd0.0008487666178636331, 32'sd-0.003285538799302869, 32'sd-0.017447653030920524, 32'sd-0.0023024352873985865, 32'sd4.9373126090236935e-124, 32'sd-2.825467905571447e-119, 32'sd-5.267865533036402e-124, 32'sd-1.7069816610224897e-120, 32'sd8.288954684805044e-127, 32'sd-1.0369537082952142e-121, 32'sd0.018723430894570004, 32'sd0.022631893958170033, 32'sd0.06923888850657962, 32'sd0.010189356752011583, 32'sd0.011820137204871477, 32'sd-0.037233352732485854, 32'sd0.00827864495073126, 32'sd-0.02965011609264007, 32'sd-0.05066657309742128, 32'sd-0.013477786911756709, 32'sd0.007871803509324267, 32'sd-0.025334078840830925, 32'sd-0.0064397852662436625, 32'sd-0.06846879670913374, 32'sd-0.00010793085872922215, 32'sd-0.09560541713441652, 32'sd-0.1799051408330532, 32'sd0.018239845948348037, 32'sd0.0992715260433721, 32'sd-0.011375078116673395, 32'sd0.10083888594514043, 32'sd-0.03127871668902253, 32'sd-0.01325761318227831, 32'sd-0.004894999484939121, 32'sd2.5321701482668914e-126, 32'sd-3.8588577112220143e-115, 32'sd-9.594722614435749e-121, 32'sd-3.2225708265345676e-122, 32'sd-0.030992166810273235, 32'sd-0.08971084203253817, 32'sd0.022179976804773866, 32'sd-0.11834886168076421, 32'sd-0.0335953214028351, 32'sd-0.09290803446263216, 32'sd0.040959866188554864, 32'sd0.03463401415410106, 32'sd0.004375892333079101, 32'sd-0.0026413126783552438, 32'sd-1.2016800391987905e-05, 32'sd0.05803350762979245, 32'sd0.19887381597027723, 32'sd0.11345847587002202, 32'sd0.029838633288970354, 32'sd-0.021854538551266577, 32'sd0.03676983106005575, 32'sd-0.13152924117757633, 32'sd-0.1647230368042932, 32'sd-0.028479387069800043, 32'sd-0.05854829407387508, 32'sd-0.11606783005719022, 32'sd0.002078135767070449, 32'sd0.0438355976429806, 32'sd0.015435497459759315, 32'sd-5.082198401746852e-119, 32'sd8.620180619776188e-117, 32'sd0.06946025596698359, 32'sd0.03621326998243114, 32'sd0.07772418509154594, 32'sd0.029951711186815423, 32'sd0.037327606292255136, 32'sd0.01042680591345986, 32'sd0.036142154040580424, 32'sd-0.13675604262215169, 32'sd-0.026426984592940888, 32'sd-0.0821876786854352, 32'sd0.026875480525317106, 32'sd-0.025811228934035587, 32'sd0.004420804775882853, 32'sd0.03810383713156898, 32'sd-0.07006347692053687, 32'sd0.11676902404387458, 32'sd0.023130577378849625, 32'sd-0.007377935493017835, 32'sd0.02715586337180581, 32'sd-0.07407774811830468, 32'sd-0.013632720915118964, 32'sd-0.12316359437681419, 32'sd-0.10562966949159368, 32'sd-0.10590181898088633, 32'sd0.04993974081132052, 32'sd-0.08254712441379464, 32'sd0.029650741212795935, 32'sd-8.487330649307075e-117, 32'sd-0.04172832332717237, 32'sd-0.03769625248547299, 32'sd0.06974996694886805, 32'sd-0.02122161456197123, 32'sd-0.012683918111982084, 32'sd-0.07667971388842788, 32'sd0.05914009341878967, 32'sd-0.12150886652762277, 32'sd0.03639569145215364, 32'sd0.010856854341128782, 32'sd0.02938975329384739, 32'sd0.05186460825884665, 32'sd0.10186266384072636, 32'sd-0.030376245846268152, 32'sd0.04772637997437744, 32'sd0.03132267620413758, 32'sd0.09896806288318366, 32'sd-0.10202517013329596, 32'sd0.05735621705903754, 32'sd-0.0120141524713076, 32'sd-0.1772896666773891, 32'sd-0.04075854157963656, 32'sd0.006019174466133303, 32'sd-0.08741652249022386, 32'sd-0.06838038314878789, 32'sd0.06568754150654184, 32'sd-0.03219530641260393, 32'sd-4.295388993012967e-124, 32'sd0.022521860613690756, 32'sd-0.13140148827971693, 32'sd0.00559286452361873, 32'sd0.012020818162636076, 32'sd0.008010622789247942, 32'sd-0.026608653151098064, 32'sd0.11017884460399753, 32'sd0.03678270244691464, 32'sd0.11202878642246009, 32'sd0.07565984621053069, 32'sd0.10006944169723292, 32'sd0.16284770460162015, 32'sd0.08243377599031806, 32'sd-0.009774250904410928, 32'sd-0.06231252209657289, 32'sd0.0031691799780290113, 32'sd0.08443962734502015, 32'sd-0.01358724195999852, 32'sd-0.16289505772418766, 32'sd-0.17165279416771875, 32'sd-0.1289208608933757, 32'sd-0.19919181663429839, 32'sd-0.10914670526129379, 32'sd-0.03552780360802868, 32'sd-0.13897101268988124, 32'sd-0.08947852332771493, 32'sd0.023394406164529546, 32'sd-0.015715664291268455, 32'sd0.017023883232910066, 32'sd-0.01079139066391468, 32'sd-0.15302843067939573, 32'sd-0.0368031644418531, 32'sd-0.1323178586222344, 32'sd-0.028520299051145455, 32'sd-0.06581959752865088, 32'sd0.0075861152113856425, 32'sd0.0328448441703366, 32'sd0.09609967895793761, 32'sd0.09928579127527397, 32'sd0.004818396228891919, 32'sd0.07855609150617891, 32'sd0.0238129880871059, 32'sd-0.06341419083677806, 32'sd-0.03710918259535584, 32'sd-0.10825821982034552, 32'sd-0.05272370666558939, 32'sd-0.014194373710168825, 32'sd-0.003915511659220428, 32'sd-0.009898957638354824, 32'sd-0.07547521450276433, 32'sd-0.03275266883689949, 32'sd-0.18864985087003436, 32'sd-0.16317681868855066, 32'sd-0.04085710378664014, 32'sd-0.028687382194339542, 32'sd-0.017753719282680745, 32'sd-0.0739148719462027, 32'sd0.1010737984339856, 32'sd-0.027311812751330385, 32'sd0.043787342519294635, 32'sd0.025281219484366985, 32'sd-0.04107154360631209, 32'sd0.010115550782110395, 32'sd0.18823406286351382, 32'sd0.01821820786214457, 32'sd-0.023769445537912447, 32'sd0.04458668072898276, 32'sd0.06070129973316678, 32'sd0.018852584047060233, 32'sd-0.09732100745686696, 32'sd-0.06468096051578774, 32'sd-0.010221563433421517, 32'sd-0.08053216832626792, 32'sd0.08847681326998301, 32'sd0.055879682595830975, 32'sd0.012478861673218905, 32'sd-0.04777264812809828, 32'sd0.03319736447898439, 32'sd-0.10733494309773005, 32'sd-0.17690391113016254, 32'sd0.014570342756181255, 32'sd-0.0929749127376049, 32'sd0.040303835606006554, 32'sd-0.01401119886969269, 32'sd-0.012497828579381118, 32'sd0.11152907077807467, 32'sd-0.041537687901526045, 32'sd-0.006694888857300731, 32'sd-0.02143978909184438, 32'sd-0.013835046520538321, 32'sd-0.018541774237071092, 32'sd0.044349141517087486, 32'sd0.05125184704102149, 32'sd0.06458227842862778, 32'sd-0.02555457949207709, 32'sd-0.07930198466205954, 32'sd0.006572422287053561, 32'sd-0.09685649307892676, 32'sd0.029560330003456634, 32'sd-0.05000733151585938, 32'sd0.17054203355896452, 32'sd0.04894570622450366, 32'sd0.06529499780419813, 32'sd0.09938511520823676, 32'sd0.04357386799506398, 32'sd-0.018515377904403503, 32'sd-0.08380758724518217, 32'sd-0.07420801150995522, 32'sd0.026589535392986856, 32'sd-0.008633210800533196, 32'sd-0.029364263132379206, 32'sd0.10685013575766897, 32'sd0.03442453119571478, 32'sd-0.030766447802251844, 32'sd-0.02140908982545065, 32'sd0.004091279387719026, 32'sd-0.019170730662206346, 32'sd0.02695078790029154, 32'sd0.06298102992011578, 32'sd-0.008457219989188004, 32'sd0.0014679677001995966, 32'sd-0.16720367023448354, 32'sd-0.07493431459457332, 32'sd-0.09218361572271842, 32'sd-0.028365278551266238, 32'sd0.07102751098990544, 32'sd-0.07989962500086338, 32'sd-0.02394382931502406, 32'sd0.16555797524890928, 32'sd0.08654627183800627, 32'sd0.150100340585523, 32'sd0.11511421063292225, 32'sd0.061463677494669064, 32'sd0.111574096978051, 32'sd-0.09189045387160492, 32'sd-0.004241801637405001, 32'sd0.04857644279834728, 32'sd-0.08333114524943183, 32'sd0.03957001325747376, 32'sd0.06622204464958918, 32'sd0.01288356278547207, 32'sd-0.17138217440451667, 32'sd-0.10483729106460885, 32'sd-0.01283315500043673, 32'sd0.029137929862473894, 32'sd0.024467257443119002, 32'sd-0.04328870550431544, 32'sd0.12642641263557702, 32'sd0.026372306088243078, 32'sd-0.11404425572619403, 32'sd-0.15592926128044454, 32'sd0.02307655375236896, 32'sd0.16912051460079364, 32'sd0.15006761010736672, 32'sd0.05605511642948211, 32'sd-0.06846085230286492, 32'sd0.15477854678390834, 32'sd0.08475011430304148, 32'sd0.14134486623614162, 32'sd0.08982264525288423, 32'sd0.0016678544439280645, 32'sd-0.0328553346926737, 32'sd0.02204123260476447, 32'sd-0.09648360951642117, 32'sd0.06995411361095313, 32'sd-0.059013511858688555, 32'sd-0.0055707471840174575, 32'sd-0.0185017551927651, 32'sd-0.018465683608946473, 32'sd-0.06818479540215988, 32'sd-0.1100572961890717, 32'sd0.0059538025800056505, 32'sd0.012123988079961736, 32'sd0.04596222485466191, 32'sd-0.04692165770122874, 32'sd-0.016413248616856814, 32'sd-0.1663605756616132, 32'sd-0.10913374357750585, 32'sd-0.01639543468348604, 32'sd-0.037668668485384034, 32'sd0.15789361052866735, 32'sd0.05735452551241211, 32'sd0.13206381788781507, 32'sd0.02775332380433831, 32'sd0.08590715345745832, 32'sd0.0726954594539714, 32'sd-0.05253689537442115, 32'sd-0.01854698449729967, 32'sd0.034942567986969514, 32'sd-0.08049615718855171, 32'sd0.08597509048175764, 32'sd-0.06859163082605935, 32'sd-0.12689832528439768, 32'sd-0.02833752191247639, 32'sd-0.056590492648603205, 32'sd-0.01865291465238719, 32'sd0.045373883682605136, 32'sd0.02596344283568045, 32'sd-0.08033641456114662, 32'sd-0.06457396743967377, 32'sd0.014057422675911512, 32'sd0.11408978405152378, 32'sd0.0010117201020375995, 32'sd-0.06759092038824527, 32'sd-0.07533481590996946, 32'sd-0.055140677298817276, 32'sd0.027380516110611056, 32'sd0.04311033102339305, 32'sd0.031597155880727555, 32'sd0.0037924068153823787, 32'sd-0.03522190269430091, 32'sd-0.034295337581741324, 32'sd-0.036397574261467, 32'sd-0.06010799893249461, 32'sd-0.06598094821719726, 32'sd-0.055153925530453604, 32'sd-0.06580182016941617, 32'sd-0.013377350515578102, 32'sd-0.16789817456125963, 32'sd-0.07288461975999437, 32'sd-0.049147927856447914, 32'sd-0.07027198408831364, 32'sd0.03265460843465744, 32'sd0.06905707250157121, 32'sd0.02829348523377433, 32'sd-0.0801743656800455, 32'sd-0.045195359285321174, 32'sd0.060959796911776484, 32'sd-0.07800941490414524, 32'sd-0.05784366836393327, 32'sd-0.05077981004958966, 32'sd-0.07019829052099921, 32'sd-0.003291121954148828, 32'sd-0.043443505396743125, 32'sd0.12724122899748325, 32'sd0.023947843971003444, 32'sd0.15683628810486813, 32'sd-0.06965211938936303, 32'sd0.1029280979214071, 32'sd-0.03550179210895914, 32'sd0.050425308868584935, 32'sd-0.038361880766596565, 32'sd-0.08659589576512985, 32'sd0.033146812266985765, 32'sd-0.0369833335041186, 32'sd0.05198147121887482, 32'sd-0.05986493702669921, 32'sd-0.2179195774817335, 32'sd-0.11586954486554744, 32'sd0.033799720871350095, 32'sd-0.037865861415990916, 32'sd0.04946532495419514, 32'sd0.020298050129710084, 32'sd0.0333478375595587, 32'sd-0.02698994077584741, 32'sd-0.0714264229554559, 32'sd-0.022023006318698243, 32'sd-0.057212507734583244, 32'sd-0.14822549835750867, 32'sd-0.11464693421936141, 32'sd-0.12034403784622948, 32'sd-0.012640660315419551, 32'sd0.0021538915409031406, 32'sd0.10492671100121961, 32'sd0.07633789645297136, 32'sd0.13250210331967327, 32'sd0.0729826091423716, 32'sd0.0017054366104456457, 32'sd0.12773376270544948, 32'sd0.04765386122769205, 32'sd-0.06257612817257431, 32'sd0.013095501751507947, 32'sd-0.047815232258558674, 32'sd-0.06624986460953723, 32'sd-0.030375517020180487, 32'sd-0.1441788874643159, 32'sd-0.03530940347579815, 32'sd-0.055824712314547206, 32'sd0.013230423905604652, 32'sd0.053084191586511766, 32'sd-0.05777204066328456, 32'sd0.0416434030465116, 32'sd0.029292657952237774, 32'sd0.020847714897156172, 32'sd-0.019603002037245708, 32'sd-0.12351875762342637, 32'sd-0.1949695275315092, 32'sd-0.2137091134873236, 32'sd-0.13390325729444047, 32'sd0.12177812584871517, 32'sd-0.0018798106293079102, 32'sd-0.017330765736836517, 32'sd-0.04485084218586911, 32'sd-0.0405370333036627, 32'sd-0.01606851650577484, 32'sd0.13926922309319112, 32'sd0.12027892649350312, 32'sd0.0788953945367281, 32'sd-0.10256196842703127, 32'sd-0.12879833178682265, 32'sd-0.26922943248639997, 32'sd-0.18398700320625921, 32'sd-0.12385103550253358, 32'sd-0.14658452526975957, 32'sd-0.08983300013040103, 32'sd-0.025101262654303458, 32'sd0.02701300266360449, 32'sd-7.214914208733941e-115, 32'sd-0.0036333176124641237, 32'sd-0.022935880121920507, 32'sd-0.042451948606980025, 32'sd0.04992724809177435, 32'sd-0.01949951894921775, 32'sd-0.10007062700988067, 32'sd-0.15303479614924656, 32'sd-0.23628012009666094, 32'sd-0.2231204730402058, 32'sd-0.20679387201884514, 32'sd-0.04134712257016033, 32'sd-0.0047062271905326586, 32'sd0.10156998652497914, 32'sd-0.0771610168042053, 32'sd-0.008416195432559503, 32'sd0.11925624236435906, 32'sd0.12125315322707055, 32'sd-0.0029830373582424587, 32'sd-0.019494592864369668, 32'sd-0.13642440151451937, 32'sd-0.05497889250421163, 32'sd0.0031470300997341726, 32'sd-0.030571499416074593, 32'sd-0.009370662755209215, 32'sd0.051220242268185265, 32'sd0.0552243558079988, 32'sd0.020924331942983262, 32'sd0.018362842318198604, 32'sd0.045451633734823464, 32'sd-0.03551169844633979, 32'sd-0.032295097965101036, 32'sd-0.01318309978569662, 32'sd-0.09830215105620073, 32'sd0.010864444073847838, 32'sd-0.11463517182408721, 32'sd-0.15098264438004574, 32'sd-0.19669016014374086, 32'sd-0.1274760609766705, 32'sd-0.05305862088947089, 32'sd0.0025466630312816784, 32'sd-0.0034438497394872632, 32'sd-0.16071259239484867, 32'sd-0.14769740012219393, 32'sd0.17144050834084312, 32'sd0.10610989041868849, 32'sd0.0741329917384239, 32'sd0.023690617882879076, 32'sd-0.22282769016195317, 32'sd-0.1411319115316229, 32'sd-0.08996502362497125, 32'sd-0.09359950286075884, 32'sd0.0245193786581726, 32'sd-0.0014236244893794541, 32'sd0.03996010715525651, 32'sd-0.03829793468757434, 32'sd0.033404580128437, 32'sd-0.052403470321496656, 32'sd0.031930130668703684, 32'sd0.044859560851788945, 32'sd-0.06183781304473641, 32'sd0.010268413786325979, 32'sd0.08412379728577356, 32'sd0.050539549910975846, 32'sd0.0561992806748841, 32'sd-0.021756832545829354, 32'sd-0.14747982311836721, 32'sd-0.03073392646800233, 32'sd-0.06558887840798021, 32'sd-0.19958552032499632, 32'sd-0.09824420188138644, 32'sd-0.02704057832517635, 32'sd0.062226501728854265, 32'sd0.12455060125900656, 32'sd0.11859280253464358, 32'sd0.022795581579074513, 32'sd-0.21437840467990735, 32'sd-0.13876900587353225, 32'sd-0.08239796321613849, 32'sd-0.10946656041561006, 32'sd-0.07989576596186275, 32'sd0.07312956709200855, 32'sd-0.025372989618529778, 32'sd0.03766608415521614, 32'sd6.209671591491241e-115, 32'sd-0.07988948637353624, 32'sd-0.00818188035113786, 32'sd-0.11031857342833246, 32'sd-0.03659601809535705, 32'sd-0.014851809865519828, 32'sd0.07199746916817079, 32'sd0.023154934114614705, 32'sd-0.08491627275786666, 32'sd0.027074091158873916, 32'sd0.018213942169580777, 32'sd-0.11554502507060503, 32'sd-0.1893196018479776, 32'sd-0.1294575196626861, 32'sd-0.03681388431009711, 32'sd-0.060853441036838644, 32'sd0.001519634818519966, 32'sd-0.018667113900891867, 32'sd-0.051432336020372574, 32'sd-0.11449984979872276, 32'sd-0.1093823587665997, 32'sd-0.17556610551663682, 32'sd-0.06207254184373726, 32'sd-0.13111189498871284, 32'sd-0.17760796718885805, 32'sd-0.010487235430428777, 32'sd0.06789301326885483, 32'sd-0.04163642967448719, 32'sd0.036694166203111174, 32'sd0.05726940717783419, 32'sd-0.01589672864272168, 32'sd-0.0693996468479781, 32'sd-0.034730862529123836, 32'sd0.03503134497310055, 32'sd0.1033772449590346, 32'sd-0.021567202847463603, 32'sd-0.02461016208058663, 32'sd-0.15592490830386355, 32'sd-0.058851047835223144, 32'sd-0.11935476338341981, 32'sd-0.07749286281795034, 32'sd-0.17923517829455005, 32'sd-0.02069370026447308, 32'sd-0.011492375884854869, 32'sd0.06445138233763197, 32'sd-0.017651270276742317, 32'sd-0.029779615083005195, 32'sd-0.24715268313270433, 32'sd-0.27268690005530505, 32'sd-0.22350052115890687, 32'sd-0.058859161325629177, 32'sd-0.04665248259040002, 32'sd0.04339058813215229, 32'sd-0.13350743998844114, 32'sd0.001970336962789733, 32'sd0.06081149706227838, 32'sd0.07439552252927738, 32'sd0.03884619776204006, 32'sd0.02068200015796288, 32'sd-0.024567114724795766, 32'sd0.04265853362723856, 32'sd0.04763691418691218, 32'sd0.10123027106594061, 32'sd0.09615288410385839, 32'sd-0.0652328834058292, 32'sd-0.10229292105247441, 32'sd-0.01934393511211149, 32'sd-0.049081989400962395, 32'sd-0.048614946958804965, 32'sd-0.1397546905675297, 32'sd0.055677057173284764, 32'sd-0.02943109490006905, 32'sd-0.0018009345429844793, 32'sd-0.03254375743597849, 32'sd-0.07809267654545939, 32'sd-0.0819615731595053, 32'sd-0.2496777320102945, 32'sd-0.2462623187568388, 32'sd-0.026139712278820778, 32'sd-0.09298960216168752, 32'sd0.07145060500214678, 32'sd-0.08616090458795699, 32'sd-0.07328748540177367, 32'sd0.01719086559640246, 32'sd4.7182687210279496e-119, 32'sd0.059309601692798475, 32'sd0.07736208165527149, 32'sd0.030903019069792415, 32'sd0.019256057062953004, 32'sd0.05001934639692306, 32'sd-0.054738868479193306, 32'sd0.03511877929023325, 32'sd-0.031898261919832284, 32'sd-0.07099517380963462, 32'sd-0.005548978195426836, 32'sd0.11038189276472157, 32'sd0.05332440967086821, 32'sd-0.03913212698489073, 32'sd0.055426289745356454, 32'sd-0.0056120864080279964, 32'sd-0.020197646429091914, 32'sd-0.06885098685174995, 32'sd-0.016813196404782897, 32'sd-0.015268396460457582, 32'sd-0.1948094562679215, 32'sd-0.17040260241165736, 32'sd-0.10480365272555515, 32'sd0.03484263180666682, 32'sd-0.05683579251610823, 32'sd-0.013587215948597959, 32'sd-0.038895532232668596, 32'sd9.32910365556693e-128, 32'sd-1.0498141000457043e-121, 32'sd-3.305356224172651e-119, 32'sd0.059915743005770766, 32'sd0.042112214535662884, 32'sd-0.02182858036050503, 32'sd0.10330429110421581, 32'sd0.06496149176035308, 32'sd0.021551859011148398, 32'sd0.02878298105812987, 32'sd0.03926951994095141, 32'sd-0.031666054709527165, 32'sd-0.02089774954733382, 32'sd-0.1206039528875821, 32'sd0.035708265453839226, 32'sd-0.014250489630712095, 32'sd-0.023187358945065673, 32'sd0.13158043190063645, 32'sd-0.06264096467875503, 32'sd5.575857361966852e-05, 32'sd-0.09366378496449357, 32'sd-0.1380961774008531, 32'sd-0.1690652344641318, 32'sd-0.1200867470562308, 32'sd-0.037650807007840334, 32'sd0.041124367101591904, 32'sd0.00011197940819501805, 32'sd0.02294992011473717, 32'sd-2.9561540430957305e-118, 32'sd1.902871670643165e-120, 32'sd-1.3566090112186332e-118, 32'sd-0.025845001934915773, 32'sd-0.03135640756449409, 32'sd-0.0026116979652766933, 32'sd-0.07436698932977298, 32'sd-0.015930402339392365, 32'sd-0.035054403727098254, 32'sd-0.010279214784272375, 32'sd-0.1392642290505201, 32'sd0.11413791205237642, 32'sd-0.06601007398731794, 32'sd-0.11625362468043705, 32'sd-0.07374772172601401, 32'sd-0.08940830242778515, 32'sd-0.03458620234682096, 32'sd-0.08824255293302521, 32'sd-0.04461409919700628, 32'sd0.08315913691646117, 32'sd0.052124561613452865, 32'sd-0.09230951402419238, 32'sd-0.030362803335191195, 32'sd-0.19194511954763072, 32'sd-0.03540238511759545, 32'sd0.00801945238658286, 32'sd0.05773611520723698, 32'sd-0.08453805940891038, 32'sd9.173982572347082e-125, 32'sd-1.1131397715344343e-115, 32'sd-7.514061712493041e-120, 32'sd-5.296863817646066e-118, 32'sd0.021356217986208535, 32'sd-0.10300085604588477, 32'sd0.053054830629881713, 32'sd-0.01697098111482214, 32'sd-0.09279988913973766, 32'sd-0.09111507959278847, 32'sd-0.10016732116371754, 32'sd0.03678644832937018, 32'sd-0.05654392497470673, 32'sd-0.08843831663003976, 32'sd0.006636596801122924, 32'sd0.0469587939066966, 32'sd-0.001080070689701484, 32'sd0.10525174547866006, 32'sd0.10165754330458827, 32'sd0.1500114363684944, 32'sd0.04351391585208638, 32'sd0.10201451764647043, 32'sd0.15660662504579345, 32'sd-0.10058153822904015, 32'sd0.016760561621579854, 32'sd0.06965060498052858, 32'sd0.025463198214636718, 32'sd5.29959575295304e-128, 32'sd-7.274818580599269e-115, 32'sd-4.1974212280137315e-123, 32'sd8.403960211255983e-120, 32'sd1.3959199485452043e-117, 32'sd-1.3910745039877518e-126, 32'sd-0.015983529469431167, 32'sd0.0532570277164938, 32'sd-0.06643177385997495, 32'sd0.06910503939043632, 32'sd-0.0011124265118322653, 32'sd-0.054444944881703365, 32'sd-0.12802203564566428, 32'sd0.033276004391246894, 32'sd-0.025666003644043825, 32'sd-0.06713223228274123, 32'sd-0.03834105774364707, 32'sd0.059624916997254376, 32'sd0.0788687718350788, 32'sd0.04380402226367124, 32'sd-0.020452207447989965, 32'sd-0.019807025212444228, 32'sd-0.1139123819991803, 32'sd-0.038632406739417036, 32'sd0.022137845895090907, 32'sd0.005958797928365486, 32'sd-1.6540896961980567e-125, 32'sd1.0377060188633053e-115, 32'sd3.5331187859690265e-125, 32'sd8.351223470350373e-119},
        '{32'sd2.5065566434627838e-117, 32'sd-1.6331578561468406e-115, 32'sd-2.014432463863553e-127, 32'sd-1.2060830125249386e-117, 32'sd1.4113457966283619e-118, 32'sd6.554715125593487e-124, 32'sd-1.0677643118848885e-119, 32'sd1.5266788176801879e-115, 32'sd6.545664284072585e-124, 32'sd-1.7666365290916613e-125, 32'sd-3.789176864307695e-126, 32'sd1.0614178993704372e-122, 32'sd0.01967086683807658, 32'sd0.12506055142611902, 32'sd0.07468275510945624, 32'sd0.06014516030332823, 32'sd1.6886926759200468e-122, 32'sd2.2857814843256778e-121, 32'sd-2.379430901064502e-127, 32'sd-1.6132793042190606e-115, 32'sd9.544466516288093e-124, 32'sd7.342553783511437e-117, 32'sd3.655469247018386e-129, 32'sd1.1591875913778514e-118, 32'sd-5.4019887175274165e-118, 32'sd-6.582334005369538e-128, 32'sd1.1733537534031258e-118, 32'sd6.937134143935215e-117, 32'sd-4.726900636510415e-123, 32'sd2.5994008417497163e-123, 32'sd-5.773648728225539e-127, 32'sd2.9942378682482037e-123, 32'sd0.017100169274652494, 32'sd0.06249490295280298, 32'sd0.01891989691538293, 32'sd0.1130270179240945, 32'sd0.08606919857801291, 32'sd0.07498755061464141, 32'sd0.0952397707451418, 32'sd0.07372994005696468, 32'sd0.05004123113377734, 32'sd0.032364225096068316, 32'sd0.05024360033034817, 32'sd0.03041597035286762, 32'sd0.07145007712229519, 32'sd0.01713190942949129, 32'sd0.04029053413322798, 32'sd-0.016775351942250914, 32'sd0.03918417140214949, 32'sd-0.008849708030034806, 32'sd0.030770307023169914, 32'sd0.016073337126373835, 32'sd4.140815730938701e-124, 32'sd1.5517310160318283e-115, 32'sd6.5332896744885055e-124, 32'sd-2.0105501149527107e-116, 32'sd-8.794506492178869e-119, 32'sd6.962786056454646e-117, 32'sd0.10336736756966, 32'sd-0.0023767384897531757, 32'sd-0.0010213997423932498, 32'sd0.06914004117016619, 32'sd0.06767304215086746, 32'sd-0.02374343415112422, 32'sd-0.012473644359518556, 32'sd0.003426354128436317, 32'sd0.022681493686617517, 32'sd-0.012219987076195246, 32'sd0.00983757729573269, 32'sd-0.1634543265810143, 32'sd-0.0639941861258812, 32'sd-0.047005317794081077, 32'sd0.0011800743082547476, 32'sd0.05303184203222185, 32'sd0.03941642324576761, 32'sd0.022973797037920896, 32'sd0.01879782464257156, 32'sd0.11674688865456408, 32'sd0.10113255530025196, 32'sd0.057018599866507085, 32'sd0.09253390143316832, 32'sd0.07160833862655976, 32'sd-7.315228004367427e-117, 32'sd3.6697708915256454e-116, 32'sd1.678130856012654e-122, 32'sd1.62125420861142e-125, 32'sd0.07730860075261575, 32'sd-0.0014181127095076527, 32'sd-0.003410443815756558, 32'sd-0.03727843343801616, 32'sd-0.007617516183743709, 32'sd-0.06068197298781837, 32'sd-0.08406831499676341, 32'sd0.06338233806833746, 32'sd-0.027435448286338208, 32'sd-0.020429930355703625, 32'sd0.0863925466825028, 32'sd-0.010466850958828239, 32'sd-0.019438211365953396, 32'sd-0.062138667394166215, 32'sd-0.04601425302444249, 32'sd-0.14433850377833612, 32'sd-0.09685975146262578, 32'sd0.04699357395294425, 32'sd0.03738089108175904, 32'sd0.12383052013412094, 32'sd-0.017057761796009412, 32'sd-0.0063989251829274915, 32'sd0.08714809786254835, 32'sd0.055995075446586766, 32'sd-0.021609687782637655, 32'sd2.4503272682292995e-126, 32'sd1.5255380712841514e-123, 32'sd0.01290884178258344, 32'sd-0.08100877679765645, 32'sd0.02566681945257406, 32'sd0.0700790409871342, 32'sd-0.008886853462345778, 32'sd0.10513246438137666, 32'sd0.030440931134405446, 32'sd-0.005921078036013148, 32'sd-0.07439098824870768, 32'sd-0.06200097263510491, 32'sd-0.016818377266954596, 32'sd-0.08699063503838166, 32'sd-0.00582303193356199, 32'sd0.0023430157469992437, 32'sd-0.05546757786899762, 32'sd0.043365498465276826, 32'sd0.07393083444643027, 32'sd0.13179367387390387, 32'sd0.10708589415737313, 32'sd0.11251644579515903, 32'sd0.135588204246076, 32'sd-0.03937011892718788, 32'sd0.009274500399186644, 32'sd0.13478732735355978, 32'sd-0.042226442293403256, 32'sd0.039750498662669685, 32'sd0.025583423659621657, 32'sd1.3404548893746617e-118, 32'sd-0.012047669401086768, 32'sd0.14083301625923453, 32'sd-0.049470116348060526, 32'sd-0.019456529757126466, 32'sd0.035794138740867086, 32'sd-0.06148052240146678, 32'sd-0.04057015108481621, 32'sd0.01965762078935961, 32'sd-0.017824184412094147, 32'sd0.09707874431712654, 32'sd0.07604296333913091, 32'sd-0.04954000692002036, 32'sd-0.07313978088249487, 32'sd-0.09758013705607457, 32'sd0.04362202848670598, 32'sd-0.05332821906364289, 32'sd0.1077297235670147, 32'sd-0.027805185510407636, 32'sd0.018842388129336394, 32'sd0.04100710813150494, 32'sd0.12453303152305226, 32'sd0.11344417166178089, 32'sd-0.00979444602004469, 32'sd0.08403317491144327, 32'sd0.025355213208688738, 32'sd-0.00993622592554992, 32'sd0.018146578402822813, 32'sd-7.898743057212212e-127, 32'sd0.025059206678808534, 32'sd0.03064013588287674, 32'sd-0.05668275621130273, 32'sd0.023830299990109004, 32'sd0.0432860183620002, 32'sd-0.02666232315704948, 32'sd-0.06769293553057733, 32'sd0.008715406025045808, 32'sd0.028807044712068235, 32'sd-0.012550211949977609, 32'sd-0.026006208089405923, 32'sd-0.03385354087413589, 32'sd-0.024638007052338307, 32'sd-0.036345223935384634, 32'sd-0.08031619480415923, 32'sd0.03042596919417823, 32'sd0.014820021490569931, 32'sd0.007317710632841198, 32'sd-0.003978327130784845, 32'sd0.07009264511442276, 32'sd0.024859843170561065, 32'sd0.011463972120052766, 32'sd0.0007705678764118703, 32'sd0.07658546319939506, 32'sd0.04678206867031306, 32'sd0.032000941258372544, 32'sd-0.058735037052783684, 32'sd0.056503749882504554, 32'sd-0.058212300952419346, 32'sd0.012260437055960385, 32'sd0.06838662877066179, 32'sd0.023441903589842748, 32'sd-0.0014041085366409886, 32'sd0.00592728285917398, 32'sd0.01122701945737408, 32'sd0.11864573479007086, 32'sd-0.08874454223969035, 32'sd-0.0037137351845097297, 32'sd-0.11706327889632978, 32'sd-0.06796332271724859, 32'sd0.08226523054583526, 32'sd-0.04019071642072397, 32'sd0.03868860989522457, 32'sd-0.03963485208704607, 32'sd-0.02651941453476996, 32'sd0.0022477692711335294, 32'sd-0.009993247582169169, 32'sd-0.03395763687290502, 32'sd-0.06153763459857213, 32'sd0.12542030363177675, 32'sd-0.08789888585041078, 32'sd0.004064830801802977, 32'sd-0.02072802087555721, 32'sd0.07422508857145446, 32'sd0.028764532562292836, 32'sd0.011215679768040176, 32'sd0.07261872170075896, 32'sd0.04272634782605983, 32'sd0.08380726443895498, 32'sd0.17175425147347337, 32'sd0.06170399496078271, 32'sd-0.08526442048861851, 32'sd-0.009372456137264258, 32'sd0.04947553387900151, 32'sd-0.045186292117513814, 32'sd0.04733056993134393, 32'sd0.04693062818243131, 32'sd0.01932900054068017, 32'sd0.09724111308507435, 32'sd0.06908655696519027, 32'sd0.005721228218866139, 32'sd0.04515222569360141, 32'sd-0.12129687455961755, 32'sd-0.04380112662474427, 32'sd0.04804332366773786, 32'sd0.014005681525332003, 32'sd-0.09461185875592687, 32'sd-0.07855353490063274, 32'sd0.041000016433825635, 32'sd0.03525660985714101, 32'sd-0.0667106528099303, 32'sd0.03012597958745522, 32'sd0.021763982255231726, 32'sd0.03702902798429964, 32'sd0.025977425016896143, 32'sd0.006634964574275928, 32'sd0.08322095940418855, 32'sd0.05356597987392695, 32'sd-0.024537038213357745, 32'sd-0.04947618893271178, 32'sd0.064681032591282, 32'sd0.07282786135238807, 32'sd0.03719383946161939, 32'sd0.198682826084517, 32'sd0.04552629189141368, 32'sd0.1760288940514277, 32'sd0.16903271218295987, 32'sd0.15796793963106917, 32'sd0.01042432820535212, 32'sd0.10905581629066995, 32'sd0.05976950398336023, 32'sd0.03392079334311613, 32'sd0.01542578428510256, 32'sd0.03349196588918721, 32'sd-0.006354293427965096, 32'sd-0.026504202618879126, 32'sd0.11887978439839174, 32'sd0.0439285177063544, 32'sd0.004969920817117029, 32'sd0.13796407737913507, 32'sd0.07383146560654705, 32'sd-0.05144090759466352, 32'sd0.021765682274261962, 32'sd0.11906739147817014, 32'sd0.15869926717716462, 32'sd-0.01535081347249872, 32'sd-0.017557406337423965, 32'sd0.07334782182593358, 32'sd0.08053459626308157, 32'sd0.05621969040376493, 32'sd0.09975749621412688, 32'sd0.20954310074079655, 32'sd0.18628058123170851, 32'sd0.012548216497173937, 32'sd-0.03909516836980973, 32'sd-0.12976259861762487, 32'sd0.018822931932270724, 32'sd0.00033998019199470234, 32'sd-0.09057453041770576, 32'sd0.001310535300587643, 32'sd-0.044090093089022286, 32'sd0.09764155422259908, 32'sd-0.0014844097617978142, 32'sd-0.06500773197969757, 32'sd0.010764919783286184, 32'sd-0.04786379906712615, 32'sd0.07180611852679697, 32'sd0.16866440113217945, 32'sd-0.038271075189985, 32'sd0.06655277896304251, 32'sd-0.034360035373366314, 32'sd0.06790528862642943, 32'sd0.052192486341134034, 32'sd-0.03987419983421867, 32'sd0.13458433244548898, 32'sd0.07545899216417461, 32'sd0.13589276568823175, 32'sd-0.05212803823061767, 32'sd0.16474671867370771, 32'sd0.06988422667729646, 32'sd0.07694369692068247, 32'sd-0.0892401277789906, 32'sd-0.29305364307310444, 32'sd-0.24999780467565413, 32'sd-0.022954476490069823, 32'sd0.14101717337463696, 32'sd-0.04714894276961938, 32'sd-0.039444247833332356, 32'sd0.043488231672416965, 32'sd-0.008862626079574795, 32'sd0.04138281046558026, 32'sd-0.02808812730213222, 32'sd-0.007528094908837944, 32'sd-0.0577262583278245, 32'sd0.07627247463346815, 32'sd0.06383487451462665, 32'sd0.05249450350241491, 32'sd0.014565024270765718, 32'sd-0.043631886836847364, 32'sd0.06533498130553822, 32'sd0.078630899682838, 32'sd0.05228687534771083, 32'sd0.08740410407310678, 32'sd0.055200743822131304, 32'sd0.13147747737275395, 32'sd-0.027860486677032358, 32'sd-0.03997413239635444, 32'sd-0.15957235678413462, 32'sd-0.1028573726538387, 32'sd-0.07717842591278988, 32'sd-0.2686718937637175, 32'sd-0.29393018359476913, 32'sd-0.12267465784917629, 32'sd-0.06564084101173194, 32'sd-0.008394819396727593, 32'sd0.025449103896051713, 32'sd5.746142518240741e-05, 32'sd0.05870009144717244, 32'sd-0.05033787924518255, 32'sd-0.03676688476060399, 32'sd-0.07928887488702237, 32'sd0.061282463237945915, 32'sd0.04281300499909384, 32'sd-0.03821822127179426, 32'sd-0.062397884836273475, 32'sd0.059422679825434525, 32'sd0.047832617649458314, 32'sd0.019165210835287234, 32'sd0.020803205502277922, 32'sd0.016156806395748652, 32'sd-0.08144115685641011, 32'sd-0.017089468869752458, 32'sd-0.05709815354489937, 32'sd-0.04520949152020781, 32'sd-0.005910726313517187, 32'sd-0.19537501054995093, 32'sd-0.14501938793748062, 32'sd-0.11979993324240679, 32'sd-0.1503051414109186, 32'sd-0.11496135631569714, 32'sd-0.07155322409423559, 32'sd-0.1922560793787191, 32'sd-0.022961125532651214, 32'sd-0.06868977518596273, 32'sd0.010163225944029325, 32'sd-0.06253506095548583, 32'sd-0.027444431193355552, 32'sd-0.07921256554268488, 32'sd0.048821390368250235, 32'sd0.09517545885527347, 32'sd-0.04844225296244915, 32'sd0.08174669222867018, 32'sd0.003550142413529422, 32'sd0.01267006536441776, 32'sd-0.0010261535315906898, 32'sd0.08180335476559833, 32'sd0.007672294175545082, 32'sd-0.0034441707110874384, 32'sd-0.04458642086352072, 32'sd-0.13358052214681568, 32'sd-0.1955149025454664, 32'sd-0.33218331630630976, 32'sd-0.23517594930505464, 32'sd-0.11582009685394896, 32'sd-0.1624204051236999, 32'sd-0.18919083545077733, 32'sd-0.004329374015258795, 32'sd-0.10596980257687744, 32'sd-0.07802858304243535, 32'sd-0.22461460602435562, 32'sd-0.08789574114121906, 32'sd-0.1070603104109046, 32'sd-0.054566499159740156, 32'sd0.039510382609316594, 32'sd-0.04013973323941113, 32'sd-0.04392332678447821, 32'sd-0.06936846139711128, 32'sd-0.007787952971123754, 32'sd-0.06063561048048959, 32'sd0.00662235407626571, 32'sd0.011458880013245331, 32'sd0.04617259006586585, 32'sd-0.027629413799831762, 32'sd0.040864256973841336, 32'sd-0.08610416258024922, 32'sd-0.14023733974833535, 32'sd-0.17097885254464135, 32'sd-0.22241822890305996, 32'sd-0.17202829433581132, 32'sd-0.27515367483025255, 32'sd-0.20084836833406275, 32'sd-0.12678421558960598, 32'sd-0.1766010061220163, 32'sd-0.08417991111472921, 32'sd0.11450442894529321, 32'sd-0.0011005593938808542, 32'sd-0.15308298592795103, 32'sd-0.17440615803545098, 32'sd-0.11348083299972565, 32'sd-0.10479167298592779, 32'sd-0.041726847021471794, 32'sd-0.12878442753230898, 32'sd-0.1416053051863285, 32'sd-0.03720426181346117, 32'sd-0.004979591636099863, 32'sd0.06366484083955083, 32'sd-0.015549687945066129, 32'sd-0.01904598208720631, 32'sd0.03750647434247164, 32'sd0.060182362441846354, 32'sd0.02955776346712202, 32'sd0.03502863426671076, 32'sd-0.13006659019748057, 32'sd-0.19796291976878166, 32'sd-0.24792019252645892, 32'sd-0.2567279312724047, 32'sd-0.155577330839299, 32'sd-0.17717748510791706, 32'sd-0.05451789090932761, 32'sd-0.11992934509850267, 32'sd-0.01068004600639096, 32'sd0.10648283538270005, 32'sd0.03711284185611657, 32'sd0.16693672860474298, 32'sd-0.011796165014911795, 32'sd-0.0067165754486304035, 32'sd-0.06625488459869516, 32'sd-0.03358352070436307, 32'sd-0.038469664054581375, 32'sd-0.2240659595398122, 32'sd0.002216605800872573, 32'sd0.07284719103075803, 32'sd0.024959572853560544, 32'sd-0.03209918651376077, 32'sd0.0826726951440153, 32'sd-0.016438367175691332, 32'sd0.08374268349776035, 32'sd-1.0365198263887466e-123, 32'sd0.065889547300192, 32'sd-0.008942809414612686, 32'sd-0.09145136066175129, 32'sd-0.01777572046944657, 32'sd-0.0747694637973014, 32'sd-0.13036803467977964, 32'sd-0.12315867864232365, 32'sd-0.06410849178219616, 32'sd0.08351677341934051, 32'sd0.1378062064459963, 32'sd0.08033134710919895, 32'sd0.11464103773795847, 32'sd0.15839156334298196, 32'sd0.06752597579100043, 32'sd-0.054021210639127175, 32'sd-0.01295619038669651, 32'sd-0.11539492503153155, 32'sd-0.09432246266923669, 32'sd-0.08569387333948941, 32'sd-0.14701198035870597, 32'sd5.471072544699596e-05, 32'sd-0.01118466989862166, 32'sd0.039465569279507826, 32'sd0.11505881506561284, 32'sd0.18301755554461752, 32'sd-0.02304320640875565, 32'sd0.046017250167727494, 32'sd0.03423714245754365, 32'sd-0.038571094768243594, 32'sd0.09069047524299449, 32'sd0.029791766936454394, 32'sd0.08409747098471149, 32'sd-0.08755157661080992, 32'sd0.026605481054213037, 32'sd-0.11784030491629591, 32'sd0.05138233442784331, 32'sd0.06752102027859348, 32'sd0.21334965760151076, 32'sd-0.013007549987198365, 32'sd0.0383460963473165, 32'sd0.10106288879714088, 32'sd0.05438518136336267, 32'sd0.13782358126485827, 32'sd-0.01955341938734844, 32'sd-0.06119101800655389, 32'sd-0.05060406399108897, 32'sd-0.006202230106475588, 32'sd0.01119422951207453, 32'sd0.04337611011129592, 32'sd-0.037937881977591834, 32'sd-0.14000666742069412, 32'sd-0.026266334003598783, 32'sd0.023940049369472832, 32'sd0.10837590862269084, 32'sd0.011880967249630102, 32'sd0.04662815967647275, 32'sd-0.054336520429582, 32'sd0.012545536922942281, 32'sd-0.00589113376290186, 32'sd0.08979141979888638, 32'sd-0.013528136888793486, 32'sd-0.08781132840913593, 32'sd0.11274804223358494, 32'sd0.17613447999881038, 32'sd0.14658207932629477, 32'sd0.02266142784560357, 32'sd0.026391710056259492, 32'sd0.038917876856792044, 32'sd0.0392180610356374, 32'sd0.049188391832513625, 32'sd0.09182303150301455, 32'sd0.16845575541693084, 32'sd0.1538595688209108, 32'sd0.07974339941932128, 32'sd0.0029024718824564645, 32'sd0.08010839809643705, 32'sd-0.04694322078707173, 32'sd-0.03369990431594527, 32'sd-0.03088119048046591, 32'sd0.09897565539602715, 32'sd0.1049349985691415, 32'sd0.08809768295499955, 32'sd0.012759201308173346, 32'sd2.1163508862399218e-125, 32'sd-0.0041015681422058425, 32'sd0.010783940335000963, 32'sd0.04602323969319826, 32'sd0.0019369726731480062, 32'sd-0.024938601647427814, 32'sd0.057390775875626056, 32'sd0.0942977493089759, 32'sd0.20535317832261235, 32'sd0.10814201295743116, 32'sd0.055772041451700394, 32'sd-0.007798440452080424, 32'sd0.08884638408039651, 32'sd0.12638958666859668, 32'sd0.10984413867915639, 32'sd0.16455378918558944, 32'sd0.03131859147689003, 32'sd0.1644463869065323, 32'sd0.010090122833920015, 32'sd0.0871125235256109, 32'sd-0.04391636348396524, 32'sd0.04316128300018069, 32'sd-0.10625879635015512, 32'sd-0.054635831457969956, 32'sd0.027454228831090454, 32'sd0.019111402423642995, 32'sd0.08094525512323933, 32'sd0.015204022661105513, 32'sd0.06597432106796954, 32'sd0.042283523841491456, 32'sd0.010226784668750868, 32'sd0.15788817640015654, 32'sd0.07829954537232789, 32'sd0.13271232970535787, 32'sd0.11917631144636719, 32'sd0.04625479788051278, 32'sd0.031014005132712155, 32'sd0.059605062567783605, 32'sd0.03361326329364942, 32'sd0.05113482048698225, 32'sd-0.0118849744432795, 32'sd0.12490243821918877, 32'sd0.10124347787867505, 32'sd0.1586144284882458, 32'sd0.1316775233355461, 32'sd0.1498931858708951, 32'sd0.13621199213405175, 32'sd0.13350041182104486, 32'sd0.01818155994200628, 32'sd-0.06200947207685376, 32'sd-0.052344642071825626, 32'sd0.05533461757272561, 32'sd0.10515599078373418, 32'sd0.06349918134730721, 32'sd0.11209176199527565, 32'sd-0.05885620518832055, 32'sd0.004378571233679162, 32'sd-0.013463324689728615, 32'sd0.02931785627861329, 32'sd0.04263466026348642, 32'sd0.09990877887736313, 32'sd0.0035672273601629893, 32'sd0.05274720384059821, 32'sd0.08192643635885151, 32'sd0.03417201461640292, 32'sd0.02409894321440308, 32'sd0.0346940251232237, 32'sd0.04763854547271233, 32'sd-0.051626463151248046, 32'sd0.11357798655002513, 32'sd-0.045882208810795376, 32'sd0.147423571584377, 32'sd0.10243849949249305, 32'sd0.15429875350901773, 32'sd0.07822028409746956, 32'sd0.018691581690705953, 32'sd-0.008524241160000057, 32'sd-0.03559781075057494, 32'sd-0.038396275024029605, 32'sd0.0407202404082955, 32'sd-0.033407332027904156, 32'sd0.057779330344540025, 32'sd0.07252328359506144, 32'sd0.04156840913411428, 32'sd-7.239531916196943e-127, 32'sd0.02695763035708694, 32'sd0.056347703975272244, 32'sd0.06384340636088873, 32'sd-0.0050825331975211845, 32'sd0.07730824144133779, 32'sd0.09479772613475645, 32'sd0.041768961361970766, 32'sd0.10945583541356407, 32'sd0.0849104723354169, 32'sd0.08510771958300047, 32'sd-0.01742395615191402, 32'sd0.11671204974648271, 32'sd0.11086337191068085, 32'sd-0.021732149934230942, 32'sd0.04488637178372462, 32'sd0.11335883177673185, 32'sd0.019472974587522417, 32'sd0.05176184072274844, 32'sd0.01897736889020355, 32'sd0.10156839770016148, 32'sd-0.06472447673148976, 32'sd-0.03488156699556167, 32'sd0.04992156186351922, 32'sd-0.04700573124926184, 32'sd-0.06458813451710678, 32'sd-0.01949178958129905, 32'sd-2.0862943470043798e-127, 32'sd8.137282428857634e-116, 32'sd1.1671415077185723e-115, 32'sd0.015655258745598696, 32'sd-0.06415971722329204, 32'sd0.08421581374395411, 32'sd0.026211796557021164, 32'sd0.045618560589893324, 32'sd0.039057942224190983, 32'sd0.06554858345020942, 32'sd0.0878079290830564, 32'sd0.06333993761886746, 32'sd0.06431022265006998, 32'sd0.006942627416081896, 32'sd0.07938216958435322, 32'sd-0.028899397050491906, 32'sd0.06921554668128614, 32'sd0.07086837088294255, 32'sd0.06382375452545702, 32'sd0.08669326215020885, 32'sd0.14626187073594127, 32'sd0.11134602419811858, 32'sd-0.009027610863685124, 32'sd0.018072522964433013, 32'sd-0.018694914172166174, 32'sd0.07636567025429775, 32'sd0.03283499590804261, 32'sd-0.07774035724431723, 32'sd-1.36499837270795e-119, 32'sd1.0232581137958617e-119, 32'sd6.539939835880898e-125, 32'sd-0.07712796743697464, 32'sd-0.02746219518448954, 32'sd-0.06695934734916163, 32'sd0.05525109214206573, 32'sd-0.00360035903800219, 32'sd-0.00032372028650739935, 32'sd0.04701728050728201, 32'sd0.08371214213737055, 32'sd-0.005857351698669587, 32'sd0.01219934147587016, 32'sd0.08339532477692857, 32'sd0.09089716236900003, 32'sd0.01204008875469627, 32'sd-0.05505569882979711, 32'sd0.0430964394463212, 32'sd0.04601484256339358, 32'sd0.04640714297493252, 32'sd0.04501032584149589, 32'sd-0.0021344220199796212, 32'sd0.038574826358586924, 32'sd-0.031922413269221094, 32'sd-0.0830846660428967, 32'sd0.03801413083571425, 32'sd0.00603962483486975, 32'sd0.034475809000367154, 32'sd-1.0787188268694218e-124, 32'sd1.2121008113567365e-122, 32'sd-7.401092530305053e-127, 32'sd-7.565159431026828e-127, 32'sd0.023900298211176108, 32'sd-0.08173011057028051, 32'sd-0.018072796365748097, 32'sd-0.015418673758031173, 32'sd0.11883556076894039, 32'sd0.09908843141763876, 32'sd0.0465215490878963, 32'sd-0.04116100005383184, 32'sd0.028346537932406678, 32'sd-0.05945395383117285, 32'sd0.0883704462929625, 32'sd0.021992164683156065, 32'sd0.0751789927150503, 32'sd-0.00224564311685691, 32'sd0.038338789974335964, 32'sd0.009872394021417057, 32'sd0.08452299100431619, 32'sd-0.0007491058642230866, 32'sd-0.04089960856580768, 32'sd0.004865314667537181, 32'sd-0.09661620190654695, 32'sd0.058174148263142815, 32'sd0.022255609213874875, 32'sd6.443646924847904e-126, 32'sd-5.584791588676611e-117, 32'sd2.284439692732397e-117, 32'sd-1.5790279595257889e-117, 32'sd8.380078511857366e-127, 32'sd6.273240765738313e-125, 32'sd0.06977399364047614, 32'sd0.0510066723578961, 32'sd0.04894066432519655, 32'sd-0.030008286034827115, 32'sd-0.028670710210372922, 32'sd0.043015677519035525, 32'sd0.10137266259885239, 32'sd-0.010230797138398475, 32'sd-0.0569306917125255, 32'sd0.12150028113132093, 32'sd0.0711420873266896, 32'sd-0.03603050427355687, 32'sd0.09151524033870645, 32'sd0.09338156720637815, 32'sd-0.006974328724979777, 32'sd-0.06310842883109263, 32'sd0.08688064082728038, 32'sd-0.05437245381854916, 32'sd-0.00873839635336929, 32'sd0.03483053555871218, 32'sd5.17286603508694e-122, 32'sd-1.6955981493672928e-123, 32'sd-3.663620194858193e-119, 32'sd3.0087026528752203e-118},
        '{32'sd-1.0824531129427174e-125, 32'sd2.320401586376534e-121, 32'sd-2.7182625000461214e-127, 32'sd-8.138250830637774e-115, 32'sd1.2231527002611445e-120, 32'sd1.0865247313567512e-123, 32'sd-1.8646236495298538e-128, 32'sd-1.7238805143900923e-116, 32'sd3.3270918529690066e-125, 32'sd3.4009028828804007e-127, 32'sd9.348602062835759e-122, 32'sd9.756956574057083e-129, 32'sd0.08182370492071336, 32'sd0.030259922596976664, 32'sd0.017592857200553178, 32'sd-0.01481346758750429, 32'sd-1.2298752886645467e-120, 32'sd2.3811306198113117e-128, 32'sd-6.60007021211031e-115, 32'sd-8.163178047925346e-127, 32'sd-1.9458769636408444e-123, 32'sd-6.149173965701447e-121, 32'sd2.616855052086665e-126, 32'sd9.94439198973549e-121, 32'sd1.531924059218788e-123, 32'sd6.829472866811606e-124, 32'sd1.933558250776897e-118, 32'sd-5.891384771946825e-124, 32'sd8.55359900009355e-125, 32'sd1.398610182176949e-123, 32'sd-3.054724240291539e-126, 32'sd-2.1092779302786526e-117, 32'sd0.01758955374164752, 32'sd-0.040373110169590845, 32'sd-0.036597427156780105, 32'sd-0.07505040279987636, 32'sd0.04519354861026124, 32'sd-0.021893198017701652, 32'sd-0.05313717497591069, 32'sd0.03321839471264586, 32'sd0.03587177307678256, 32'sd-0.03134680937383637, 32'sd-0.040365009817895633, 32'sd0.06171778219409745, 32'sd-0.054856190677841976, 32'sd0.00017271530333443544, 32'sd0.0496880731683416, 32'sd-0.015006750038503146, 32'sd0.02681736097712095, 32'sd0.07981035156270777, 32'sd-0.003997432056012215, 32'sd0.0032475351201555515, 32'sd-1.1110981529170536e-119, 32'sd-4.6118053890325334e-119, 32'sd-9.536049612406301e-118, 32'sd6.490939508552426e-126, 32'sd2.6578615940358846e-127, 32'sd2.111045802798698e-117, 32'sd-0.01093624718561643, 32'sd-0.018399277811919756, 32'sd-0.017731812695562073, 32'sd0.005936918139943272, 32'sd-0.005756914785421467, 32'sd0.013914264853885248, 32'sd0.048729963978677016, 32'sd-0.018978939504415013, 32'sd-0.08613960638356437, 32'sd-0.0028538234731142306, 32'sd0.09097532208830919, 32'sd-0.03925928114691814, 32'sd-0.09895140895291094, 32'sd-0.1952453215236712, 32'sd-0.12665272168158231, 32'sd-0.03549257751948682, 32'sd-0.13492447301785812, 32'sd-0.0945287209375088, 32'sd-0.003021523960220128, 32'sd-0.004885151407997283, 32'sd-0.026649843825001008, 32'sd0.025036734518402284, 32'sd0.005305053675156103, 32'sd-0.0038161167748587328, 32'sd-6.8891770916238e-126, 32'sd-2.915418378495111e-116, 32'sd-1.1391503908071411e-119, 32'sd2.395718488887237e-121, 32'sd0.016482768547115056, 32'sd-0.002168875738108458, 32'sd-0.044984075840080295, 32'sd-0.12485302950480814, 32'sd-0.08587503668190193, 32'sd-0.04569292709956418, 32'sd-0.0707579251413768, 32'sd0.008335959413534766, 32'sd0.01863776873318142, 32'sd0.004921675697266, 32'sd-0.07312937316249203, 32'sd0.0453515166083879, 32'sd0.10193810397680561, 32'sd0.05875480505595048, 32'sd-0.04863614907057305, 32'sd0.06826226914853575, 32'sd0.0795458898463226, 32'sd0.14846455192322358, 32'sd0.09021921981947588, 32'sd-0.03030888313573872, 32'sd0.08443541764874637, 32'sd-0.03042699973101109, 32'sd-0.033505006494651574, 32'sd0.057556610266035986, 32'sd0.07277358894021713, 32'sd1.3716446244945173e-115, 32'sd-9.022749671505285e-124, 32'sd-0.01067156507075595, 32'sd-0.0550337020760039, 32'sd0.06871657566823225, 32'sd0.05757236447747443, 32'sd0.048137503493492766, 32'sd-0.01465165236356331, 32'sd0.014402554768012187, 32'sd-0.0669078817057435, 32'sd-0.021970012960156927, 32'sd-0.16051639720880578, 32'sd-0.024403500419355215, 32'sd-0.06944118189658713, 32'sd0.17146588290695045, 32'sd0.07895092250823707, 32'sd0.04479306955456635, 32'sd0.05125318926674153, 32'sd0.10595719002319405, 32'sd0.09080954585301082, 32'sd0.010420291688108705, 32'sd0.07221622791182628, 32'sd0.05618897433469992, 32'sd0.0442975654703126, 32'sd0.04309947340689212, 32'sd-0.07308770802308841, 32'sd-0.10917653104447146, 32'sd0.08030806720032298, 32'sd-0.009944570359645105, 32'sd3.4896114925037935e-116, 32'sd0.05934072011690929, 32'sd-0.021928233130238513, 32'sd0.03840855520434759, 32'sd-0.17083436043132483, 32'sd-0.048813628917596046, 32'sd-0.02365615542509839, 32'sd-0.1343398523534284, 32'sd-0.06475166632293335, 32'sd0.01067451828441051, 32'sd-0.10294753199782856, 32'sd-0.2172264552139226, 32'sd-0.13284873052489238, 32'sd-0.02876077549998926, 32'sd0.030522595906225265, 32'sd0.11353595917582388, 32'sd0.1371053686923159, 32'sd0.003974021604320441, 32'sd0.11757167546761375, 32'sd0.07755093152641135, 32'sd-0.03705605602853269, 32'sd0.08220704767560712, 32'sd0.021684915543976727, 32'sd-0.00831991769855909, 32'sd-0.12966728914010364, 32'sd-0.079111910964901, 32'sd0.080547707693387, 32'sd0.07174932447274741, 32'sd1.199384692871644e-117, 32'sd-0.00733015352758001, 32'sd0.03636113750061412, 32'sd0.03493416285635457, 32'sd-0.015615169336058317, 32'sd-0.08630086069872377, 32'sd-0.043679159044280755, 32'sd-0.06908616063525788, 32'sd0.047496769833208496, 32'sd-0.04689344362577878, 32'sd0.002511457474227299, 32'sd-0.07396313782219809, 32'sd-0.09108823956010353, 32'sd-0.05444261339339698, 32'sd0.03175813410503766, 32'sd-0.030699423679914673, 32'sd0.053344628899757655, 32'sd0.07359575816386923, 32'sd0.04734259918482218, 32'sd0.01957975264830931, 32'sd-0.04209663525195009, 32'sd-0.016654854099282527, 32'sd0.0665331029930702, 32'sd-0.05728398206224031, 32'sd5.953011214178917e-06, 32'sd-0.008761762298338381, 32'sd0.018403101479525136, 32'sd0.09455437367102729, 32'sd-0.01826898245761636, 32'sd-0.031087197025197657, 32'sd0.115588202748502, 32'sd0.025665039141054623, 32'sd-0.01914782484359863, 32'sd0.05051182280689988, 32'sd0.09756382887220523, 32'sd0.039046028515800864, 32'sd0.04321986428185273, 32'sd0.09558409080955546, 32'sd-0.0015617241591625725, 32'sd-0.008572554076184067, 32'sd-0.0029322661489006308, 32'sd-0.0670913432493593, 32'sd-0.0029522032465325947, 32'sd-0.07194304215362245, 32'sd0.10495525377825696, 32'sd-0.04813185671867553, 32'sd0.016676894293948502, 32'sd0.1594782702808173, 32'sd0.16333374259984743, 32'sd0.09240967780103973, 32'sd0.01867279054399996, 32'sd0.09626664084424931, 32'sd-0.0042806147527028595, 32'sd0.0003455008468878709, 32'sd0.010512191604314637, 32'sd0.06676462516827936, 32'sd-0.0018563080162274513, 32'sd0.02806632153434128, 32'sd0.05413468203705635, 32'sd-0.09778033482084855, 32'sd-0.01878686372274698, 32'sd-0.010593135941712071, 32'sd0.09566846226211932, 32'sd0.07850801909625764, 32'sd0.07379547071644328, 32'sd0.045800427835475464, 32'sd0.02564156233530969, 32'sd-0.10717758590796943, 32'sd-0.11469267465652083, 32'sd-0.06329545089640978, 32'sd0.026957761677242054, 32'sd0.13882718392259258, 32'sd0.08750685281859305, 32'sd-0.09663266044998882, 32'sd-0.09299803177539588, 32'sd0.07729569786896023, 32'sd0.06973550009407878, 32'sd0.031120599935002557, 32'sd-0.0075027724605530345, 32'sd0.03923174047070035, 32'sd-0.048388967371553585, 32'sd0.039709726654046186, 32'sd-0.08621744700506064, 32'sd0.03852067212474897, 32'sd0.019974706554688595, 32'sd-0.04739612411843727, 32'sd-0.002648232349254217, 32'sd0.05925739292298692, 32'sd0.12166834767223667, 32'sd0.028031200088057512, 32'sd-0.08838896145600475, 32'sd-0.05869674587070247, 32'sd0.035385888163351295, 32'sd0.022901535994296184, 32'sd-0.05534788757022325, 32'sd-0.1855752313893801, 32'sd-0.22517777845131445, 32'sd0.03452319556310797, 32'sd0.1328474473490667, 32'sd0.09638932134964043, 32'sd-0.05538040156683013, 32'sd-0.11235090839981685, 32'sd-0.042112159349921414, 32'sd0.10511574503072585, 32'sd0.12869317959899104, 32'sd0.036604966983448395, 32'sd0.04508254094425105, 32'sd0.07708627988998945, 32'sd-0.0758324677503093, 32'sd0.10068500047680333, 32'sd-0.05003499594211311, 32'sd0.07638158916004893, 32'sd-0.06277171728667846, 32'sd-0.09358870993083361, 32'sd0.06298058007967242, 32'sd-0.05204499069103331, 32'sd-0.002996224707277811, 32'sd-0.0736747110359615, 32'sd-0.06449675862591325, 32'sd-0.057985566100453585, 32'sd-0.018682361049955076, 32'sd0.022396132391843907, 32'sd-0.09273379673754682, 32'sd-0.16445186337431028, 32'sd-0.13572278087210934, 32'sd0.14554416954739605, 32'sd0.13437770851849035, 32'sd0.09419757485677291, 32'sd0.04839335459464441, 32'sd0.032791369349601335, 32'sd-0.007237884242623477, 32'sd0.034187111865845714, 32'sd0.11511820232565528, 32'sd0.011057043248198681, 32'sd0.19412802204863217, 32'sd0.10676936061516323, 32'sd-0.06836036549419353, 32'sd0.033142571081768955, 32'sd-0.014121505159968436, 32'sd-0.05132222238229526, 32'sd0.06157669400299866, 32'sd-0.05413639606773643, 32'sd-0.036899462592284174, 32'sd0.07982364418904853, 32'sd-0.1593303683121378, 32'sd-0.07954270626089, 32'sd-0.0970087012679695, 32'sd-0.053787379107647304, 32'sd0.023632858965719452, 32'sd0.02687128737949698, 32'sd-0.13550342432658785, 32'sd-0.14265766236783867, 32'sd-0.15725852662742248, 32'sd-0.022926593279021582, 32'sd0.042539201872512, 32'sd0.08690598596558677, 32'sd0.010654072756454953, 32'sd0.0370022507234741, 32'sd0.06506071182851667, 32'sd-0.0019009137420885477, 32'sd0.06121062837682981, 32'sd-0.0015265437717810876, 32'sd0.15103345516810468, 32'sd-0.08632414678483312, 32'sd0.00391999097212875, 32'sd-0.07066475041514815, 32'sd0.02473509067840241, 32'sd0.06781074381373829, 32'sd0.034260062636003286, 32'sd0.050644916310010606, 32'sd0.025508970965433923, 32'sd-0.09378373904323672, 32'sd-0.024588329223305935, 32'sd-0.053321664669176996, 32'sd0.026727135510688137, 32'sd-0.06272532435997037, 32'sd-0.005816333927045592, 32'sd0.00452545334773913, 32'sd-0.22916880113210103, 32'sd-0.08509571878916634, 32'sd-0.13248756679117743, 32'sd-0.023268185462432003, 32'sd0.04876911720033948, 32'sd0.0679859265719177, 32'sd0.10870158601603161, 32'sd-0.04543138219540208, 32'sd-0.06991860385127843, 32'sd-0.06551848279307694, 32'sd0.012683096698994279, 32'sd-0.001962163265931065, 32'sd0.02469685163298519, 32'sd-0.014535834694877644, 32'sd0.004759053654774026, 32'sd-0.05520143493847461, 32'sd-0.04167769097203962, 32'sd0.020847317350669997, 32'sd-0.016907400651286632, 32'sd-0.031486153963283074, 32'sd-0.025735903287864716, 32'sd0.06738495706984604, 32'sd0.0009130627630305607, 32'sd-0.00543657564534824, 32'sd-0.06177028201333773, 32'sd0.040203271075925306, 32'sd-0.01021175976203973, 32'sd-0.04176379798607472, 32'sd-0.04062953552534904, 32'sd-0.22614309322895448, 32'sd-0.16975443268705878, 32'sd0.049014855445096726, 32'sd0.10174147499063392, 32'sd0.07548263637519008, 32'sd0.04697804888428193, 32'sd0.0016010122962721086, 32'sd0.007900375872501498, 32'sd0.05526934096247311, 32'sd0.007682189265274263, 32'sd0.011529765101761012, 32'sd0.017886508468764283, 32'sd0.1089860303020299, 32'sd-0.052245469681914423, 32'sd-0.062246010559311234, 32'sd-0.04548613377649659, 32'sd-0.006954929143227755, 32'sd-0.015690868604725548, 32'sd0.056528760732828524, 32'sd-0.04808293346505499, 32'sd-0.01431752663852303, 32'sd-0.013190379562556618, 32'sd0.0901733495342257, 32'sd0.04860271452767164, 32'sd0.07214399347477796, 32'sd0.14051181446454933, 32'sd-0.060827459587541564, 32'sd-0.10456570810305177, 32'sd-0.0846067537508728, 32'sd-0.014328122988260928, 32'sd-0.04121851632731625, 32'sd0.06093846475467207, 32'sd-0.04922581149253891, 32'sd0.005457947235559001, 32'sd0.04524050335363098, 32'sd0.06134232088452873, 32'sd0.0672975863570979, 32'sd0.1691117809860209, 32'sd0.24695580369260195, 32'sd0.1285549073169038, 32'sd0.04230520489962292, 32'sd0.05823388350973058, 32'sd-0.09464048162035482, 32'sd-0.04365624858431378, 32'sd-0.032346042559609975, 32'sd-0.015052189698435909, 32'sd0.031783766682837576, 32'sd-0.02617474883293026, 32'sd-0.05877456270537915, 32'sd0.03566318269719964, 32'sd0.11052590848393325, 32'sd0.037644669975534596, 32'sd0.04754729302838102, 32'sd-0.01205371431806623, 32'sd-0.05227533122088372, 32'sd-0.1783456500362696, 32'sd-0.05485046413426121, 32'sd0.04111546263760193, 32'sd-0.013665091621953897, 32'sd-0.007770045376408389, 32'sd-0.0952728017981969, 32'sd0.044517786415240006, 32'sd0.037524703152762275, 32'sd-0.03485739278353851, 32'sd-0.038087221244264176, 32'sd0.10258096192087111, 32'sd0.031114224658849454, 32'sd-0.005198035254157853, 32'sd0.044046718223672975, 32'sd0.031123026201952137, 32'sd-0.17963813192221834, 32'sd0.0324868473485466, 32'sd-0.01964302646473983, 32'sd-0.01845336885149711, 32'sd0.08954938458181924, 32'sd0.024115210299840383, 32'sd0.07261140655909566, 32'sd-0.021424149987420982, 32'sd0.06564647280017757, 32'sd0.08359199536244642, 32'sd0.01548432580860778, 32'sd0.04498842072795442, 32'sd-0.08094601852157932, 32'sd-0.13020406474948623, 32'sd-0.14516159146410945, 32'sd-0.0016613286304480428, 32'sd0.04017727385980194, 32'sd-0.039207013970477315, 32'sd-0.02818500263756933, 32'sd-0.06292281552178303, 32'sd-0.061912629049790585, 32'sd0.007501759972725185, 32'sd-0.0918200146337652, 32'sd0.09638332845003339, 32'sd-0.004266625603168734, 32'sd0.03938762343124969, 32'sd-0.06304529824916796, 32'sd0.08476004693941262, 32'sd0.004895616167160436, 32'sd-0.08348688670968994, 32'sd-0.027284333733844503, 32'sd-1.325626795239733e-122, 32'sd0.11573642258177019, 32'sd0.13856586228311138, 32'sd-0.0345713814653073, 32'sd0.07102938915050744, 32'sd0.12263986083492703, 32'sd-0.03085109865191554, 32'sd0.07933759009472194, 32'sd0.02506351070922249, 32'sd-0.12230432621117905, 32'sd-0.1952831560142364, 32'sd-0.11011001910170662, 32'sd-0.03418692241253418, 32'sd-0.07619705604609191, 32'sd-0.09475153232302784, 32'sd-0.02017978803828327, 32'sd0.029748695776664398, 32'sd0.0543903154695847, 32'sd0.02631592501162028, 32'sd0.002616271001704144, 32'sd0.014283462586167464, 32'sd-0.05668561798451407, 32'sd-0.031733331860100134, 32'sd0.056572974154769216, 32'sd-0.07318227709501816, 32'sd-0.02960221291765102, 32'sd0.02058871174208834, 32'sd-0.018666124620066515, 32'sd0.022193318792553176, 32'sd-0.0002612596734495165, 32'sd0.05333825431023705, 32'sd-0.01340727577678152, 32'sd-0.0028158833238477706, 32'sd0.03141691679529132, 32'sd0.076327100920814, 32'sd0.11335417363401509, 32'sd0.11304550235318846, 32'sd0.11807463650485112, 32'sd0.02342684058992791, 32'sd-0.0736776668143598, 32'sd-0.11047129491346315, 32'sd0.009169119553115456, 32'sd-0.005242004411895847, 32'sd0.019776350614797492, 32'sd-0.01916117258642907, 32'sd-0.00016713651071525293, 32'sd0.012066963152114028, 32'sd-0.05821377021829485, 32'sd-0.009420024319771242, 32'sd-0.017318650795194936, 32'sd0.03583912587929669, 32'sd0.018540447342961064, 32'sd-0.09172374550000274, 32'sd-0.09597696446630156, 32'sd0.01450390708112262, 32'sd-0.010962636929642893, 32'sd0.019814258188656352, 32'sd0.02070228457055902, 32'sd-0.09249607992202527, 32'sd0.03460611709011623, 32'sd0.11696714705073721, 32'sd0.09950153938829485, 32'sd0.1566479384716143, 32'sd0.18707924664149, 32'sd0.11156462828449915, 32'sd0.21488442659877013, 32'sd0.1045091215950018, 32'sd-0.03836773658402113, 32'sd0.14266224506207378, 32'sd0.009040148382232677, 32'sd-0.0015049464148611377, 32'sd0.08581223724003455, 32'sd-0.1525039692030609, 32'sd-0.09760203981982887, 32'sd-0.014190088765454783, 32'sd0.01786509866718124, 32'sd0.0033935387573967735, 32'sd-0.09463622210309751, 32'sd-0.04614427412700318, 32'sd-0.008107933871339741, 32'sd-0.03463910790236547, 32'sd-0.05784179536565699, 32'sd-0.027420910303908464, 32'sd-0.00922391381577349, 32'sd2.3587154562378295e-123, 32'sd0.004662743219861179, 32'sd-0.0027501803082657997, 32'sd0.13130241465097744, 32'sd0.11772516876360162, 32'sd0.00833338266878986, 32'sd0.04638469980645726, 32'sd0.051667304286163084, 32'sd0.13608396785475912, 32'sd0.15979067457747273, 32'sd0.11320833245342797, 32'sd0.053140574067157574, 32'sd0.1054106204330683, 32'sd0.15658021655258114, 32'sd0.0030253136097502507, 32'sd-0.15430694718016297, 32'sd-0.08356296577178114, 32'sd-0.1700870452780607, 32'sd-0.18130035975800912, 32'sd-0.10448056649464664, 32'sd0.00982347733328839, 32'sd0.03259695094135894, 32'sd-0.023918514815816246, 32'sd-0.10539154165404759, 32'sd0.024725598025778745, 32'sd0.08316555768924899, 32'sd-0.008825054059633415, 32'sd0.1213535272348302, 32'sd-0.023396414477322897, 32'sd0.048719556292443573, 32'sd0.004266742774464263, 32'sd0.0380107924706081, 32'sd0.09412670336532065, 32'sd-0.10154836857145723, 32'sd-0.02400921962852324, 32'sd0.07028157233327632, 32'sd0.18352909837096731, 32'sd0.19781092457127347, 32'sd0.19928452025767102, 32'sd0.22145288933815482, 32'sd0.1477302636485659, 32'sd0.07439239192245359, 32'sd0.03473424348539423, 32'sd-0.08256174937553756, 32'sd-0.053932743810897014, 32'sd0.038496928177315634, 32'sd-0.08595713074158105, 32'sd0.0005819067485280353, 32'sd0.03900846129144958, 32'sd-0.010925845696122967, 32'sd-0.1157443471219283, 32'sd-0.11817982627928413, 32'sd-0.08370687954318078, 32'sd-0.03191991606033071, 32'sd0.11332466970385253, 32'sd0.04689999729393315, 32'sd-0.0572445814268601, 32'sd0.027955588988374202, 32'sd0.09585784886812192, 32'sd0.0808188784580506, 32'sd0.08954331850454464, 32'sd0.019418708619222517, 32'sd0.02160167312634573, 32'sd0.013586735208401346, 32'sd0.13505246310091412, 32'sd0.14892504241998028, 32'sd0.2946188357337511, 32'sd0.12662149791613173, 32'sd0.19597626409584223, 32'sd0.19949667981106772, 32'sd0.09197874600072202, 32'sd0.041793480708351184, 32'sd0.09369201861914946, 32'sd-0.0004817099254151298, 32'sd-0.06152411256520906, 32'sd0.05853886738396226, 32'sd0.022979990367685416, 32'sd0.016784728996562626, 32'sd0.0024267157693578364, 32'sd-0.13324024422077632, 32'sd0.027132036877532347, 32'sd-0.004132448249227941, 32'sd0.029476626110025054, 32'sd0.07819825155210212, 32'sd-2.9632033003502465e-119, 32'sd0.04581648505339143, 32'sd0.11884646382464992, 32'sd0.021946638399878756, 32'sd-0.02022769135259381, 32'sd0.04186089942221092, 32'sd0.1077911444136135, 32'sd-0.01900529923041419, 32'sd-0.05423711298142528, 32'sd0.10294889728656346, 32'sd0.18043414024362225, 32'sd0.18147474237698216, 32'sd0.07363513030973731, 32'sd0.06102290931912039, 32'sd0.012446965334068489, 32'sd-0.001416347179115048, 32'sd0.06087624689903733, 32'sd0.08631584285330646, 32'sd-0.05805658561874318, 32'sd-0.22322054854257245, 32'sd-0.15234363626866268, 32'sd-0.003967057834572299, 32'sd-0.05006334788181464, 32'sd-0.009377187421124058, 32'sd-0.0387884895521838, 32'sd-0.050205012129608526, 32'sd-0.04108979535442075, 32'sd-4.4614616919432886e-123, 32'sd-5.517252928250058e-124, 32'sd6.378162499805465e-126, 32'sd0.015528429515743214, 32'sd0.097201449368232, 32'sd0.1087342557654227, 32'sd0.032622973445349146, 32'sd0.09412468939456382, 32'sd0.016777371211653586, 32'sd0.11259492205388211, 32'sd-0.08712035469883886, 32'sd-0.10174367542675132, 32'sd-0.20701767821720035, 32'sd-0.12661729779202965, 32'sd-0.08778712912309611, 32'sd-0.005949260575685503, 32'sd0.05743543210318409, 32'sd-0.093532116289041, 32'sd-0.05980162600338847, 32'sd-0.0816030963021175, 32'sd-0.17570217447226993, 32'sd0.002209611496271959, 32'sd-0.020640640051794522, 32'sd0.012909102962024094, 32'sd-0.031781532528557005, 32'sd0.05305720044953063, 32'sd0.06484899868753011, 32'sd0.08828632703902957, 32'sd-9.562952164207162e-120, 32'sd2.17594825575836e-125, 32'sd-3.237593156644011e-121, 32'sd0.08333765304996715, 32'sd-0.014283409246998446, 32'sd0.022865261210758134, 32'sd-0.024275034944464736, 32'sd-0.13702921063665666, 32'sd-0.12553342658614128, 32'sd0.049816052279545435, 32'sd0.05810362185526958, 32'sd-0.12675538511470272, 32'sd-0.1568237409460808, 32'sd-0.2200816409844836, 32'sd-0.08331330600752579, 32'sd-0.06947118480965982, 32'sd-0.058456800311039704, 32'sd-0.11101965051564243, 32'sd-0.19222158021567332, 32'sd-0.07319161164307518, 32'sd-0.0039541975946392515, 32'sd-0.021826881589536464, 32'sd-0.07010096434384881, 32'sd0.025978460117823704, 32'sd-0.006948879785206838, 32'sd0.09665292408782833, 32'sd-0.0434003571799891, 32'sd0.04493638646426893, 32'sd-2.673468804873837e-116, 32'sd-1.5243101476355195e-115, 32'sd6.612695861665095e-117, 32'sd-1.058787476118311e-124, 32'sd-0.01603247954761493, 32'sd-0.05208174996792416, 32'sd-0.10837140672681671, 32'sd-0.06881952185197297, 32'sd-0.03458190652766648, 32'sd-0.1386765254435737, 32'sd-0.09525883730282994, 32'sd-0.03293138466811066, 32'sd-0.04105801399816786, 32'sd0.060407785036095014, 32'sd-0.06540028380528166, 32'sd-0.045771238279573766, 32'sd-0.11152639752482371, 32'sd-0.09035845623067411, 32'sd-0.03974756973564693, 32'sd-0.0625190281286176, 32'sd-0.019294434179518698, 32'sd-0.08056459507087216, 32'sd0.008941097961224671, 32'sd0.03010163367074711, 32'sd-0.0614221076331407, 32'sd0.021970094077718005, 32'sd0.007597299190884685, 32'sd8.603863813980262e-116, 32'sd3.516664832728111e-122, 32'sd2.46971331274842e-114, 32'sd2.226983218482257e-114, 32'sd-8.619895702809474e-125, 32'sd1.3381028554547085e-122, 32'sd0.0335568964510559, 32'sd-0.037045249767194546, 32'sd-0.019579978226193097, 32'sd0.008921572254268284, 32'sd0.03516016219634829, 32'sd-0.0185113797800851, 32'sd-0.038666765357505954, 32'sd0.008538736819900191, 32'sd0.09096886176598538, 32'sd0.07621623259055521, 32'sd-0.04084624158739669, 32'sd-0.05437500673737072, 32'sd-0.0672946430691555, 32'sd-0.016389547845195616, 32'sd0.01003716734164787, 32'sd0.0471253549120077, 32'sd0.04445994327944448, 32'sd-0.053266174619081216, 32'sd0.00846845708781136, 32'sd-0.01886905337120127, 32'sd2.49375080976168e-124, 32'sd-2.4844384007959134e-124, 32'sd3.042282005144524e-122, 32'sd9.700312225082795e-121},
        '{32'sd3.5627385613225834e-118, 32'sd-1.076319429917413e-124, 32'sd-3.323681153903594e-119, 32'sd7.81629081990073e-123, 32'sd7.28475395662103e-122, 32'sd-1.0045994340322249e-120, 32'sd-1.481487149618548e-126, 32'sd-6.118753601226762e-127, 32'sd4.3012526703827783e-125, 32'sd5.353645889792516e-126, 32'sd1.1615092914463078e-115, 32'sd2.6085333237852938e-124, 32'sd-0.05241465297046943, 32'sd0.05292503655792024, 32'sd-0.013038640546805466, 32'sd0.09476349344031525, 32'sd9.715089908148993e-128, 32'sd2.7107094165134687e-124, 32'sd5.896669835611275e-125, 32'sd-6.949974563564655e-124, 32'sd-9.200423605375604e-125, 32'sd3.801908933809092e-122, 32'sd4.239225800791358e-123, 32'sd-4.0655649732592054e-123, 32'sd-9.291773065690837e-118, 32'sd-1.4908636693548465e-127, 32'sd6.876931488430664e-126, 32'sd-6.794230162995436e-116, 32'sd-1.6452804415278355e-116, 32'sd8.440743822703241e-120, 32'sd-1.1743470161406617e-119, 32'sd-1.3733704512741262e-116, 32'sd-0.008361047905468695, 32'sd0.026953109169445967, 32'sd-0.027527451956528552, 32'sd0.05119662732023329, 32'sd-0.07427026870784384, 32'sd0.0069489614601626355, 32'sd-0.03952398429350133, 32'sd-0.015862601929470938, 32'sd-0.06041862928534155, 32'sd-0.05709718591613809, 32'sd-0.026842126721390767, 32'sd0.06603418219495918, 32'sd-0.022755237393661785, 32'sd0.026737441475293087, 32'sd-0.023758807990368242, 32'sd-0.0004625431672128575, 32'sd0.05144422049157361, 32'sd0.007183108592125106, 32'sd0.000678233770361715, 32'sd0.009494721834903434, 32'sd1.4329742275551226e-119, 32'sd3.1394245666008054e-126, 32'sd2.564777217785e-126, 32'sd-1.0419821295645922e-125, 32'sd2.8245129255755976e-115, 32'sd4.33545658903929e-123, 32'sd0.04933565856026376, 32'sd-0.0020241942106402895, 32'sd-0.06252678215951242, 32'sd-0.009677980951083267, 32'sd-0.05484253912003991, 32'sd0.0025178710664733317, 32'sd-0.021200586587920598, 32'sd-0.10043357895947153, 32'sd-0.020794588731721166, 32'sd0.0005255223579150461, 32'sd-0.09821789442789246, 32'sd-0.11203756553901861, 32'sd-0.08302068133727465, 32'sd-0.029257098733501935, 32'sd-0.03827965448419611, 32'sd-0.0030789976534079323, 32'sd-0.02511707183900635, 32'sd-0.03779099671968939, 32'sd-0.0823044677606959, 32'sd0.03006607039982223, 32'sd0.04797355611807275, 32'sd0.041531267005788866, 32'sd0.062152450898082155, 32'sd-0.03528935984519814, 32'sd-3.599739311176532e-123, 32'sd-1.0127676527990188e-122, 32'sd-4.857147988087191e-124, 32'sd-1.8751244132228958e-120, 32'sd0.03522709355415992, 32'sd-0.0035655723172089322, 32'sd0.03778135836535797, 32'sd0.07632969064156009, 32'sd-0.01858509694490223, 32'sd-0.05627266459134806, 32'sd-0.13401629661542117, 32'sd-0.04232264184533548, 32'sd0.0448538452689725, 32'sd0.04867873994742883, 32'sd0.11494506160651546, 32'sd0.019483152851144173, 32'sd-0.035476895593441034, 32'sd-0.13360823242129438, 32'sd0.029128984179439644, 32'sd-0.027959068187407905, 32'sd-0.16406781850075122, 32'sd-0.22652659882530582, 32'sd-0.14866911388600637, 32'sd-0.06647389431700582, 32'sd-0.0798499235443858, 32'sd-0.05625936017303529, 32'sd0.06702190335578406, 32'sd0.028374023695531488, 32'sd-0.06034928939240105, 32'sd4.617055035980879e-118, 32'sd-3.200739110034914e-118, 32'sd-0.011144470457525072, 32'sd0.010799384001350764, 32'sd0.06918501560277626, 32'sd-0.06108822098591801, 32'sd0.03229029763011796, 32'sd0.0563942568389822, 32'sd0.0811293526143773, 32'sd0.012739600119949, 32'sd0.03796037475944533, 32'sd-0.020546420497546253, 32'sd0.05580573039049859, 32'sd-0.05791537507540756, 32'sd0.01920917573571315, 32'sd0.026457723064476964, 32'sd-0.021170594129175446, 32'sd-0.012152239967132944, 32'sd0.023437930599997915, 32'sd-0.03377765011338545, 32'sd-0.13843576017241357, 32'sd-0.062270742056779564, 32'sd-0.09607336368103943, 32'sd-0.07237598579071274, 32'sd-0.08788315078934077, 32'sd0.036400755661156574, 32'sd-0.025851427545188894, 32'sd-0.02437426684832447, 32'sd0.03600389847707921, 32'sd-1.1360086755089271e-121, 32'sd0.02218578369922138, 32'sd-0.017658491610050682, 32'sd-0.10991921688901726, 32'sd-0.15292572944315155, 32'sd-0.030116794526747755, 32'sd-0.03656139947812318, 32'sd-0.05977038020861685, 32'sd-0.006799666569016539, 32'sd0.1087796004452387, 32'sd0.0654833790245914, 32'sd0.03583087107300974, 32'sd0.0815306859897754, 32'sd-0.005465256231324743, 32'sd0.003973138158122615, 32'sd-0.02365059003078301, 32'sd0.00014819073487848364, 32'sd-0.004496618637905223, 32'sd0.16059923977182541, 32'sd0.05298096708519989, 32'sd-0.06190747233099054, 32'sd-0.06639701832692375, 32'sd-0.003490289537134957, 32'sd-0.019888227815314366, 32'sd-0.02285328070694319, 32'sd-0.04583632562310124, 32'sd0.09189133823083705, 32'sd0.024713990691180875, 32'sd-1.5942951109835808e-115, 32'sd0.0017779980849575165, 32'sd-0.023190352931806952, 32'sd-0.00827124680288653, 32'sd0.02270644717133577, 32'sd-0.09893006106199319, 32'sd-0.07037863629806435, 32'sd0.051513703995198244, 32'sd0.024888868513211922, 32'sd0.04489329342270805, 32'sd0.010975061363838589, 32'sd-0.06332452492366113, 32'sd-0.04731430702311546, 32'sd-0.0025364080516083157, 32'sd0.007300300601650967, 32'sd0.036362530915919185, 32'sd0.12383918579734546, 32'sd0.12681132636150477, 32'sd0.09932536083996873, 32'sd0.09089672362840143, 32'sd-0.021952717584952666, 32'sd0.06099704094916286, 32'sd-0.0009455644401240287, 32'sd-0.03361079352257668, 32'sd-0.058939873690455974, 32'sd0.12201057980230018, 32'sd0.016628905607929345, 32'sd-0.08665171263208518, 32'sd0.009615018910598487, 32'sd0.06178645036674143, 32'sd0.03251021266221615, 32'sd0.00015473906653362806, 32'sd-0.008963088661297958, 32'sd0.04453190007691563, 32'sd-0.0632595708790255, 32'sd-0.04749529493813527, 32'sd0.009091559798361147, 32'sd-0.021544025487275142, 32'sd-0.06948843670774632, 32'sd-0.08944541541943718, 32'sd-0.008414049203370617, 32'sd0.19102648838963537, 32'sd0.11072467495094213, 32'sd0.24351082751008923, 32'sd0.13262236322474458, 32'sd-0.04367090733806316, 32'sd0.10927081635561406, 32'sd-0.03444722903750805, 32'sd0.015412791634391718, 32'sd-0.008303338762774575, 32'sd-0.0030448987493735965, 32'sd-0.03321409541092998, 32'sd0.04428235457809944, 32'sd0.11608594549777872, 32'sd-0.03444528326811005, 32'sd0.0658198490548936, 32'sd0.06340610563793683, 32'sd0.046468000405622406, 32'sd-0.0018859267112065498, 32'sd-0.013088791477240153, 32'sd0.08333889751568378, 32'sd-0.07437861055807447, 32'sd-0.05920709317315331, 32'sd-0.19233392057227158, 32'sd-0.08951841154328821, 32'sd-0.13813455290995058, 32'sd-0.07119793720451587, 32'sd0.06571024773460424, 32'sd0.06762817662780969, 32'sd0.141477128223921, 32'sd0.008030381451200065, 32'sd-0.013275886641842406, 32'sd0.07576643587830723, 32'sd-0.04775550540609002, 32'sd-0.05855429524040902, 32'sd0.08606164045663536, 32'sd-0.052251527293174484, 32'sd0.09245891615091473, 32'sd-0.004927829700791638, 32'sd-0.016150353814228195, 32'sd0.011140037948164063, 32'sd-0.001583831620988691, 32'sd0.1290932789755163, 32'sd-0.0061509578809356945, 32'sd0.010345297025603361, 32'sd0.02307344868561898, 32'sd0.006732664913989652, 32'sd0.038887773981799933, 32'sd-0.08171257729325246, 32'sd-0.03748239595631664, 32'sd-0.14719277657253577, 32'sd-0.12232608991966049, 32'sd-0.056979443292795105, 32'sd-0.013420176466672776, 32'sd-0.048689796163803395, 32'sd0.016416051148344865, 32'sd0.020512148363090826, 32'sd-0.12737928307497384, 32'sd-0.12343908925198709, 32'sd-0.14008015246649563, 32'sd-0.12939027753851168, 32'sd0.0451458048949058, 32'sd-0.13393975376350845, 32'sd0.04990301003099544, 32'sd0.03273471237973236, 32'sd0.029967440193044658, 32'sd0.014013568857203514, 32'sd-0.045400538755209136, 32'sd0.005875400775205761, 32'sd0.00012502249853558542, 32'sd0.07260937370230766, 32'sd0.033285609265461875, 32'sd0.014763806178241851, 32'sd-0.06122763679547837, 32'sd-0.04222992290541268, 32'sd-0.14915471962004928, 32'sd-0.025074699143466585, 32'sd-0.050396895441044885, 32'sd-0.08712938599709902, 32'sd-0.021305090991427626, 32'sd-0.04635654030078691, 32'sd-0.02676526928018895, 32'sd-0.060099269840401065, 32'sd-0.10508585110687944, 32'sd-0.18117180970060273, 32'sd-0.228526986221814, 32'sd-0.22417379699555082, 32'sd-0.18312360903143557, 32'sd0.021172564454901472, 32'sd0.055207556603675156, 32'sd0.04041228854737302, 32'sd-0.02465244758704664, 32'sd0.00019096868313939568, 32'sd0.08585816882407662, 32'sd-0.05402968189889039, 32'sd-0.0323448011312137, 32'sd-0.07453160132195585, 32'sd-0.05263326033062747, 32'sd0.010230202967006182, 32'sd0.06668788601294118, 32'sd0.005877026744115198, 32'sd-0.01756223937318061, 32'sd-0.00021773592490597048, 32'sd0.009827472069822743, 32'sd0.06720937184872115, 32'sd0.08039212573980142, 32'sd0.019342771672651093, 32'sd0.021503174810012002, 32'sd0.14246719150822987, 32'sd0.06695987995921368, 32'sd-0.11685440509540476, 32'sd0.05785499102082235, 32'sd0.011261008220850728, 32'sd-0.10235846363904999, 32'sd0.00832287173069264, 32'sd-0.005937597176167561, 32'sd0.04837677781422307, 32'sd0.08111553190219319, 32'sd-0.013981075783167669, 32'sd0.03060296493670046, 32'sd0.04517488372921984, 32'sd0.02100589082550872, 32'sd0.05324431177080284, 32'sd0.11448843399020411, 32'sd-0.172426126954488, 32'sd-0.06461547270907984, 32'sd-0.015132480460584727, 32'sd0.021774511094507783, 32'sd-0.006982145758394186, 32'sd-0.019501080184323106, 32'sd0.0479275853302608, 32'sd0.10103468477912343, 32'sd0.002335400618094315, 32'sd-0.015101631029650942, 32'sd0.061064621680311536, 32'sd0.03252388038488784, 32'sd0.1845402814941104, 32'sd0.0375638992632353, 32'sd0.04161061663314266, 32'sd0.0354526596013162, 32'sd-0.04152650236653949, 32'sd0.09755516455522338, 32'sd-0.045454949379657876, 32'sd-0.07576460037282624, 32'sd0.07124462724562655, 32'sd0.10149264360941984, 32'sd-0.00882376204729335, 32'sd0.05829475797325072, 32'sd-0.03386293285790314, 32'sd0.09961161975271336, 32'sd0.004673305588822261, 32'sd0.00044896532426226825, 32'sd-0.09319360325905025, 32'sd0.04729489943907045, 32'sd-0.0219182831585944, 32'sd-0.011669063447397416, 32'sd-0.015475095518869247, 32'sd0.009630932933546645, 32'sd-0.04613781227846027, 32'sd-0.02429837847037704, 32'sd0.028884151695317294, 32'sd-0.00033992094181721575, 32'sd0.07233083763552829, 32'sd-0.12085253786429799, 32'sd-0.043457190288043526, 32'sd0.0349300135728839, 32'sd0.039139322779436055, 32'sd0.00765138904316727, 32'sd-0.006923763772558513, 32'sd0.08536770191342988, 32'sd-0.06544440668844836, 32'sd-0.08652285577938498, 32'sd0.02490767893150641, 32'sd-0.025142596858205482, 32'sd-0.009202421096928471, 32'sd-0.1172926372262131, 32'sd0.05284150467634418, 32'sd0.05699612402401933, 32'sd-0.0029778102202956016, 32'sd-0.09547837727565704, 32'sd-0.014257707234132454, 32'sd0.08328539057401489, 32'sd0.07798181453935174, 32'sd0.10104641322192644, 32'sd0.05290725021222022, 32'sd0.05876365601308291, 32'sd0.040089230117821506, 32'sd-0.009568506711758813, 32'sd0.057854663374275264, 32'sd0.09839218550848557, 32'sd0.13906451256876565, 32'sd-0.04337138398043916, 32'sd-0.21233915430991515, 32'sd-0.3001959649458569, 32'sd-0.12906314493595586, 32'sd-0.015356090449394316, 32'sd0.012401387979937417, 32'sd0.03028917992926311, 32'sd-0.058071722304972415, 32'sd-0.054274893449987774, 32'sd-0.07682105132293891, 32'sd-0.12332666399635855, 32'sd-0.1325137162930139, 32'sd-0.10913792598523706, 32'sd0.06458663337295324, 32'sd-0.0068345444679830825, 32'sd-0.18475488301716328, 32'sd-0.10814288366933231, 32'sd-0.03762851197494848, 32'sd-0.07543552126860716, 32'sd-0.051958230606443966, 32'sd0.054232853695401054, 32'sd0.0039672758550089535, 32'sd0.0243297910731258, 32'sd-0.11905828888553055, 32'sd0.002298793344752748, 32'sd-0.03245573504206729, 32'sd0.04861202415987018, 32'sd0.186408181401171, 32'sd0.0859925076425797, 32'sd0.02251542561371347, 32'sd-0.18071993579972032, 32'sd-0.033128333775828314, 32'sd-0.06759226711970169, 32'sd-0.14519100722010392, 32'sd-0.11404636443641317, 32'sd-0.12868690693292145, 32'sd-0.08157545967667935, 32'sd-0.0773596716996728, 32'sd-0.051044779535007835, 32'sd-0.07531254491236859, 32'sd-0.1504497077220074, 32'sd-0.01860762971792103, 32'sd-0.09628187566735892, 32'sd-0.06720370184056317, 32'sd-0.07568398508407087, 32'sd-0.09209912460387189, 32'sd-0.16761095546369256, 32'sd0.05292486346101759, 32'sd-0.025025396528650722, 32'sd0.012376492641567665, 32'sd0.042453311580167255, 32'sd-0.041179383726283804, 32'sd0.01984728686353284, 32'sd0.039398385286100054, 32'sd0.027307086396188417, 32'sd0.04829721149865208, 32'sd0.04943825565973898, 32'sd0.11168401012721643, 32'sd0.0633515228218664, 32'sd0.06914897506807913, 32'sd0.01646825674840219, 32'sd-0.041392702668612745, 32'sd-0.07750831238679394, 32'sd-0.06798190271518409, 32'sd-0.07456042609152695, 32'sd-0.11276033675342136, 32'sd-0.1370753386219598, 32'sd-0.11183824053332313, 32'sd-0.10403221238247172, 32'sd-0.01461728739985311, 32'sd0.03263782214015922, 32'sd-0.07625352795347705, 32'sd-0.11858224681215203, 32'sd-0.1387824938080959, 32'sd-0.056390183962887634, 32'sd-0.03760700573764327, 32'sd-0.020639692197591705, 32'sd1.2329403414011463e-122, 32'sd-0.00536469979492096, 32'sd-0.08311824637382713, 32'sd0.015527628928582443, 32'sd-0.07073267284804455, 32'sd-0.042885434126031595, 32'sd-0.06896198475953436, 32'sd-0.048463137106758654, 32'sd0.07505930713980753, 32'sd0.08266093574270043, 32'sd0.04396833342390774, 32'sd0.04064893325717104, 32'sd0.2109013779697223, 32'sd0.16251936852808288, 32'sd0.07768501637155595, 32'sd0.12039652951426077, 32'sd0.04570739848723518, 32'sd-0.019090467585084214, 32'sd-0.044340903053652306, 32'sd-0.16954039539968557, 32'sd-0.0642502144645164, 32'sd-0.14906744759545118, 32'sd-0.14104573957329303, 32'sd-0.06713680685971063, 32'sd-0.0475387825665137, 32'sd0.12018323893793455, 32'sd-0.03376586085730558, 32'sd0.03368456278925711, 32'sd-0.059258340682518396, 32'sd-0.05764369940637689, 32'sd-0.10312536445896847, 32'sd0.0008910473298172501, 32'sd0.06140368534015334, 32'sd0.037285997352511806, 32'sd0.010955554497163796, 32'sd0.046179675313024096, 32'sd0.020147556723459695, 32'sd0.08940175226559245, 32'sd0.11786406871301257, 32'sd0.006140542287400678, 32'sd0.14490236892157485, 32'sd0.04654424441137707, 32'sd-0.03807630567327579, 32'sd0.10270174108119472, 32'sd-0.017230611289213993, 32'sd-0.09828089109537692, 32'sd-0.06646997848345282, 32'sd0.040594648896228165, 32'sd-0.0010951641051654513, 32'sd-0.03479610875142483, 32'sd-0.07194234635928454, 32'sd0.024876138086627995, 32'sd-0.03868391133308762, 32'sd0.007039720938729517, 32'sd-0.05697841124541753, 32'sd0.055028089767989966, 32'sd0.046312856272626476, 32'sd-0.0892290780982285, 32'sd-0.02833622412501969, 32'sd-0.04471377008164537, 32'sd-0.07811093647855107, 32'sd0.06098562816455807, 32'sd0.04335452699713418, 32'sd0.026152073150974044, 32'sd-0.04055823668706065, 32'sd0.001728968645573602, 32'sd0.006701502607744986, 32'sd-0.07024961225444779, 32'sd0.04007672248043993, 32'sd0.0034578337312062037, 32'sd0.01849779213641443, 32'sd-0.07685198583684576, 32'sd-0.13943522069244996, 32'sd0.026172699341054366, 32'sd-0.01852526274863788, 32'sd0.02325536714569228, 32'sd-0.003829630492508995, 32'sd-0.0010823891757956623, 32'sd-0.06174346027828388, 32'sd-0.018548400569407576, 32'sd0.057078125161098295, 32'sd0.13559328128833942, 32'sd0.010006432206891203, 32'sd-0.09017250830970201, 32'sd1.706908155317735e-125, 32'sd-0.0014710925050534843, 32'sd0.050076897119656065, 32'sd-0.032276440044385596, 32'sd-0.09583077836651521, 32'sd-0.03085226518916393, 32'sd0.07401112808614552, 32'sd-0.056852026588706236, 32'sd-0.08488930634435968, 32'sd0.03318730510886382, 32'sd-0.04423938518651879, 32'sd0.0023261106041642093, 32'sd0.06870251085181422, 32'sd-0.024640426967699698, 32'sd0.05289402715384847, 32'sd0.025473226103859214, 32'sd0.027601911161526393, 32'sd0.1031536508895715, 32'sd0.02461483531426504, 32'sd0.11553701819003696, 32'sd-0.01909994117526356, 32'sd-0.044110417725602716, 32'sd-0.08829082493506345, 32'sd-0.025937486520363186, 32'sd0.05236885991209124, 32'sd0.11051296910965334, 32'sd-0.018501265963977113, 32'sd0.04392271406542741, 32'sd-0.0060027729742761805, 32'sd-0.07230925562666732, 32'sd0.10072565687790799, 32'sd-0.1370579000236875, 32'sd-0.0412640477142713, 32'sd0.028818953034266646, 32'sd0.028860160815215856, 32'sd-0.06264325235998891, 32'sd-0.13888243099949169, 32'sd-0.023177075435073632, 32'sd-0.04408557416331901, 32'sd-0.10136054868977831, 32'sd-0.10388841444181382, 32'sd0.022694763542517826, 32'sd-0.13325971527169364, 32'sd0.05112088100564227, 32'sd0.1393473215969914, 32'sd0.1250563834370209, 32'sd0.04615089089054368, 32'sd0.011316621944539168, 32'sd0.10874960990841932, 32'sd0.11705556934829443, 32'sd0.1473638227465185, 32'sd0.07267825128549459, 32'sd-0.00298145261767441, 32'sd0.13101560679779772, 32'sd0.01405945005103003, 32'sd0.006006487625463794, 32'sd-0.010747192054357193, 32'sd-0.02330109636693115, 32'sd-0.06532137282503965, 32'sd-0.07067217260549927, 32'sd-0.05266602200934097, 32'sd0.028877389845481386, 32'sd0.037824591014113416, 32'sd0.04054419534979562, 32'sd-0.04208722520910164, 32'sd-0.15369894908244483, 32'sd-0.013969947654642679, 32'sd-0.015394425114709034, 32'sd-0.004564011466373501, 32'sd-0.14641701166291413, 32'sd-0.08540503937052965, 32'sd-0.044579287842462796, 32'sd-0.009826956754423759, 32'sd0.08534234099436264, 32'sd0.04250640482371, 32'sd-0.05234970161546544, 32'sd0.0718869329856943, 32'sd0.06509687874014482, 32'sd0.16551250929884037, 32'sd0.05729893596242254, 32'sd0.0816306289105862, 32'sd-0.0032963604223283415, 32'sd-0.013704106627739007, 32'sd-0.007678026366487728, 32'sd-5.186786429567342e-128, 32'sd0.03201354079576668, 32'sd0.016450817407962417, 32'sd-0.12378444164407088, 32'sd-0.06050259623067474, 32'sd0.0072685192382723265, 32'sd-0.0126181336069062, 32'sd-0.0034628898679820116, 32'sd0.0510578185253037, 32'sd-0.06513666202048446, 32'sd-0.0033237128545354666, 32'sd0.081502713673956, 32'sd-0.06336871009571539, 32'sd-0.09029315854043761, 32'sd0.07669631465197882, 32'sd0.05463821284689801, 32'sd0.04868189284895234, 32'sd0.11883895949600319, 32'sd0.1059058674445516, 32'sd-0.005960436089594981, 32'sd-0.028255086196498934, 32'sd0.06540642310692948, 32'sd0.06828986027625365, 32'sd0.05010847866962544, 32'sd-0.1069294700150652, 32'sd0.07945286334908865, 32'sd-0.0723278859460148, 32'sd2.1330911010135245e-126, 32'sd-1.69133177412588e-117, 32'sd2.9175868760800848e-120, 32'sd0.014499825495901357, 32'sd0.007880020737477426, 32'sd-0.0795087685911101, 32'sd-0.10275632154384984, 32'sd-0.009997603957353194, 32'sd0.0026799710914323757, 32'sd0.005462457921643945, 32'sd-0.01345425863369787, 32'sd-0.010890744404047716, 32'sd-0.032177602985571756, 32'sd0.10571690955757833, 32'sd0.18784566432848354, 32'sd0.11075508377242689, 32'sd0.059586921204840056, 32'sd0.13423781238133392, 32'sd0.08931953325574993, 32'sd0.07677969555409256, 32'sd0.07007279961534463, 32'sd-0.03953573291521566, 32'sd0.02675316077777659, 32'sd0.0575020766122778, 32'sd0.0637385810716164, 32'sd-0.018685838475471665, 32'sd0.042930662849459164, 32'sd0.06403337837679829, 32'sd3.3794014846167623e-116, 32'sd-8.836447172108375e-123, 32'sd-5.297107123147212e-116, 32'sd-0.02645999894764383, 32'sd-0.024948281592820053, 32'sd-0.033012872055537656, 32'sd-0.07352785513404266, 32'sd-0.019050576394236463, 32'sd0.05314367505576293, 32'sd0.11088347994411427, 32'sd-0.02993581783585343, 32'sd-0.0022301792211069636, 32'sd0.01841731090667377, 32'sd0.04516281658068985, 32'sd0.16854475289154305, 32'sd-0.041875918436609885, 32'sd0.14948384365308048, 32'sd0.09031534944784207, 32'sd0.17922399802016792, 32'sd0.004374001997152525, 32'sd-0.07244761843303797, 32'sd0.0232451328316494, 32'sd-0.057107114640868026, 32'sd0.09262558408812255, 32'sd0.03695285132787878, 32'sd-0.026341808357338615, 32'sd-0.05871342936069369, 32'sd-0.029396922465605522, 32'sd-3.997289257580743e-126, 32'sd-1.297728119454667e-122, 32'sd8.137143886686402e-117, 32'sd-5.0747231935022696e-126, 32'sd0.03536087414186089, 32'sd0.040950120193349315, 32'sd0.04437971122195005, 32'sd-0.043213278481483396, 32'sd0.06629137796693824, 32'sd0.052373454076208276, 32'sd0.04541211223216003, 32'sd-0.0023322368826131814, 32'sd0.03373795265766292, 32'sd0.16807349676992683, 32'sd0.057828663530189596, 32'sd0.10639334975944849, 32'sd0.13725576613263996, 32'sd-0.01405136191575967, 32'sd0.07266308828995285, 32'sd0.06286093624166697, 32'sd0.02343123907757049, 32'sd0.058422369070772875, 32'sd0.005051063391638866, 32'sd-0.017117112490620617, 32'sd0.1173462343460104, 32'sd0.049359072690066605, 32'sd0.07691348192493808, 32'sd3.6757128864181857e-116, 32'sd-4.275982024464553e-124, 32'sd-1.9116099295947076e-126, 32'sd4.171605689856587e-119, 32'sd2.0033766443717286e-127, 32'sd6.759818656437419e-127, 32'sd-0.0023587500831931943, 32'sd0.08442463705517247, 32'sd-0.026318608472565907, 32'sd0.015344567616782268, 32'sd0.007154122207844463, 32'sd0.014824196886585653, 32'sd-0.0681223579878736, 32'sd0.019464832712068357, 32'sd0.08012298373184616, 32'sd-0.012235892423660716, 32'sd0.038411442169787306, 32'sd0.06512453233507368, 32'sd0.0008490403909594283, 32'sd-0.04097115034907202, 32'sd0.034476612843706324, 32'sd0.013199136021057583, 32'sd-0.038014661833935016, 32'sd0.09430012932880183, 32'sd0.18424045745974996, 32'sd-0.009384747915979421, 32'sd1.0222331383659674e-120, 32'sd2.0369528644707806e-127, 32'sd1.7175854123169825e-125, 32'sd1.676644033600722e-120},
        '{32'sd-6.230952105322304e-119, 32'sd-5.526959720013149e-116, 32'sd-6.277522507094955e-125, 32'sd-7.910848491667046e-124, 32'sd-9.451518041876405e-123, 32'sd-8.011479389490515e-127, 32'sd-2.9003640768782346e-130, 32'sd6.642376083087674e-124, 32'sd-1.0422137159013875e-124, 32'sd1.0490380885368915e-120, 32'sd-2.7422268524448624e-121, 32'sd3.870059302703391e-124, 32'sd0.009815087065373406, 32'sd-0.05374821658025198, 32'sd0.09015509035039419, 32'sd0.03200575558701223, 32'sd-2.147939140670183e-120, 32'sd-4.239327038977327e-118, 32'sd-8.556958900820866e-118, 32'sd1.277667542424291e-127, 32'sd5.48925091860404e-124, 32'sd8.08307980204241e-122, 32'sd5.573472247802717e-118, 32'sd1.0314778921142496e-121, 32'sd-4.7800892211770697e-119, 32'sd1.9067411522348783e-114, 32'sd1.3110569207743449e-122, 32'sd-1.9820525858180504e-121, 32'sd2.486907633223905e-121, 32'sd1.5179401944010226e-124, 32'sd-1.9574724303667745e-126, 32'sd-1.7984709789899622e-123, 32'sd0.030503649173780043, 32'sd-0.0664642977357508, 32'sd-0.0174240437490283, 32'sd0.007576285304194964, 32'sd0.023639803383215134, 32'sd-0.052825512236102615, 32'sd-0.010843950601450138, 32'sd-0.016315038109824022, 32'sd-0.018977183189945897, 32'sd-0.08400081563669363, 32'sd0.04075678498011015, 32'sd0.012196989470934932, 32'sd0.07566625607615418, 32'sd-0.03226619154370901, 32'sd0.002342059521742328, 32'sd-0.07280485343128747, 32'sd0.06671124915213568, 32'sd0.017009534276710092, 32'sd-0.03442336481345723, 32'sd0.0015970885194149364, 32'sd3.2323640481394828e-121, 32'sd-1.0967653363007293e-125, 32'sd1.5164388827477366e-127, 32'sd-1.67894100186939e-126, 32'sd4.7776749882633776e-120, 32'sd-2.840522756992865e-119, 32'sd-0.02485142257166576, 32'sd-0.023891092478389334, 32'sd0.02130690940669095, 32'sd-0.02905124147596137, 32'sd0.011537517136019452, 32'sd-0.0442803768719611, 32'sd-0.0691059338349297, 32'sd-0.05015520633464314, 32'sd-0.052629339226182854, 32'sd-0.09049145356231135, 32'sd-0.1214207528550577, 32'sd-0.011461409903649048, 32'sd0.0459673979368145, 32'sd0.010864433541865712, 32'sd0.029045809450078487, 32'sd0.03344623886380853, 32'sd-0.013638982441187003, 32'sd-0.101302771348608, 32'sd-0.10603046682255625, 32'sd-0.06687541724202299, 32'sd0.050034197744054494, 32'sd0.023565534127450802, 32'sd-0.059769669330654814, 32'sd-0.025666728645365112, 32'sd2.71277362065423e-120, 32'sd-5.50199231988819e-124, 32'sd7.864880528900095e-125, 32'sd1.1948310142444831e-122, 32'sd0.006279093367801738, 32'sd-0.06702797349844042, 32'sd-0.004730165311968622, 32'sd-0.08624012373275963, 32'sd-0.09233283586357985, 32'sd0.015832580718434755, 32'sd-0.08948803616970392, 32'sd-0.1411648068073134, 32'sd-0.1358024925491031, 32'sd-0.07233691145734146, 32'sd-0.12458734926290176, 32'sd-0.14304062359085357, 32'sd-0.09679208530352763, 32'sd-0.048526648335796924, 32'sd0.04856422354361264, 32'sd0.22778506511662627, 32'sd0.18040954314378313, 32'sd0.043801324529345945, 32'sd0.007939722128089103, 32'sd-0.05175130781437812, 32'sd0.03903769018513119, 32'sd-0.03279008703202773, 32'sd-0.028182597697878592, 32'sd0.03964655264413592, 32'sd-0.040967174199824465, 32'sd4.870093107889975e-123, 32'sd-1.0097909722925758e-119, 32'sd0.017170084074274207, 32'sd0.030858484547493695, 32'sd0.06658539034246644, 32'sd-0.0019972500359067683, 32'sd0.013955207180300008, 32'sd-0.07881367310909104, 32'sd0.0025672486872897714, 32'sd-0.12893726191383423, 32'sd-0.017363641755295735, 32'sd0.06472030663695098, 32'sd0.021229178417039543, 32'sd-0.007351231663138817, 32'sd0.029557915893734577, 32'sd-0.07920524240883359, 32'sd-0.06209987717850756, 32'sd-0.016708071083699014, 32'sd0.077769518776913, 32'sd0.19847512521008057, 32'sd0.07252544008304224, 32'sd-0.016418621806982416, 32'sd-0.008294107491507673, 32'sd-0.07457030365534054, 32'sd-0.028346970860658325, 32'sd-0.02078854219038759, 32'sd-0.05178593419224635, 32'sd-0.07423654058347232, 32'sd0.030177780119267087, 32'sd-6.613083322924114e-115, 32'sd0.03170376558804501, 32'sd-0.007899143729192008, 32'sd-0.05611178459530783, 32'sd-0.004261970758980321, 32'sd-0.007877305919463026, 32'sd-0.0406823401375809, 32'sd-0.12738082927777214, 32'sd-0.03224822528743365, 32'sd-0.11259655953929475, 32'sd-0.008979641533751628, 32'sd-0.012235799559398523, 32'sd0.022960402840987472, 32'sd-0.08732970983624944, 32'sd-0.051524551775767126, 32'sd-0.09160688801976227, 32'sd-0.029337108610781298, 32'sd-0.06692764362177325, 32'sd0.15163266134416467, 32'sd0.22451047535907911, 32'sd0.21584199488883307, 32'sd0.0366675267590653, 32'sd-0.047940580361714516, 32'sd-0.08730592135311536, 32'sd0.0008116295563957048, 32'sd-0.07872930075372905, 32'sd-0.08621472402827468, 32'sd-0.02705997115244432, 32'sd-1.2657994032965693e-124, 32'sd0.056808980249365, 32'sd-0.09852997579742515, 32'sd0.05401604418792108, 32'sd-0.0011901717439439436, 32'sd0.03760677031116684, 32'sd-0.04470766621930201, 32'sd-0.09573039211371401, 32'sd-0.11210984447671346, 32'sd-0.008825796084178968, 32'sd-0.023647630080157613, 32'sd0.09241229085348417, 32'sd0.11372083095821041, 32'sd-0.05325284707910989, 32'sd-0.1570024759577854, 32'sd-0.014594716400022932, 32'sd-0.036712307048412225, 32'sd-0.10547440540989078, 32'sd0.006851842198932678, 32'sd0.017781768701326143, 32'sd0.2350343075391153, 32'sd0.02147764207036689, 32'sd-0.08356179119639691, 32'sd0.03063718260762269, 32'sd0.014780070415122132, 32'sd-0.1595003382586489, 32'sd0.021591118048487148, 32'sd-0.03523023146791191, 32'sd0.00748395550711728, 32'sd-0.04595837804087985, 32'sd0.08600291750405145, 32'sd0.0052561609821765885, 32'sd0.07811027647486753, 32'sd-0.035586206658541585, 32'sd0.07676705200669648, 32'sd0.023674613316142807, 32'sd-0.08943292970617758, 32'sd0.05937006370720679, 32'sd0.03471132008022747, 32'sd0.048519980206103173, 32'sd0.08162555990612304, 32'sd-0.12747696101282005, 32'sd-0.06431875289468822, 32'sd-0.05382601627314152, 32'sd0.050490720010402446, 32'sd-0.05011437012691078, 32'sd0.06282715833641611, 32'sd0.0706626415929936, 32'sd0.06268048230060629, 32'sd0.06897528398952367, 32'sd0.034910032416924835, 32'sd-0.019181660055262645, 32'sd0.0007945432289339721, 32'sd-0.204336731548129, 32'sd0.01334061252779939, 32'sd-0.02000806686050324, 32'sd-0.0012431616475812243, 32'sd0.022502789377645816, 32'sd0.08745982663123793, 32'sd0.10137161771633738, 32'sd0.11018580438383115, 32'sd0.04192355964699128, 32'sd0.08381660151974536, 32'sd0.0024955796733982924, 32'sd0.10296752995534773, 32'sd0.05733623293143058, 32'sd-0.02604895703254064, 32'sd-0.07415606448822572, 32'sd-0.11452395902357913, 32'sd-0.14333520188826254, 32'sd-0.12277853500681843, 32'sd-0.15222515380813878, 32'sd-0.05642329248106295, 32'sd-0.04413845116684072, 32'sd0.06860755010580682, 32'sd0.22309927346635366, 32'sd0.09006448808761715, 32'sd0.09281067532007807, 32'sd-0.03274111871289309, 32'sd-0.1084506567832118, 32'sd-0.012409918333530072, 32'sd-0.029106765030116354, 32'sd-0.027042267834130548, 32'sd-0.0937751048268233, 32'sd-0.02791678720807276, 32'sd0.04216379037630127, 32'sd-0.0035067002470128648, 32'sd0.0668576992788932, 32'sd0.08398787909751627, 32'sd0.10745761938880105, 32'sd0.16719300911370977, 32'sd0.10655370912846593, 32'sd0.020820061165697616, 32'sd-0.11337627380114272, 32'sd-0.2569843296626764, 32'sd-0.13269758941242157, 32'sd-0.1736375780466734, 32'sd-0.05804848044772207, 32'sd-0.18535161816513543, 32'sd-0.03264521718486147, 32'sd-0.07435745743672892, 32'sd0.1209103479630839, 32'sd0.2832956644223392, 32'sd0.16119073641305767, 32'sd0.14449202260390837, 32'sd-0.011123532196401708, 32'sd-0.12125018867601874, 32'sd-0.01854517237098055, 32'sd-0.22756650119648952, 32'sd-0.17282472459154152, 32'sd-0.04398904326170851, 32'sd0.041182535149604245, 32'sd0.001748205705956228, 32'sd0.025527976869468914, 32'sd0.02196150110721665, 32'sd0.03378871639910624, 32'sd0.011278038867475651, 32'sd0.04396332677005936, 32'sd0.0850597803648393, 32'sd-0.027814088495040305, 32'sd0.04128466462680471, 32'sd-0.12582220989118564, 32'sd-0.20898880466405884, 32'sd-0.18025613235589846, 32'sd-0.00037579347495892763, 32'sd-0.15402559602178278, 32'sd-0.13827977660856625, 32'sd-0.17312577049065792, 32'sd-0.06539987326375203, 32'sd0.14437462089845407, 32'sd0.30798934397031935, 32'sd0.1257000561767773, 32'sd0.030406995813387346, 32'sd0.0030608689683019586, 32'sd-0.052138009559018456, 32'sd-0.10569197497713104, 32'sd-0.13510240131951845, 32'sd0.0003057483037526398, 32'sd0.008461913990301537, 32'sd0.03284420193510162, 32'sd0.012552380281110628, 32'sd-0.03415032647669396, 32'sd-0.008096706186512804, 32'sd-0.026810225197711993, 32'sd0.013439562317295886, 32'sd0.08615149423887901, 32'sd0.05018638619149366, 32'sd0.05111333767532126, 32'sd-0.14192374108972447, 32'sd-0.19563415113620744, 32'sd0.009482060475988425, 32'sd0.03456589171407036, 32'sd0.025748768495169248, 32'sd-0.16228190198778347, 32'sd-0.10686346357988423, 32'sd-0.0030728608676028435, 32'sd0.06461666384534137, 32'sd0.1215822655436104, 32'sd0.1470895959738886, 32'sd0.03653039251585532, 32'sd-0.12658425570834578, 32'sd-0.16179274880838776, 32'sd-0.2618659534486817, 32'sd-0.1543247206661141, 32'sd-0.02975461651318015, 32'sd0.10476072006024241, 32'sd0.054112367771994435, 32'sd0.04660386334644183, 32'sd0.007776805913822018, 32'sd-0.021707717974178385, 32'sd0.021327225184242335, 32'sd-0.032980392406149896, 32'sd0.00380065023105592, 32'sd0.0463098968712895, 32'sd0.05439301913010857, 32'sd0.08717704669146377, 32'sd-0.11005611350348855, 32'sd-0.13502334471064914, 32'sd0.06729347640677572, 32'sd0.0034661471240399226, 32'sd0.11797057886162442, 32'sd-0.03613681846132863, 32'sd0.036757094423381376, 32'sd-0.04255856743148234, 32'sd0.21253009123878466, 32'sd0.09947891019381731, 32'sd0.14593164029020958, 32'sd-0.10283706293292602, 32'sd-0.1813901195818745, 32'sd-0.1929015402923679, 32'sd-0.21480816701637104, 32'sd-0.059594067008238424, 32'sd-0.09832590277976289, 32'sd-0.023689479994520295, 32'sd-0.03616599084325928, 32'sd0.008375296883898618, 32'sd0.0017002076909358745, 32'sd-0.00479878656172116, 32'sd-0.08598381424666925, 32'sd0.043402238989478294, 32'sd0.08627228335039552, 32'sd-0.033683047777759406, 32'sd0.0036107389926912214, 32'sd0.09964901396571751, 32'sd0.08067154642378624, 32'sd0.007993785352931429, 32'sd0.1852370853395724, 32'sd0.20963947106293718, 32'sd0.05091784328244275, 32'sd0.09128504956263508, 32'sd0.019850067697391862, 32'sd-0.014914893249198086, 32'sd0.11935477112927377, 32'sd0.15253939262667465, 32'sd0.08223562987047907, 32'sd-0.13101570762965584, 32'sd-0.14062962506039775, 32'sd-0.036467397271212, 32'sd-0.0953031113945971, 32'sd-0.06828608236002597, 32'sd-0.04144723922484354, 32'sd-0.031207023147439325, 32'sd0.037097320807460275, 32'sd-0.04802182110181066, 32'sd-0.025323602790313274, 32'sd0.03802745899432727, 32'sd-0.10233927168437741, 32'sd0.0757589999742484, 32'sd-0.056468356039578095, 32'sd0.06538398234637192, 32'sd0.07993434176077496, 32'sd0.110191827652705, 32'sd0.16425537068038007, 32'sd0.193420017985075, 32'sd0.2250009653213976, 32'sd0.13370141798156712, 32'sd0.05919597008608874, 32'sd0.019411182221047953, 32'sd-0.027265385508186857, 32'sd0.07901489180936187, 32'sd0.12923704700943478, 32'sd0.16378819545200698, 32'sd-0.07332648509482384, 32'sd-0.05911733607369902, 32'sd0.07549099432567383, 32'sd0.01707688341291581, 32'sd-0.038567274506237884, 32'sd0.03552454818259394, 32'sd-0.044230092471645735, 32'sd-0.04712627158477395, 32'sd-0.046855496155646034, 32'sd-0.026883705803291195, 32'sd-0.0020044116824902954, 32'sd0.05389816263346141, 32'sd0.01799802620074296, 32'sd0.07457763134380757, 32'sd0.04072149247025328, 32'sd0.019141728506560728, 32'sd0.0068142813970727785, 32'sd0.04083344455092452, 32'sd0.12586439405300762, 32'sd0.1648312334711579, 32'sd0.17576550324200296, 32'sd0.07918754416652256, 32'sd0.13245567306200806, 32'sd0.22823892205913257, 32'sd0.052468535369859626, 32'sd0.0958279584927598, 32'sd-0.04325608049867412, 32'sd0.052066612278535394, 32'sd-0.04187671447771313, 32'sd0.12433865007052071, 32'sd0.09663471325295842, 32'sd-0.028499636151989024, 32'sd0.09228045390091462, 32'sd0.06754256532289046, 32'sd-0.03795367362429748, 32'sd0.015051090586892435, 32'sd-0.10107956927300275, 32'sd0.010571893242310776, 32'sd0.02182844773677162, 32'sd-0.04935028447019454, 32'sd-0.03257485506960187, 32'sd-0.0594857464874438, 32'sd0.10929293713455333, 32'sd-0.0072117062119284705, 32'sd-0.023633429521254936, 32'sd0.020225728486091325, 32'sd0.008979272221120277, 32'sd0.09564178048101002, 32'sd-0.06725041979808943, 32'sd0.09206359043833569, 32'sd0.12846915415041496, 32'sd0.12421959098049455, 32'sd0.06951521471284729, 32'sd0.08890640743409671, 32'sd-0.02820393912613459, 32'sd-0.0017466368339826971, 32'sd0.15509581195151328, 32'sd0.08391494711027406, 32'sd0.06555744077181636, 32'sd0.14926033640889283, 32'sd0.036402791277527165, 32'sd-0.015001753200148595, 32'sd0.10918550411868956, 32'sd0.07312439666718719, 32'sd-0.16455458666101208, 32'sd0.03338165953902582, 32'sd1.567820271621567e-123, 32'sd0.041569761723526714, 32'sd0.013000607693882343, 32'sd-0.00581032447476734, 32'sd0.006435769888651897, 32'sd0.010945313042985254, 32'sd0.057761121096492826, 32'sd0.037218155335492664, 32'sd-0.03664463468657434, 32'sd-0.1715951579030247, 32'sd-0.07796589740254174, 32'sd-0.07050921265401103, 32'sd0.0013745162490286058, 32'sd0.03732024813848072, 32'sd0.05017740233884835, 32'sd0.11119072969163368, 32'sd-0.07479748138805574, 32'sd-0.014324597444329725, 32'sd0.09139963241836616, 32'sd-0.03330838000245779, 32'sd-0.008409558914212197, 32'sd0.10978903271166722, 32'sd0.12804225124551533, 32'sd0.016602685203312238, 32'sd0.06091131701368074, 32'sd-0.013675618556414205, 32'sd-0.04211801655675872, 32'sd-0.039335732025618464, 32'sd0.03904530651118565, 32'sd-0.006787829675212304, 32'sd0.041139693575677136, 32'sd0.11833177369054074, 32'sd0.03056333687691064, 32'sd0.06471642848389521, 32'sd-0.0401720961118402, 32'sd-0.0610223004232705, 32'sd-0.09220335599692832, 32'sd-0.05904745256315546, 32'sd-0.15267261766972934, 32'sd-0.03874959499327928, 32'sd-0.04796803802853104, 32'sd-0.10172007862811003, 32'sd-0.06590771038854866, 32'sd-0.0566253862316552, 32'sd0.04769303834875895, 32'sd0.10651867223224504, 32'sd0.011044011330471533, 32'sd-0.046297428398150646, 32'sd-0.022798077275384375, 32'sd0.020355717475911087, 32'sd0.09269364482376152, 32'sd-0.15524287206422674, 32'sd-0.09956460540409191, 32'sd-0.088341747217428, 32'sd-0.019211597186497828, 32'sd-0.05801996316695539, 32'sd-0.009483207579875572, 32'sd-0.010073876399610061, 32'sd0.07705424869208466, 32'sd0.1425903290844295, 32'sd0.018278048171546095, 32'sd0.15207714583467868, 32'sd0.07085811144362952, 32'sd-0.10074412224800715, 32'sd-0.16632302984871883, 32'sd-0.18674645781453234, 32'sd-0.12741844075935205, 32'sd-0.019070225694153817, 32'sd-0.18509248327472572, 32'sd-0.11165595086106408, 32'sd0.036245381557006844, 32'sd0.001900795486270289, 32'sd0.011593204434911271, 32'sd0.08222786142117691, 32'sd-0.013627200206451875, 32'sd0.015963316817840432, 32'sd-0.03224852623198172, 32'sd0.04042877583806673, 32'sd-0.03407582160787237, 32'sd-0.01929348985782261, 32'sd-0.09427921765833856, 32'sd-0.015877028449434873, 32'sd0.012915610070803494, 32'sd-0.007836508733303207, 32'sd-4.867176078232302e-115, 32'sd0.08385266853880223, 32'sd0.01677149893086561, 32'sd0.04609011330618909, 32'sd-0.011481955789489755, 32'sd0.012331366189980203, 32'sd-0.01530319590518171, 32'sd-0.0855709545099129, 32'sd-0.10790896866482173, 32'sd-0.12126254782209235, 32'sd-0.19352431894943878, 32'sd-0.16083523510134815, 32'sd-0.1622998061148475, 32'sd-0.10816115206660963, 32'sd-0.15624088066841538, 32'sd-0.12842870899904982, 32'sd-0.12309225309180206, 32'sd0.058474445270151276, 32'sd-0.008020304092308226, 32'sd0.0333555057657663, 32'sd0.0030766307807707453, 32'sd-0.02982725193620011, 32'sd0.10609308927729892, 32'sd0.008016934673013936, 32'sd0.0772490880317369, 32'sd-0.06495291965119297, 32'sd0.013739882043571246, 32'sd0.027819218984282686, 32'sd0.039810418957586885, 32'sd-0.021092773504235184, 32'sd0.040235708212587484, 32'sd-0.024402432897838548, 32'sd-0.04863293155687738, 32'sd0.11944882686574722, 32'sd0.07985892052441516, 32'sd0.06199123811851447, 32'sd0.03598625295158385, 32'sd-0.044738630785612216, 32'sd-0.147570219765873, 32'sd0.019813564335844802, 32'sd-0.032161483644763865, 32'sd-0.08132024840192394, 32'sd-0.021946380930604192, 32'sd0.0035435496192606636, 32'sd0.010679707985066095, 32'sd0.04546516197867142, 32'sd0.05871152168146117, 32'sd0.07630376133569797, 32'sd0.013367131578623083, 32'sd0.08247059696327955, 32'sd0.07600341337220212, 32'sd-0.00793885901320215, 32'sd0.13427631265427822, 32'sd0.13242106754611555, 32'sd-0.012365071586585993, 32'sd-0.009024067306248908, 32'sd0.008431831415894465, 32'sd0.06115006844110835, 32'sd0.016885584082359326, 32'sd0.006413979903155545, 32'sd-0.04758476137837506, 32'sd-0.09624361488113833, 32'sd-0.03822955811001334, 32'sd-0.016510332041203214, 32'sd-0.030651722044027493, 32'sd-0.10517654977895168, 32'sd-0.0505386755795864, 32'sd0.08278707107390569, 32'sd-0.024023666691919337, 32'sd0.0445490416338157, 32'sd-0.06664190942565279, 32'sd-0.05357915267702286, 32'sd0.0938228225644677, 32'sd0.13615085018072448, 32'sd0.13168106382007172, 32'sd0.08403232940098462, 32'sd0.10511501383097993, 32'sd0.029854766438630942, 32'sd-0.032334335230562734, 32'sd-0.07352180938117188, 32'sd0.06056872725547918, 32'sd-0.018484947596271152, 32'sd0.0949177420514835, 32'sd0.0006339694751404222, 32'sd1.3552064104202624e-118, 32'sd0.04911079234715557, 32'sd0.02033371340798327, 32'sd0.11230658974531231, 32'sd0.06907549463121057, 32'sd-0.023339717822408578, 32'sd-0.030006022114058156, 32'sd0.0765258181172947, 32'sd-0.025826111681015576, 32'sd-0.029189871688864822, 32'sd0.042741372304091835, 32'sd0.09586084609106796, 32'sd0.00409761369323091, 32'sd0.12000306924752933, 32'sd0.08141633463101855, 32'sd0.011085821798195334, 32'sd0.04038249523551009, 32'sd0.04348304309868624, 32'sd-0.04181821436209539, 32'sd-0.015792400789174942, 32'sd0.05183372048722444, 32'sd0.011335868857876137, 32'sd0.02796491062385562, 32'sd0.021281323202352754, 32'sd0.022005085983839705, 32'sd-0.0503594916601035, 32'sd0.07941611901809797, 32'sd1.7167669734863565e-125, 32'sd4.316438206503977e-119, 32'sd-9.081328169180933e-122, 32'sd0.05678682053140397, 32'sd0.059803516420220006, 32'sd0.042151161761009324, 32'sd-0.06464645218908106, 32'sd0.05067396260309748, 32'sd-0.023305896922628386, 32'sd-0.08244476942789918, 32'sd-0.016696547339799382, 32'sd0.06816113195193588, 32'sd0.04545742206954346, 32'sd-0.029660986891338868, 32'sd-0.04068911452992422, 32'sd0.010646018431932448, 32'sd-0.023893532897299688, 32'sd0.012486661026876551, 32'sd-0.048181520643250965, 32'sd0.0441438235100722, 32'sd-0.0011231876911860965, 32'sd0.03949573208135375, 32'sd0.030960844346683117, 32'sd-0.040214882312125506, 32'sd-0.07844982792775201, 32'sd0.030167371271065255, 32'sd-0.05274797482733554, 32'sd-0.010311433080123314, 32'sd5.35743758591156e-118, 32'sd-2.8637402470742363e-119, 32'sd-6.84040693886542e-126, 32'sd0.027080109080600018, 32'sd-0.07682772175024054, 32'sd-0.021473640920529228, 32'sd-0.015113154169181594, 32'sd0.09996828021816449, 32'sd0.05902526292708046, 32'sd-0.0577142304413684, 32'sd-0.09062686139164645, 32'sd-0.06047471380557497, 32'sd0.0027040579520684112, 32'sd-0.12937837262111979, 32'sd-0.04957664798715876, 32'sd0.0021591189812125685, 32'sd-0.08981945732254044, 32'sd-0.05850627621055924, 32'sd-0.00280314402369307, 32'sd0.15823551835758687, 32'sd0.12809875911483093, 32'sd-0.04023502334161842, 32'sd-0.08803352518928569, 32'sd-0.014757301975216392, 32'sd0.01665835890127834, 32'sd-0.05784945729541889, 32'sd0.016588327663415274, 32'sd-0.02831815317156228, 32'sd3.5523724138987283e-116, 32'sd5.460020940957135e-122, 32'sd3.144046593823616e-119, 32'sd1.8190170022348177e-123, 32'sd-0.03813836035869424, 32'sd0.009616797492747794, 32'sd-0.07745808440808218, 32'sd-0.0329619241154335, 32'sd0.12782061232434147, 32'sd-0.07482070171488474, 32'sd-0.03486483462399421, 32'sd-0.037639984959832375, 32'sd0.03299711973767558, 32'sd0.12846582491119132, 32'sd0.05814412906137768, 32'sd0.03396248647807631, 32'sd0.035050123842412094, 32'sd-0.05148044417864031, 32'sd-0.09087178418914775, 32'sd-0.010406847967627052, 32'sd-0.11207431665523834, 32'sd-0.03289999879300003, 32'sd0.0013982509043002297, 32'sd-0.06002924092481583, 32'sd-0.008314616481910838, 32'sd-0.05097953440512187, 32'sd0.025851689017496127, 32'sd-8.830637099213915e-116, 32'sd-7.443907077477178e-115, 32'sd1.3635217953733825e-121, 32'sd6.526952079399573e-122, 32'sd2.4190412102336626e-115, 32'sd-3.1106152557238726e-117, 32'sd0.019461893648082103, 32'sd0.011194571521196727, 32'sd0.06256240439302277, 32'sd0.003372483533126032, 32'sd-0.03217068089256806, 32'sd-0.06354693293797892, 32'sd0.006903397588939215, 32'sd-0.022456675851209112, 32'sd-0.0109943837533196, 32'sd0.002450637089874245, 32'sd0.008097834310645547, 32'sd0.043367729135622854, 32'sd0.004591656637021053, 32'sd0.044429881269448065, 32'sd0.08213548679322484, 32'sd-0.018115144282478214, 32'sd-0.017425019745532948, 32'sd-0.01299865269262113, 32'sd-0.06143717029173824, 32'sd0.010086472553105052, 32'sd4.160460380535551e-122, 32'sd-1.0603307280382949e-125, 32'sd9.420218051132695e-120, 32'sd-2.71515317005049e-122},
        '{32'sd-1.0782555016947535e-118, 32'sd-7.344131188772271e-116, 32'sd-2.100605663089919e-126, 32'sd-4.086705610801683e-117, 32'sd5.633910790785955e-121, 32'sd4.1958451123511726e-123, 32'sd3.898514258658169e-119, 32'sd3.676832919200718e-116, 32'sd-2.973455275429761e-116, 32'sd2.0743969546869403e-127, 32'sd-1.124678068711404e-127, 32'sd-2.447684581928867e-123, 32'sd-0.06951990762416878, 32'sd0.04866689118756126, 32'sd-0.021316619188607264, 32'sd0.016764456187048662, 32'sd-3.3696328495295927e-125, 32'sd7.998004787503602e-118, 32'sd-3.4572589379035e-122, 32'sd-3.907627472535235e-124, 32'sd2.1883077480264564e-125, 32'sd1.2939224305257032e-118, 32'sd-6.237947890861989e-128, 32'sd1.3527953489521447e-119, 32'sd-1.362902211672622e-123, 32'sd-5.406068841106726e-118, 32'sd7.465430509952406e-118, 32'sd1.3088569741869739e-118, 32'sd-3.4357766474878125e-118, 32'sd1.2573924327736995e-125, 32'sd7.424892799140864e-128, 32'sd-7.209673121913351e-115, 32'sd0.02421522904890127, 32'sd-0.03581800838265752, 32'sd-0.013963480364801243, 32'sd0.034739950734853045, 32'sd-0.023893231137944542, 32'sd0.04276049907148842, 32'sd0.008989090990953545, 32'sd-0.03468506292042971, 32'sd0.00638707997818643, 32'sd-0.016420549538874566, 32'sd-0.029443455545338913, 32'sd0.045763967233956065, 32'sd0.01139166818199959, 32'sd0.0001320934983952259, 32'sd-0.06559509118274379, 32'sd0.02140329651743805, 32'sd-0.04209294761854081, 32'sd-0.04054551129197957, 32'sd-0.0811127506339478, 32'sd0.0252287613722144, 32'sd-1.7742120381394343e-123, 32'sd-1.548518409899346e-127, 32'sd7.565286867824375e-115, 32'sd-3.281835220927456e-125, 32'sd2.6746202856622092e-114, 32'sd-2.0183563927328428e-127, 32'sd0.009355185772222531, 32'sd-0.008950264366429164, 32'sd0.08208555828145278, 32'sd0.012614783450045308, 32'sd-0.05648464557926286, 32'sd-0.011067763389070888, 32'sd-0.016216950950089373, 32'sd-0.0709928949049129, 32'sd0.009253345459671358, 32'sd0.004978847598551877, 32'sd-0.16449569667861155, 32'sd-0.1778054782566247, 32'sd-0.03090576465131526, 32'sd-0.06323412020791402, 32'sd-0.0507392765466349, 32'sd-0.02737959121149412, 32'sd0.07902170279901269, 32'sd0.007642317394291327, 32'sd0.09430257415355099, 32'sd0.07500504585633869, 32'sd0.03475649703073666, 32'sd0.06014600849338596, 32'sd0.009484138778483257, 32'sd0.01294857380119628, 32'sd1.5722220570660485e-125, 32'sd-4.217903842309998e-118, 32'sd-4.945836833981578e-117, 32'sd-1.78716875017493e-117, 32'sd-0.045372186730856606, 32'sd-0.024680173966652952, 32'sd0.03666134779659312, 32'sd0.05924308328401727, 32'sd0.04925757306211585, 32'sd0.022712654417003354, 32'sd0.06864885309139349, 32'sd-0.11013200323314569, 32'sd-0.06407498089492601, 32'sd0.0325303077461497, 32'sd-0.10633262652008305, 32'sd-0.021485080058345086, 32'sd-0.08017791522625549, 32'sd0.02099804318764796, 32'sd0.0920594872582818, 32'sd0.03539611001240683, 32'sd-0.0746783533987844, 32'sd-0.13389445386524762, 32'sd0.010787719036649771, 32'sd-0.11544538566359802, 32'sd-0.10489792236103247, 32'sd-0.007256754507173272, 32'sd0.03527009035343547, 32'sd-0.039578066104916265, 32'sd-0.01681708574072328, 32'sd2.185057940687533e-126, 32'sd2.138802343147013e-118, 32'sd0.015881034350025844, 32'sd0.03013006918191208, 32'sd-0.11754591206942852, 32'sd-0.0507988193300713, 32'sd0.06105140448194873, 32'sd-0.08124232125713512, 32'sd-0.033102168191115944, 32'sd0.05326582169343432, 32'sd0.05409856286692061, 32'sd-0.09843176027933848, 32'sd0.11264513251250798, 32'sd0.050774044172281284, 32'sd0.026458218040459097, 32'sd-0.04091846221977011, 32'sd-0.10625868380515624, 32'sd0.05102176225494609, 32'sd0.0020738556056548673, 32'sd-0.0834992074731193, 32'sd0.00874480404231535, 32'sd-0.010985032434660428, 32'sd0.02861277019896743, 32'sd0.050238180513956766, 32'sd-0.003761434222509624, 32'sd-0.0374264963463957, 32'sd-0.018422551516237673, 32'sd0.03587674693088418, 32'sd-0.026320440491292164, 32'sd-3.8662666785451417e-121, 32'sd-0.020808699165086236, 32'sd-0.04308013220430234, 32'sd-0.015309760365637208, 32'sd-0.007065353371206928, 32'sd0.0726209388249587, 32'sd-0.03604110526612239, 32'sd-0.03660175513484182, 32'sd-0.005808503965790975, 32'sd-0.09041989020790414, 32'sd-0.00903840649694767, 32'sd0.04502828764415582, 32'sd0.13464567343506947, 32'sd-0.05129797405255403, 32'sd-0.005738899044420806, 32'sd0.11638108990829887, 32'sd0.10533274200758524, 32'sd-0.028495270152331317, 32'sd-0.10920160698655734, 32'sd-0.09291848911236435, 32'sd0.02976959839766171, 32'sd0.017558830446291845, 32'sd-0.03322905041354354, 32'sd0.010300980675700653, 32'sd0.033307923630762216, 32'sd0.04068537852764387, 32'sd0.029092595506716248, 32'sd-0.041297117894700704, 32'sd-6.751702011315161e-116, 32'sd0.03959316091801844, 32'sd0.04656599786267415, 32'sd-0.010796200776480983, 32'sd-0.047210339835543014, 32'sd0.09194592527662206, 32'sd0.00378797063566274, 32'sd0.027068191223484136, 32'sd-0.031764337655782016, 32'sd-0.06601376311798599, 32'sd-0.02092318443365422, 32'sd0.12308404835715979, 32'sd0.010072766193989573, 32'sd-0.005035458973461972, 32'sd0.08673048821697557, 32'sd-0.01211727337659977, 32'sd0.023471315064863836, 32'sd-0.036022733422600206, 32'sd-0.1593117597136796, 32'sd-0.17113439979993283, 32'sd-0.039972756699321495, 32'sd0.08360642694596536, 32'sd0.03679180902457917, 32'sd0.11991755783421894, 32'sd-0.07228415908685279, 32'sd-0.15861220767963782, 32'sd0.1026225904773504, 32'sd-0.09487038602741447, 32'sd0.014572974525935041, 32'sd-0.04909835984371544, 32'sd-0.05540991356893485, 32'sd-0.14002719136211234, 32'sd-0.04420316592581426, 32'sd0.09617102130049415, 32'sd-0.07882733309667903, 32'sd0.1136357726983433, 32'sd0.06243411201316228, 32'sd-0.055740818755649596, 32'sd0.0984914930722389, 32'sd0.16699649480464068, 32'sd0.0895674991720293, 32'sd0.09397407518388463, 32'sd-0.042584999196574, 32'sd-0.1849860317084042, 32'sd-0.1106833346372037, 32'sd-0.08015086475506183, 32'sd-0.11272972035709264, 32'sd-0.07156600584142007, 32'sd-0.08154010014035958, 32'sd0.0217864675444687, 32'sd0.031090223849468676, 32'sd-0.04552702256093733, 32'sd0.025228536089758547, 32'sd0.02293482777021299, 32'sd0.005404397955634151, 32'sd-0.10579934420275211, 32'sd0.014395622281298034, 32'sd-0.08039001294175452, 32'sd-0.033252787713289066, 32'sd-0.03717948499760366, 32'sd-0.07561547128903091, 32'sd-0.02120586874186452, 32'sd-0.11971113171690191, 32'sd0.051175682324286965, 32'sd-0.027486582458838938, 32'sd0.014567892013782223, 32'sd0.04687158532332496, 32'sd0.07309294128510911, 32'sd0.19865772804298243, 32'sd0.018842871855851238, 32'sd0.03448065299714715, 32'sd0.014130755585447756, 32'sd-0.12875602238523173, 32'sd-0.03824844404745668, 32'sd-0.02934068973002028, 32'sd-0.0500842871127142, 32'sd0.025749624642079937, 32'sd0.08547285921388617, 32'sd0.09396766225205126, 32'sd0.03325670047024158, 32'sd-0.013225104569515003, 32'sd0.08971990951024622, 32'sd-0.05105999391228201, 32'sd0.00203143472285073, 32'sd0.005273617645865185, 32'sd0.09448758121025501, 32'sd0.10475608188013698, 32'sd-0.00509199217377795, 32'sd0.012703428176440861, 32'sd-0.06261075465281708, 32'sd-0.0013189406870869652, 32'sd-0.05896611842903558, 32'sd0.031436545753403954, 32'sd0.059247661660471185, 32'sd0.09451002375797694, 32'sd0.022710089396476656, 32'sd0.01585364414831471, 32'sd0.1280574460689756, 32'sd-0.014594282194863155, 32'sd-0.11484041148283136, 32'sd0.0230710818283432, 32'sd-0.03354345911465926, 32'sd0.07102316797092445, 32'sd0.021549474217056372, 32'sd0.014801128925465685, 32'sd0.15769590062955677, 32'sd0.10374802017871426, 32'sd0.11028374616540282, 32'sd-0.050660378483325795, 32'sd0.019297073751394063, 32'sd0.07381202145178123, 32'sd-0.04821022397399063, 32'sd0.09692781188885202, 32'sd0.0653822182920871, 32'sd0.1181418938227906, 32'sd0.0679515644085178, 32'sd-0.007388561388201551, 32'sd0.04380618621638058, 32'sd-0.06673525410053668, 32'sd-0.09069650034248437, 32'sd-0.12253827342402833, 32'sd-0.1750349090699134, 32'sd-0.004417423196777138, 32'sd0.033652961054724935, 32'sd0.1432349464525756, 32'sd0.02769979144919134, 32'sd0.05573831751925321, 32'sd-0.05054139352728871, 32'sd-0.09116729955048851, 32'sd-0.028224716478241874, 32'sd0.015189151148108098, 32'sd0.08824816284107016, 32'sd0.12113036571481327, 32'sd0.14884765585051316, 32'sd0.0944098268971086, 32'sd0.14712382813715755, 32'sd0.0468884677915749, 32'sd0.12425819752543822, 32'sd0.0763015696409162, 32'sd0.06211444830702363, 32'sd-0.011159643349056007, 32'sd0.06245640581558412, 32'sd0.05748875285682882, 32'sd0.09291278187030283, 32'sd0.014902175605618224, 32'sd0.04233233104458782, 32'sd0.023327129773458386, 32'sd-0.07970993710518483, 32'sd0.011382960014709433, 32'sd-0.1097431617823711, 32'sd-0.03459298490697496, 32'sd0.0614665276026196, 32'sd0.08340478632827271, 32'sd-0.08948433929333592, 32'sd0.026871534970722935, 32'sd-0.17598938133837894, 32'sd-0.11980275219209993, 32'sd-0.06574279806852784, 32'sd-0.033223271425440064, 32'sd0.06974633622622592, 32'sd0.0622728883091608, 32'sd0.04823724565757727, 32'sd-0.03467816344344911, 32'sd-0.035855364136717444, 32'sd-0.013977472337757157, 32'sd-0.018537137774266146, 32'sd-0.05548680650406084, 32'sd-0.11660583767414258, 32'sd0.012448753377974978, 32'sd0.09242322866316316, 32'sd0.04551492628019557, 32'sd0.0441203244647563, 32'sd0.0991631726514996, 32'sd0.08488448478892713, 32'sd-0.029331318831552124, 32'sd0.0008612820054442514, 32'sd0.008019478172988145, 32'sd-0.0017249138633625698, 32'sd0.1924758793238145, 32'sd0.07926879693994465, 32'sd0.16513790446618837, 32'sd0.0693145947172163, 32'sd-0.030769121603486577, 32'sd-0.11098925538342283, 32'sd-0.016978136415236315, 32'sd0.011871210141419897, 32'sd0.07468362515864377, 32'sd-0.011591811552933736, 32'sd0.06944051823644792, 32'sd0.10860115127501219, 32'sd0.0918100385874253, 32'sd-0.02689025663137479, 32'sd0.04489242213907069, 32'sd0.058357349509900895, 32'sd0.05762494856991403, 32'sd-0.07427076973913116, 32'sd0.06128568540492477, 32'sd0.06117194656393617, 32'sd0.016998763897178564, 32'sd0.03569728692187274, 32'sd0.06302814612789039, 32'sd-0.05950867738542445, 32'sd-0.03059770310264893, 32'sd-0.008276769934370563, 32'sd0.009393239991372046, 32'sd0.18841185637849103, 32'sd0.23590771029774057, 32'sd0.22484953176028818, 32'sd0.17330482429182287, 32'sd0.015830461936087177, 32'sd0.018907575350129633, 32'sd0.05621095023279208, 32'sd-0.02013070776928124, 32'sd0.07814899159006945, 32'sd0.11330659131995248, 32'sd0.020158700029813886, 32'sd0.09560381314702297, 32'sd0.08045286900532544, 32'sd-0.011915507743573122, 32'sd0.003825028788149054, 32'sd-0.03575458448752525, 32'sd-0.02595502549191223, 32'sd-0.05834265387121371, 32'sd0.017535911836671664, 32'sd0.0006786474282317312, 32'sd-0.0050906988912818, 32'sd0.04458250736906067, 32'sd0.022842947427381192, 32'sd-0.027315230785867894, 32'sd0.05542834888115848, 32'sd-0.06035012865299416, 32'sd-0.027370802370343807, 32'sd0.12411956313671527, 32'sd0.21767018354946915, 32'sd0.14621498703822913, 32'sd0.19506331803494742, 32'sd0.21109228622457998, 32'sd0.2093922157856795, 32'sd0.19346991673779604, 32'sd0.18173195608611162, 32'sd0.020846014258414005, 32'sd0.08899594816719344, 32'sd0.046673753673311336, 32'sd-0.001099367644790909, 32'sd0.0008753716642663817, 32'sd0.1565929541194116, 32'sd0.00504345518195419, 32'sd-0.049942926686244955, 32'sd0.031982271632734524, 32'sd-0.00825289179556844, 32'sd-0.04827021230367897, 32'sd0.03794065581691679, 32'sd-0.024021760375880996, 32'sd-0.010853461749954833, 32'sd0.08067033249925686, 32'sd-0.024681279257368745, 32'sd0.030598500430282897, 32'sd0.016306661707939197, 32'sd-0.08774821768890556, 32'sd-0.06294841541832716, 32'sd0.013263083558951711, 32'sd-0.01154971798126306, 32'sd0.16048815229187177, 32'sd0.20113812153841104, 32'sd0.16584799463085428, 32'sd0.17288528293441102, 32'sd0.13318360265013426, 32'sd0.07495556795746497, 32'sd0.08458356869203615, 32'sd0.13320685725668557, 32'sd-0.03628501556653907, 32'sd-0.018469173755465973, 32'sd0.019768848009763362, 32'sd-0.00613174382491245, 32'sd-0.0006289963460761294, 32'sd-0.08810004400085761, 32'sd-0.07582161846282903, 32'sd0.004128551172212175, 32'sd0.04727270796064813, 32'sd0.012030598307728594, 32'sd0.021678343317362455, 32'sd-0.023707790593417006, 32'sd-0.06452286541823259, 32'sd0.05747023877979589, 32'sd0.07866499290028443, 32'sd0.013092468810593045, 32'sd-0.04600036862107571, 32'sd-0.11765757759945748, 32'sd-0.04613434766005665, 32'sd-0.03532858278099251, 32'sd0.0041047393538359575, 32'sd0.03850914356667557, 32'sd0.1663517996809514, 32'sd0.21376623442876014, 32'sd0.05084021721998967, 32'sd0.009221556599216682, 32'sd-0.015887978124921296, 32'sd-0.08474343022516084, 32'sd-0.09787705682791761, 32'sd-0.21816345005662313, 32'sd-0.1059782090084641, 32'sd0.05043548082006151, 32'sd0.03695829444904631, 32'sd-0.06178681410611651, 32'sd0.09313068970657985, 32'sd-0.18288233555182967, 32'sd-0.015519396967103687, 32'sd-0.015894727143775756, 32'sd1.322161417199774e-122, 32'sd0.0808724363927475, 32'sd0.012874496470967325, 32'sd-0.09842578236487166, 32'sd-0.002371127375546923, 32'sd-0.021616873550402427, 32'sd-0.17075269632047427, 32'sd-0.051922251209388905, 32'sd-0.2254571242588566, 32'sd-0.289166171875869, 32'sd-0.35410847174426274, 32'sd-0.17655754754937453, 32'sd-0.09159635389965146, 32'sd0.021304515047195938, 32'sd0.06454791487199749, 32'sd-0.052350807444066914, 32'sd-0.03815510717081631, 32'sd-0.047562155905497734, 32'sd-0.12719486526350496, 32'sd-0.16298030120732898, 32'sd0.02510764874765339, 32'sd0.013415931784442682, 32'sd0.09412121607952938, 32'sd0.02895961752547053, 32'sd0.1259692125631393, 32'sd-0.050087655060276855, 32'sd0.0914761803486046, 32'sd-0.0636878822690096, 32'sd-0.01817997084226162, 32'sd0.07614196115750861, 32'sd-0.08779876495357827, 32'sd-0.010232918438061327, 32'sd-0.05422817410439141, 32'sd-0.13284990737734767, 32'sd-0.11090149492036892, 32'sd-0.14741624241277565, 32'sd-0.15026689155706355, 32'sd-0.3381843020991072, 32'sd-0.3170522239606078, 32'sd-0.15319363454146886, 32'sd-0.10127895772471165, 32'sd-0.006674769793951384, 32'sd-0.031745208946863425, 32'sd-0.11367913949579231, 32'sd-0.018871366134620888, 32'sd-0.15883321585630336, 32'sd-0.1931411731129495, 32'sd-0.22046354770969553, 32'sd-0.13350667639403982, 32'sd0.03680861994130133, 32'sd0.04696155513086808, 32'sd0.013281747045704544, 32'sd-0.04963914229512582, 32'sd0.038897351032065805, 32'sd0.05345749654194791, 32'sd-0.03613639971358887, 32'sd0.009732933662517316, 32'sd0.008272817937063184, 32'sd-0.0025217485167997322, 32'sd0.03024138660626485, 32'sd0.03358266830772625, 32'sd-0.1710103367491599, 32'sd-0.18743147750154857, 32'sd-0.15900094353395858, 32'sd-0.25496493287414623, 32'sd-0.09905535717081974, 32'sd-0.1403184963017549, 32'sd-0.1402844197050135, 32'sd-0.1857041625107605, 32'sd-0.12775453334456754, 32'sd0.006031735856454292, 32'sd0.005078130953720499, 32'sd0.037538674706325166, 32'sd-0.00762782358351598, 32'sd-0.06761277209121562, 32'sd-0.07706170635873678, 32'sd-0.12207963084598297, 32'sd0.10290978876092469, 32'sd0.073211925050937, 32'sd-0.07362353540862909, 32'sd0.013522908613565946, 32'sd0.10481830487649411, 32'sd0.008751625501694912, 32'sd-0.0324972495158736, 32'sd-1.5875226081652678e-115, 32'sd0.0815466544958913, 32'sd0.034433815582475116, 32'sd-0.042607767700815674, 32'sd0.07535636960763063, 32'sd-0.13193807980708175, 32'sd-0.10711343221658269, 32'sd-0.08993562993959614, 32'sd-0.18169886048114622, 32'sd0.07527429684751635, 32'sd0.03628754641663764, 32'sd0.005069292581475334, 32'sd-0.09847658968704982, 32'sd0.031231867781985074, 32'sd0.10370710546488665, 32'sd-0.04118954748401278, 32'sd-0.013303219410730675, 32'sd0.03623935809500583, 32'sd-0.018871646186727375, 32'sd-0.07728096858158194, 32'sd-0.0888715230651524, 32'sd-0.03421807353088545, 32'sd0.11709027581470374, 32'sd0.07807577524191264, 32'sd-0.0650959789209149, 32'sd-0.058303740609689444, 32'sd-0.020394504996208755, 32'sd0.02460326087499044, 32'sd0.056842082302906764, 32'sd0.04385238099069663, 32'sd-0.039972382860727684, 32'sd0.00671173711209911, 32'sd0.11973416755596043, 32'sd-0.08106853844213456, 32'sd0.07744021560745853, 32'sd0.036870818309987334, 32'sd0.12549531533254352, 32'sd-0.002487338695447311, 32'sd0.043261166004414, 32'sd0.06035068195425282, 32'sd0.015814451817992032, 32'sd-0.08795918749202901, 32'sd-0.08805764626255926, 32'sd-0.006924914188930936, 32'sd-0.01111727261227012, 32'sd-0.14222238879762553, 32'sd-0.00830478550374749, 32'sd-0.12961146196586748, 32'sd-0.056174244767698674, 32'sd0.007561227703465725, 32'sd-0.025520252682785394, 32'sd0.042246671026884064, 32'sd0.011932671245884001, 32'sd-0.1018515827968461, 32'sd0.04607834373040811, 32'sd-0.011387287683450778, 32'sd0.03549730943375925, 32'sd0.09162155181778649, 32'sd-0.005961688397101261, 32'sd-0.00036251186455785574, 32'sd0.17373245963341272, 32'sd-0.02654934613436734, 32'sd0.00886657343395435, 32'sd0.12564487105345296, 32'sd0.1114412527821872, 32'sd0.02555078359714682, 32'sd-0.0048516916811781625, 32'sd0.08305476356808474, 32'sd0.10184303153632787, 32'sd0.06950802075907364, 32'sd0.029523470539494202, 32'sd0.002739013839051595, 32'sd-0.07437041322007387, 32'sd-0.008516139737916983, 32'sd0.007626916383793931, 32'sd-0.023520590915655653, 32'sd-0.0248061626279656, 32'sd0.012743548986313028, 32'sd0.05111570919863536, 32'sd0.05684319884924519, 32'sd0.04475006958873601, 32'sd-0.1416346060624707, 32'sd-0.11745860182834013, 32'sd-0.03531122921857621, 32'sd-6.0238472037503545e-124, 32'sd0.04399029417468718, 32'sd-0.04712932172190775, 32'sd-0.06903810458193156, 32'sd-0.04351508639094509, 32'sd0.02298651894443913, 32'sd0.07272263275164416, 32'sd-0.003579428532060625, 32'sd0.15748311879191515, 32'sd0.04413953179351527, 32'sd0.10406811817776626, 32'sd0.03658304570009093, 32'sd0.008249500759800943, 32'sd0.11754060794619223, 32'sd0.09788536043073776, 32'sd-0.12668001821196748, 32'sd-0.03433291323460694, 32'sd0.05412352203836324, 32'sd-0.06530252231208329, 32'sd-0.008267694798992484, 32'sd-0.03904989878228391, 32'sd-0.005556383825377396, 32'sd0.03325071499111365, 32'sd0.02311507594244041, 32'sd-0.013060199867835943, 32'sd0.017352419446318393, 32'sd-0.05342257927038555, 32'sd4.31902126255651e-123, 32'sd-1.275596557060797e-127, 32'sd-1.0537919910110947e-118, 32'sd-0.022762641694015248, 32'sd-0.009420986005900087, 32'sd-0.009989564669245882, 32'sd-0.047675302171230664, 32'sd-0.08977710568342726, 32'sd0.013107233024649447, 32'sd-0.02298497865915461, 32'sd-0.04335964608854593, 32'sd0.012586051280409478, 32'sd0.030711634766014222, 32'sd0.0036923087783244397, 32'sd0.028926752539009233, 32'sd0.16368493128385134, 32'sd-0.10044006791603471, 32'sd-0.1101695909479643, 32'sd-0.05711544850111367, 32'sd-0.029856367087159063, 32'sd0.09009525571121026, 32'sd-0.018091147183523552, 32'sd0.06844141518071653, 32'sd0.005054180850878065, 32'sd-0.06392761130910783, 32'sd0.05781666443748534, 32'sd-0.02288422879129933, 32'sd0.04781429212067923, 32'sd1.8674180076102548e-120, 32'sd-1.3592281179001095e-121, 32'sd-3.0726176123093516e-125, 32'sd-0.0321037322993422, 32'sd0.0016036543148626953, 32'sd0.06411393540367824, 32'sd0.038703958399927865, 32'sd-0.00867758753120524, 32'sd-0.036723707110672535, 32'sd0.06912373783128574, 32'sd-0.014595217263927075, 32'sd-0.05770815493437163, 32'sd0.008007025775148571, 32'sd-0.08077771309737321, 32'sd-0.012200363416657303, 32'sd0.06240632700235573, 32'sd-0.0656436881256149, 32'sd-0.1512440693689137, 32'sd-0.09399296560433797, 32'sd0.09516301069087577, 32'sd0.04694704092986383, 32'sd0.03661002863783795, 32'sd-0.06478022366699267, 32'sd-0.01143886332414356, 32'sd0.03188506145209057, 32'sd0.03186511871024359, 32'sd0.024967482188677902, 32'sd-0.021940039618320483, 32'sd1.732481098717147e-123, 32'sd3.6684237104680075e-116, 32'sd1.1262588521574872e-115, 32'sd-6.740110460227296e-123, 32'sd0.0016055226838064948, 32'sd0.1025023517384206, 32'sd-0.0730099123500156, 32'sd0.05284973809838978, 32'sd-0.006070817424693702, 32'sd0.013899849608560168, 32'sd-0.017147570980445836, 32'sd-0.03356610942115513, 32'sd-0.09966274813586237, 32'sd-0.06393813988266038, 32'sd-0.038544209910151325, 32'sd-0.12469161469745843, 32'sd-0.06681938691419984, 32'sd-0.006592494722805474, 32'sd0.02216285292390117, 32'sd-0.06811711604608431, 32'sd-0.02529359184144447, 32'sd0.016154453946744425, 32'sd-0.04759017326883574, 32'sd-0.09354329452562747, 32'sd0.05526613193780969, 32'sd-0.03350973312851544, 32'sd0.022694518888226236, 32'sd2.555501754661522e-120, 32'sd3.3342725065452456e-121, 32'sd-6.608528064958185e-118, 32'sd7.328560375494092e-122, 32'sd-7.647682486674366e-118, 32'sd-2.7378815063625123e-116, 32'sd-0.030375769876505705, 32'sd-0.00751883654564149, 32'sd-0.041795358440109565, 32'sd-0.03994681873926982, 32'sd0.0583825758824684, 32'sd0.010554284402002399, 32'sd0.0013492517746486396, 32'sd-0.06758703817148667, 32'sd-0.08613133730470927, 32'sd0.0068456437088655975, 32'sd-0.045655720401592687, 32'sd0.020819305549833265, 32'sd-0.053989599941819254, 32'sd-0.07599118447329413, 32'sd-0.029514243575033804, 32'sd-0.026063304068373726, 32'sd0.0448494436459427, 32'sd0.08427705455954765, 32'sd-0.00425709109936775, 32'sd0.0007927934142196992, 32'sd-1.7376116552080973e-125, 32'sd-1.0516869639747648e-124, 32'sd-1.0492357679764088e-120, 32'sd1.0581614417489336e-125},
        '{32'sd1.0244013093544635e-120, 32'sd1.726750300708643e-126, 32'sd-6.626254676884664e-124, 32'sd-4.312551351061593e-125, 32'sd7.342742094629858e-127, 32'sd8.091417366258982e-125, 32'sd3.5761755422419368e-124, 32'sd1.5924414005041436e-127, 32'sd-2.026304754268551e-123, 32'sd1.6096608797795916e-125, 32'sd2.389428773619343e-114, 32'sd1.1849307572425719e-118, 32'sd-0.09087240772878598, 32'sd-0.0352452484222735, 32'sd-0.018116221291571064, 32'sd0.01375086140265373, 32'sd3.9068761780328007e-119, 32'sd3.0011086930658792e-123, 32'sd3.317353338736913e-126, 32'sd1.6404630546815783e-125, 32'sd-4.506093337337643e-125, 32'sd-1.3593708804457275e-125, 32'sd6.201214018789724e-117, 32'sd-2.217337490730259e-122, 32'sd1.6755580814696849e-125, 32'sd5.7190425576431505e-126, 32'sd1.2501512134951792e-118, 32'sd-7.564954206113812e-115, 32'sd3.415106172886138e-122, 32'sd-2.0187937929147382e-115, 32'sd1.7373430297937873e-125, 32'sd1.508146246911598e-115, 32'sd-0.002718263755927313, 32'sd-0.009010901687798589, 32'sd-0.015318952957706366, 32'sd-0.05456697657900364, 32'sd-0.008202019703958754, 32'sd-0.11064529934915568, 32'sd-0.04160361429063699, 32'sd0.019299821812682465, 32'sd-0.011181579792802935, 32'sd-0.01844923972875966, 32'sd-0.0447612869652764, 32'sd0.001271838639906003, 32'sd-0.055232462419067097, 32'sd2.6988173606296032e-05, 32'sd0.02004539627121362, 32'sd0.0687317567758147, 32'sd-0.017465075503125076, 32'sd-0.040687954200821705, 32'sd-0.05649758689936373, 32'sd0.04612380239977836, 32'sd-2.740415778740483e-118, 32'sd8.334075459665152e-120, 32'sd4.425818478171886e-126, 32'sd-3.575646140059644e-114, 32'sd3.291018161040162e-117, 32'sd9.499051584656005e-125, 32'sd-0.008324240266587925, 32'sd-0.018053650448809307, 32'sd-0.018495625597572448, 32'sd-0.05616768636418552, 32'sd-0.05989249857578963, 32'sd0.027191176227726974, 32'sd0.04098617307294869, 32'sd0.038468336150550335, 32'sd-0.08300219510262956, 32'sd-0.0438086626028311, 32'sd0.037706317790122235, 32'sd0.02259227897332166, 32'sd-0.0540108900697477, 32'sd-0.08821064860725458, 32'sd-0.08265452096557441, 32'sd-0.05703596666125697, 32'sd0.07051372286819267, 32'sd-0.057270288988983564, 32'sd-0.01514680442849009, 32'sd0.14046314834457987, 32'sd0.16084519431203928, 32'sd0.10353962805138964, 32'sd0.07245435714153456, 32'sd0.0127565642247706, 32'sd1.9289986232900494e-120, 32'sd2.6365563735378546e-117, 32'sd-1.1440287954656287e-126, 32'sd9.193620035256441e-120, 32'sd0.06276872814023544, 32'sd-0.04676379675316971, 32'sd-0.07839870330454449, 32'sd0.006106246560321095, 32'sd-0.12251038825718291, 32'sd-0.11271925445312028, 32'sd-0.10863362753746013, 32'sd-0.018893661658749217, 32'sd0.07240381915624029, 32'sd0.025066769791873143, 32'sd0.1184589428278246, 32'sd0.020006460002519457, 32'sd-0.07301420084514756, 32'sd-0.0902035373415296, 32'sd-0.028337914512292787, 32'sd0.0065901864054424214, 32'sd0.0627936914907381, 32'sd0.011373320066265034, 32'sd-0.048096713444866344, 32'sd0.08922461994593738, 32'sd-0.032417439664984546, 32'sd0.027510608534133743, 32'sd-0.042393282452403126, 32'sd-0.0570041634950249, 32'sd0.011575666751425778, 32'sd-6.232794284656353e-122, 32'sd-8.393584447407055e-117, 32'sd0.04337730861091776, 32'sd0.003970748647284478, 32'sd-0.06207974835324666, 32'sd0.01892244562775844, 32'sd-0.0230239327959007, 32'sd-0.010908260130496172, 32'sd0.06422404267201531, 32'sd0.03952237891164402, 32'sd-0.04454707044500358, 32'sd0.15532178252014478, 32'sd0.07752086793760862, 32'sd0.1275204777078849, 32'sd0.16167425566744992, 32'sd0.11024084797489231, 32'sd-0.02884339163149356, 32'sd-0.12105448883707778, 32'sd-0.04372778731479217, 32'sd-0.04274611018090129, 32'sd0.0009207507866127009, 32'sd0.08764022970868765, 32'sd0.0893181250318214, 32'sd-0.042252747683995305, 32'sd0.012296478951111696, 32'sd0.01312934465341131, 32'sd0.06360024340479893, 32'sd0.05906361328643448, 32'sd0.07864113939437226, 32'sd-9.761032099748065e-126, 32'sd-0.049793287651417883, 32'sd0.07482387487128164, 32'sd-0.04847351339442657, 32'sd0.04208659594337784, 32'sd0.012251179483755184, 32'sd0.02466418826653166, 32'sd0.09610175645270289, 32'sd0.07981842350949196, 32'sd-0.060836938624982004, 32'sd0.11177310163717512, 32'sd0.1531205179146972, 32'sd0.08986865803020914, 32'sd0.025438659855657655, 32'sd0.011368208541779865, 32'sd0.017066914911963882, 32'sd-0.003313163247099281, 32'sd0.030952175073671956, 32'sd0.056702086247007524, 32'sd-0.01044371095894341, 32'sd0.015020626351759716, 32'sd0.08994347913662905, 32'sd-0.06091719635921431, 32'sd0.10329614438559503, 32'sd-0.10577479875865954, 32'sd0.04616524166196148, 32'sd0.02004143837877358, 32'sd0.02070192091157743, 32'sd-7.719898594109379e-115, 32'sd-0.021913193182466324, 32'sd0.022691016912476988, 32'sd-0.08506238522129775, 32'sd-0.0709501000313436, 32'sd-0.18415410939099494, 32'sd-0.08086801606149069, 32'sd-0.018748681518538823, 32'sd0.031897564087921534, 32'sd0.04076405709813716, 32'sd0.1220180755656161, 32'sd0.0382529731440592, 32'sd-0.015619823647236575, 32'sd-0.11269831637846063, 32'sd0.0054273671801864385, 32'sd-0.026467964102628753, 32'sd0.11023477089725166, 32'sd0.14295826707472756, 32'sd0.03856721701878364, 32'sd-0.11557220442673623, 32'sd-0.17198405715928602, 32'sd-0.07375074776036801, 32'sd-0.006834221085539516, 32'sd0.009669913051386989, 32'sd-0.027701525860033438, 32'sd-0.0612263773339266, 32'sd0.07126529482163656, 32'sd-0.02014983479197034, 32'sd-0.020815750799410247, 32'sd-0.018107860101685455, 32'sd-0.03827045710862058, 32'sd-0.0010782591095291724, 32'sd0.011725628142348548, 32'sd-0.14162950328902352, 32'sd-0.06036907333576096, 32'sd-0.08863459366393533, 32'sd-0.028575032499132215, 32'sd0.0522956137547291, 32'sd0.20750378655232765, 32'sd-0.07130949109487228, 32'sd-0.15099039364411362, 32'sd-0.1666309286138732, 32'sd-0.013509438317293712, 32'sd0.05614289772014349, 32'sd-0.008457392378741765, 32'sd0.08041325244589002, 32'sd-0.11081676924612457, 32'sd-0.22536538922405522, 32'sd-0.08681139074822199, 32'sd-0.09713616940963335, 32'sd0.005952430005107579, 32'sd-0.0828068167294812, 32'sd0.08421673119264403, 32'sd0.09774595962252305, 32'sd-0.01548455733392649, 32'sd0.05198073848344916, 32'sd0.0056874639566306335, 32'sd-0.08206183192081846, 32'sd0.006227485211675832, 32'sd0.018418075880385527, 32'sd0.1199625367500873, 32'sd-0.13213704163964404, 32'sd0.0092224642476649, 32'sd-0.01899510022253625, 32'sd0.03615134922589063, 32'sd0.04791044949433295, 32'sd0.1419933161278699, 32'sd0.10111531375466985, 32'sd-0.06678133451582136, 32'sd-0.08008620025597908, 32'sd-0.05501879493860654, 32'sd0.055765635059182354, 32'sd-0.07861868411531085, 32'sd0.055336768485839766, 32'sd-0.10894762774847772, 32'sd-0.2004169639484351, 32'sd-0.14882968082702225, 32'sd-0.21204250474144684, 32'sd-0.1056253494101532, 32'sd0.03670755165122347, 32'sd0.06565616921384788, 32'sd0.07372411594526396, 32'sd0.01844229351272959, 32'sd-0.023670561881201212, 32'sd0.01305091969660279, 32'sd0.04752219209532359, 32'sd0.01581942948500435, 32'sd0.07523090750012673, 32'sd-0.020746344051744966, 32'sd-0.054529118759318304, 32'sd-0.032071330520064036, 32'sd-0.13394290736445785, 32'sd-0.037298823676537946, 32'sd0.12461568777135751, 32'sd0.08216504121290238, 32'sd-0.07743513845164662, 32'sd-0.05655251833422641, 32'sd-0.1333488625346051, 32'sd-0.005182973683836184, 32'sd-0.029570540043807055, 32'sd-0.16491057201823303, 32'sd-0.11986415788669395, 32'sd-0.1311410364401551, 32'sd-0.09089705301104366, 32'sd-0.09527657613883037, 32'sd-0.11056968878755266, 32'sd0.0925783293989405, 32'sd0.11757204032531841, 32'sd0.04609018794352395, 32'sd0.14388375988217153, 32'sd0.025055429461637538, 32'sd-0.04559702866293913, 32'sd0.005160456197512083, 32'sd0.02847775349973562, 32'sd0.06921134172410094, 32'sd0.04449006894987644, 32'sd0.17233296110294813, 32'sd-0.06641913191563381, 32'sd0.04229184002189378, 32'sd0.08492446315251095, 32'sd0.024350927926829344, 32'sd0.05780180973533434, 32'sd0.06596164863672288, 32'sd-0.044799711005355944, 32'sd-0.111419817172962, 32'sd-0.07246572507438427, 32'sd0.07762795369172616, 32'sd0.06531876019171222, 32'sd-0.056018610769613585, 32'sd-0.04965230332928612, 32'sd0.01089502727856286, 32'sd-0.028493792958785354, 32'sd-0.08061163509696212, 32'sd0.030622406543875935, 32'sd-0.010239966110865674, 32'sd0.023096324782070275, 32'sd0.06086534168731593, 32'sd-0.026008107523390892, 32'sd-0.057365829664941886, 32'sd0.021499103705813802, 32'sd-0.02730014460981098, 32'sd-0.01853829064563536, 32'sd0.12109310791069042, 32'sd0.039093297575568405, 32'sd0.0355145562295762, 32'sd-0.06057123063611631, 32'sd0.02673810810054683, 32'sd0.044308969311285126, 32'sd0.12346798890227348, 32'sd0.12247851492073943, 32'sd-0.06937767897881979, 32'sd0.0035227458444490327, 32'sd-0.052729707315988174, 32'sd-0.08776637029949115, 32'sd0.11676027733381861, 32'sd0.057900762284782636, 32'sd0.04581563723186395, 32'sd-0.0532760648914445, 32'sd-0.07493005852814516, 32'sd0.08290627452506724, 32'sd0.032503124428202815, 32'sd0.07652373833231103, 32'sd-0.04571420822625979, 32'sd0.05353118164004153, 32'sd0.10116893769163318, 32'sd0.08393806107963057, 32'sd0.06930894160508354, 32'sd0.04629367908022905, 32'sd-0.05517102084877263, 32'sd0.07905137107575679, 32'sd0.09125829168368904, 32'sd-0.04657851958404158, 32'sd0.00796555613490666, 32'sd-0.07189021560832695, 32'sd0.04046068860093612, 32'sd0.07672353942502479, 32'sd0.013190829055943784, 32'sd-0.012054683923715764, 32'sd0.12681902811292461, 32'sd0.003499180958257613, 32'sd-0.06917313492710989, 32'sd0.004020761991122975, 32'sd-0.023456272564663882, 32'sd0.008458895825013668, 32'sd0.052180086999557694, 32'sd0.011574624829256513, 32'sd0.043112963092607225, 32'sd0.053038708305292524, 32'sd0.22983847863623638, 32'sd0.22526106668213736, 32'sd0.14898374219107155, 32'sd0.06046921063798978, 32'sd0.09531988264994888, 32'sd0.008288335533398528, 32'sd0.05318053736964243, 32'sd0.024752037966499333, 32'sd-0.0051694961669929585, 32'sd-0.0001411516116634432, 32'sd0.06261470192969354, 32'sd-0.033850525109238, 32'sd-0.07580380702804501, 32'sd-0.048810980652446226, 32'sd-0.10823777793735917, 32'sd-0.008231522275421618, 32'sd0.10134942303819638, 32'sd0.13211763399892212, 32'sd0.03750952691800679, 32'sd0.10602787667627468, 32'sd0.12454737807070404, 32'sd-0.014048248195881402, 32'sd0.0371203922739012, 32'sd0.16644756578011785, 32'sd0.07292926007020796, 32'sd0.0006590065821742474, 32'sd0.08376298014859994, 32'sd0.17143169953910375, 32'sd0.2005423047304551, 32'sd0.20013391340157885, 32'sd0.09006072531811452, 32'sd-0.0005135323937644836, 32'sd0.142166959283964, 32'sd0.03967908926722309, 32'sd0.05819323984516046, 32'sd-0.008614663922717314, 32'sd0.07225575445209154, 32'sd-0.009390064980632796, 32'sd0.054315493423602416, 32'sd0.03873483054692385, 32'sd-0.003030767603779316, 32'sd-0.017021629420665582, 32'sd-0.07134175015120946, 32'sd-0.061361913590413764, 32'sd0.004365570459937265, 32'sd-0.03659611249749403, 32'sd0.007770937431352315, 32'sd0.07046760797137035, 32'sd0.0389750358468797, 32'sd0.016894235698544473, 32'sd0.08396969552296121, 32'sd0.1626049243552589, 32'sd0.1372908469932858, 32'sd-0.034695156154377085, 32'sd0.0722666488401965, 32'sd0.13798664604172947, 32'sd0.1479873489526663, 32'sd0.11833821788377054, 32'sd0.07605014766710333, 32'sd0.01875129654697403, 32'sd0.10875729210747163, 32'sd0.11533834282446821, 32'sd0.017250939582483093, 32'sd0.06277408531553193, 32'sd0.039459589136642735, 32'sd0.05208618397055299, 32'sd0.08572674832816182, 32'sd0.09684790605170666, 32'sd0.03693565183106269, 32'sd0.06266301592510158, 32'sd0.05590173425921421, 32'sd0.05635441492745601, 32'sd-0.07808893537005997, 32'sd-0.06974741648605744, 32'sd0.11787285065947933, 32'sd0.18027458494283163, 32'sd0.08611385256302226, 32'sd0.056188404427287966, 32'sd0.016952109753584976, 32'sd0.01944691043494687, 32'sd-0.04116685565113969, 32'sd-0.022026674166455828, 32'sd0.02951427613348927, 32'sd-0.017216862830968738, 32'sd-0.06721557029123064, 32'sd0.024892953962345133, 32'sd0.06995197057266891, 32'sd-0.05217213233617746, 32'sd-0.11106478255171448, 32'sd0.05426339569095056, 32'sd0.030001051355262584, 32'sd0.07558278299691581, 32'sd0.053670586588843064, 32'sd0.013327524682203292, 32'sd-0.07189309304174428, 32'sd0.08940081843008515, 32'sd-0.10159187194507126, 32'sd-0.008425674250219298, 32'sd0.05200474140471195, 32'sd0.027690589015821374, 32'sd0.02823952297045774, 32'sd0.12338072780091586, 32'sd0.16006925617005674, 32'sd0.03755789407941309, 32'sd-0.04535081151518121, 32'sd0.0714290799240378, 32'sd0.06077630825214467, 32'sd0.019224850428549146, 32'sd-0.11203241859477862, 32'sd-0.016745892859316887, 32'sd0.0009644986410798141, 32'sd-0.057637790366443814, 32'sd-0.013463092056626963, 32'sd0.05627853036273568, 32'sd-0.08231333410885312, 32'sd-0.011090032175149355, 32'sd-0.07876674932797537, 32'sd-0.06533077987855014, 32'sd-0.11702723634827655, 32'sd-0.009681986239086216, 32'sd3.783518330785232e-122, 32'sd0.03383953135179829, 32'sd0.007735658041224521, 32'sd-0.03910027853273446, 32'sd0.032359288848579644, 32'sd-0.00941574605693363, 32'sd0.01897038968837971, 32'sd-0.06711416603694352, 32'sd0.07113288856525271, 32'sd0.11911369384994697, 32'sd0.12745202806707656, 32'sd0.013373024101548154, 32'sd0.035886560317773146, 32'sd0.07196426505251563, 32'sd0.03424755768418318, 32'sd-0.029660373875974283, 32'sd-0.09931061038938803, 32'sd-0.18472116022586232, 32'sd-0.05254706442475321, 32'sd-0.18322473435735287, 32'sd3.569528966007623e-05, 32'sd0.05741083899493559, 32'sd0.003813929633638363, 32'sd0.04595449707069767, 32'sd0.02177171702125512, 32'sd-0.0007456787286279045, 32'sd-0.09645864597192555, 32'sd0.034325099558239786, 32'sd-0.055352257358170405, 32'sd0.03149729630378301, 32'sd0.030641827504374435, 32'sd0.0018533520362695216, 32'sd0.04222188590557037, 32'sd0.15158343638001498, 32'sd0.09684722788713493, 32'sd0.014865164877893924, 32'sd0.042793021986676914, 32'sd0.14980116432678287, 32'sd0.05695413685430264, 32'sd-0.12254797466809672, 32'sd-0.11235978689552739, 32'sd-0.13527777348792552, 32'sd0.02328660574988543, 32'sd-0.11490405563402378, 32'sd-0.1841848332482366, 32'sd-0.03876883942024255, 32'sd-0.11690428009396514, 32'sd-0.20108606619623345, 32'sd-0.06239971119342031, 32'sd0.061256503016779165, 32'sd-0.07543079539111912, 32'sd0.02305775150809456, 32'sd0.050857435880800675, 32'sd0.002638003875361666, 32'sd-0.015822443951702726, 32'sd0.031686511355093136, 32'sd-0.0008603401686708266, 32'sd-0.010912787663483501, 32'sd0.08190122743173282, 32'sd-0.11879368898887249, 32'sd0.08160072191441792, 32'sd0.0010514350939727535, 32'sd0.13810765475912962, 32'sd0.03604692709523002, 32'sd0.16783742307049676, 32'sd0.021117815360596995, 32'sd-0.13721344596802698, 32'sd-0.028571463618367293, 32'sd-0.1513703779922769, 32'sd-0.16004205216819056, 32'sd-0.16896142353914942, 32'sd-0.0969952683326896, 32'sd-0.042299797327521406, 32'sd-0.02627016255240422, 32'sd-0.14331001605158045, 32'sd-0.17790185373160616, 32'sd-0.03721943514268982, 32'sd-0.0035283197798762385, 32'sd0.12825991550577076, 32'sd-0.03463230514280856, 32'sd-0.02237650646001884, 32'sd0.0009458233158643617, 32'sd0.036443263634710385, 32'sd0.06700618987393674, 32'sd1.4434448291292033e-117, 32'sd0.0891763698164166, 32'sd0.10254360577461563, 32'sd-0.03547709084640639, 32'sd0.00013072258862176206, 32'sd0.06846271551557019, 32'sd0.006972677187981583, 32'sd0.19561518820308108, 32'sd0.18346615340524774, 32'sd0.06682659241571103, 32'sd-0.13946414331054613, 32'sd-0.1696760371649836, 32'sd0.011994461787376254, 32'sd-0.10632942312977087, 32'sd-0.012872886795807732, 32'sd0.009892857648079395, 32'sd-0.13985293655039835, 32'sd-0.04809953130949561, 32'sd-0.08175810989476477, 32'sd-0.10440260177202504, 32'sd-0.10306162498541595, 32'sd0.016982525372815086, 32'sd0.11573331737443086, 32'sd-0.03893082857772464, 32'sd-0.13235851587025593, 32'sd-0.09287422069330392, 32'sd0.07890509301879459, 32'sd-0.016274302506076446, 32'sd0.05383942866615187, 32'sd-0.006409664215216947, 32'sd0.0818947860944866, 32'sd-0.029009909538778567, 32'sd-0.10673788637569827, 32'sd-0.01677479171273987, 32'sd0.09392527934068012, 32'sd0.20805157525477766, 32'sd0.03821278163267375, 32'sd0.0010467844871994809, 32'sd0.049881669239913606, 32'sd0.12243660558564938, 32'sd0.10545276810919851, 32'sd0.08462576218044805, 32'sd0.047935445889553355, 32'sd0.002486366728313813, 32'sd-0.07487814872653861, 32'sd0.03414170927730574, 32'sd-0.041837343760621246, 32'sd-0.051516160886696916, 32'sd-0.04179372089878348, 32'sd0.07619600255450007, 32'sd0.05189940795166114, 32'sd-0.0011053017315457497, 32'sd0.04937541653232837, 32'sd-0.09648001219228323, 32'sd0.0900721647886953, 32'sd0.02201828263465004, 32'sd0.05781793075566372, 32'sd0.02565247149439829, 32'sd-0.0420600818930618, 32'sd-0.08716341883136218, 32'sd-0.008402650139443923, 32'sd-0.07380263864485904, 32'sd0.1645568137307216, 32'sd0.1765957191229147, 32'sd0.08600901624034517, 32'sd0.015769280328898724, 32'sd0.1637169817511749, 32'sd-0.02548602416125417, 32'sd0.07066031090769442, 32'sd-0.10246449582965121, 32'sd-0.1403207035265788, 32'sd-0.08074691619009727, 32'sd-0.07318355934472867, 32'sd-0.041133879812101336, 32'sd-0.03177495376873853, 32'sd0.07534773545831389, 32'sd-0.005901875338118713, 32'sd-0.041481485204390656, 32'sd0.027198246124757446, 32'sd0.045250984114804, 32'sd-0.005678109603813631, 32'sd0.05025310765689222, 32'sd0.012774536620936952, 32'sd0.027377969432278354, 32'sd-7.171563902022467e-126, 32'sd0.01945037057528255, 32'sd-0.040204533717011846, 32'sd0.036277418754877076, 32'sd-0.10340690845328326, 32'sd-0.10911489753865268, 32'sd-0.03324611675973368, 32'sd0.08396007629147925, 32'sd0.10797951504152495, 32'sd-0.08399555401753019, 32'sd-0.035575147180632455, 32'sd-0.052048563769864865, 32'sd-0.013220421527282615, 32'sd-0.12367485063495061, 32'sd-0.06547661186169464, 32'sd-0.12883040602746731, 32'sd-0.06537148226234175, 32'sd-0.19357652339579012, 32'sd-0.17484296697962984, 32'sd0.029657751028051797, 32'sd-0.1036891689322618, 32'sd-0.10770873664163921, 32'sd-0.023608949554700366, 32'sd0.04060346496343725, 32'sd0.005880402691186461, 32'sd-0.08300615706493474, 32'sd-0.007317331247184238, 32'sd-8.088152857836704e-122, 32'sd-9.828508485060267e-121, 32'sd-1.2332385343091327e-125, 32'sd0.019856002158029438, 32'sd0.03281915104975253, 32'sd-0.03715091006217844, 32'sd-0.11934037744397434, 32'sd0.01962209707297554, 32'sd0.03783264776062615, 32'sd-0.06711681308759374, 32'sd-0.07135287358362977, 32'sd0.06707062944050894, 32'sd0.011596029498137818, 32'sd0.015527146284015102, 32'sd0.13196509653309835, 32'sd0.030836272363063626, 32'sd-0.032894266477886465, 32'sd-0.03186744803065689, 32'sd0.00018087697214818618, 32'sd-0.015819110968861398, 32'sd-0.013853711784779062, 32'sd-0.06685670077141767, 32'sd-0.06562552323292827, 32'sd0.011388571447500875, 32'sd0.033072489852287015, 32'sd-0.008663254017384228, 32'sd-0.04944392089392978, 32'sd-0.021119041648797864, 32'sd5.767410881567133e-126, 32'sd-1.2580087480075641e-118, 32'sd-4.214955154062599e-124, 32'sd-0.06275980473725462, 32'sd0.05109727803216313, 32'sd0.030006471917601613, 32'sd-0.11869825948477207, 32'sd-0.02946476575676492, 32'sd-0.06381857301860895, 32'sd0.035856249005559664, 32'sd0.06698146106488113, 32'sd-0.0031162288652629338, 32'sd0.0341134134608909, 32'sd-0.019528880885687192, 32'sd0.10533655419960945, 32'sd0.10958946585772432, 32'sd0.1283249801756181, 32'sd0.20209214811380993, 32'sd0.112980381426978, 32'sd0.1661779201582526, 32'sd-0.07395614849361269, 32'sd0.03122052780292579, 32'sd-0.02446135213394253, 32'sd-0.00022139811093636275, 32'sd0.04373849655954054, 32'sd0.06664600469050685, 32'sd-0.014163393465623493, 32'sd0.008062373702813222, 32'sd2.1047839443242237e-117, 32'sd3.467129161311639e-125, 32'sd-3.620264008607455e-116, 32'sd-4.3209655118177364e-117, 32'sd0.020354683784586155, 32'sd-0.007318159811382829, 32'sd-0.027039411227398766, 32'sd-0.1572271571230572, 32'sd-0.040786074721860736, 32'sd0.08952124418206288, 32'sd0.08927344474690616, 32'sd-0.017478339970239135, 32'sd0.12907904843234985, 32'sd0.07683086307843606, 32'sd-0.05485617157306205, 32'sd0.014459135111356531, 32'sd-0.044373191071896634, 32'sd-0.08992258708557349, 32'sd-0.06938733476878242, 32'sd0.003587492636225341, 32'sd-0.08607198270655514, 32'sd0.021541552738575963, 32'sd0.033977243494194044, 32'sd0.005682851219187781, 32'sd-0.07952027496502488, 32'sd-0.03525989904956828, 32'sd-0.02680255443574825, 32'sd2.294445603428952e-126, 32'sd-7.0457891056130535e-121, 32'sd1.3861420484235672e-115, 32'sd5.999677315417494e-124, 32'sd1.196948952147716e-122, 32'sd1.2053329417709365e-115, 32'sd0.019913559602010158, 32'sd0.03366255843227899, 32'sd-0.07796615899306582, 32'sd-0.04302277224283317, 32'sd-0.049277867072365714, 32'sd-0.072851627152359, 32'sd-0.027653284098956874, 32'sd-0.08303024274688997, 32'sd-0.07826338539182172, 32'sd-0.029851398507421988, 32'sd-0.05032808952889674, 32'sd0.07327494093490093, 32'sd0.006668386662656492, 32'sd-0.01022331747033746, 32'sd-0.07137704295667444, 32'sd-0.01852072851743315, 32'sd0.06408522719764634, 32'sd0.08428799047789401, 32'sd-0.05598557516057929, 32'sd-0.002968148413325137, 32'sd-1.4474894842856929e-115, 32'sd1.1823597202913544e-115, 32'sd-2.1503309850275638e-127, 32'sd-2.720861220435011e-121},
        '{32'sd-3.725515961185996e-125, 32'sd-8.456138470404173e-117, 32'sd-1.3922954204989235e-118, 32'sd-3.139898371976817e-123, 32'sd1.356885476942952e-120, 32'sd-5.365204466337017e-118, 32'sd-7.743086118199335e-122, 32'sd-7.279593442120965e-127, 32'sd-4.3111134582631497e-116, 32'sd-7.601421984828835e-122, 32'sd3.610298464464483e-122, 32'sd3.672896465623711e-116, 32'sd0.07084639400544056, 32'sd-0.03205979616765792, 32'sd0.03399783201717839, 32'sd0.06284742695050369, 32'sd-5.690207697650078e-124, 32'sd-1.108498885631233e-121, 32'sd-2.4106379234125644e-119, 32'sd-1.3496466107977487e-118, 32'sd3.636046849123029e-119, 32'sd3.306568846404007e-120, 32'sd3.6657154689637904e-126, 32'sd-4.754351000724126e-118, 32'sd-3.3759191483655358e-124, 32'sd-6.464278883371662e-115, 32'sd1.0491251410339027e-119, 32'sd-1.1628017348596297e-123, 32'sd2.703133692744958e-119, 32'sd3.2499520283038537e-125, 32'sd-3.670005170758107e-116, 32'sd9.910083361911112e-116, 32'sd-0.019469682674429722, 32'sd0.07847425578974301, 32'sd0.047274026692134215, 32'sd0.004557957753462451, 32'sd0.10700887151260069, 32'sd0.025260099763829584, 32'sd0.10495541878241661, 32'sd0.026237240647920483, 32'sd-0.04427689454338849, 32'sd0.008524011476678793, 32'sd-0.020032640702518333, 32'sd0.05990072697818214, 32'sd0.08325200440865281, 32'sd0.049293183580750896, 32'sd0.016947227200888478, 32'sd0.06554082667448027, 32'sd0.027075353350623367, 32'sd0.027800291498784532, 32'sd0.03627468209345991, 32'sd-0.017453357575135314, 32'sd5.23197147119397e-118, 32'sd2.9167117230569426e-119, 32'sd-2.028817194207435e-124, 32'sd2.391862040180392e-126, 32'sd-5.686772641364185e-115, 32'sd-1.1318637677595803e-119, 32'sd0.04028630661755359, 32'sd0.0435366591629368, 32'sd-0.11207189690179212, 32'sd-0.037354431583901136, 32'sd0.0404348165547421, 32'sd0.04751171658311988, 32'sd-0.060551092808676626, 32'sd0.0032743376463704923, 32'sd0.03499714964746045, 32'sd0.029435695313530148, 32'sd0.06159742393769248, 32'sd0.0765943681805525, 32'sd0.000993425440375733, 32'sd0.001689839899168218, 32'sd-0.0184039454208951, 32'sd0.05601888817100042, 32'sd0.04633300319061272, 32'sd0.032841213956833155, 32'sd0.024674336929227426, 32'sd-0.011654357126784197, 32'sd-0.01783697430568708, 32'sd-0.10040880610052105, 32'sd0.1304448777393737, 32'sd0.04735012673564271, 32'sd-1.9169298172684488e-126, 32'sd-4.606644652257e-123, 32'sd1.43474135437909e-118, 32'sd-2.0368412941170683e-125, 32'sd-0.034340029641968514, 32'sd-0.027950967794071132, 32'sd0.027172433128180334, 32'sd-0.1300346779336488, 32'sd-0.02362860483378167, 32'sd-0.0029400973673584466, 32'sd-0.030844669649116092, 32'sd-0.010265360095684916, 32'sd0.08217372184166263, 32'sd0.057479899498747766, 32'sd0.05798646302620581, 32'sd0.043853270576897335, 32'sd0.0613103672149263, 32'sd0.08044003153465079, 32'sd0.04743432492553782, 32'sd-0.0719019434260718, 32'sd-0.027987379102067233, 32'sd-0.028745981533235265, 32'sd-0.11379895339185264, 32'sd-0.10711787952436194, 32'sd-0.0661921957621295, 32'sd-0.07456129796700771, 32'sd-0.0802610574183789, 32'sd-0.005363029707348688, 32'sd-0.016249975868869265, 32'sd-5.362666727921703e-128, 32'sd-3.3099056326072752e-121, 32'sd0.02745828654608485, 32'sd0.07106311435805009, 32'sd0.02249710010533564, 32'sd0.011352673325616482, 32'sd-0.0006494968746825476, 32'sd-0.06043542570882689, 32'sd0.05183119620634359, 32'sd0.08971767464022704, 32'sd0.03133744825193092, 32'sd0.024458678782385522, 32'sd0.034966064024542824, 32'sd0.12320687392427625, 32'sd0.05921097845543319, 32'sd0.16026888211155335, 32'sd0.06357991124829272, 32'sd-0.024352128434094938, 32'sd-0.08303519580651166, 32'sd-0.03876308502108367, 32'sd-0.12412076367976684, 32'sd-0.21425274605381756, 32'sd-0.16406267370195177, 32'sd-0.0010827046750338581, 32'sd-0.11715663369464506, 32'sd-0.046184405458646806, 32'sd0.007739584156230743, 32'sd-0.06144132110779476, 32'sd0.022496287377626985, 32'sd2.9144820604048566e-125, 32'sd0.019963329919421492, 32'sd0.04770589544285027, 32'sd-0.007527897115517502, 32'sd0.011588866290530965, 32'sd0.03625181971150021, 32'sd0.07436298420378457, 32'sd-0.0060121891080011525, 32'sd-0.06887788854097783, 32'sd-0.06741024842030578, 32'sd-0.003344485810699035, 32'sd0.06885369555779151, 32'sd0.08389893069422304, 32'sd0.16139451562318888, 32'sd0.10072697154096726, 32'sd0.10156915419288091, 32'sd-0.009645303833793611, 32'sd-0.09321610638862446, 32'sd0.04273312431227346, 32'sd-0.0003274624045592101, 32'sd-0.056399657085420565, 32'sd-0.24387363353985003, 32'sd-0.09422604996121324, 32'sd-0.030918787951283375, 32'sd-0.0071973069889183, 32'sd-0.013648174329992477, 32'sd-0.011352447741598114, 32'sd0.04749027605861925, 32'sd3.7616908053580906e-122, 32'sd0.018550363071030203, 32'sd-0.018229946102323903, 32'sd-0.07369134513033353, 32'sd-0.00790103685030941, 32'sd0.07370439605314445, 32'sd-0.04309382306127479, 32'sd-0.020585993997707806, 32'sd-0.09704317693183127, 32'sd-0.08754718432569686, 32'sd-0.09408416159601343, 32'sd-0.08258191881286732, 32'sd0.022363016857205056, 32'sd0.021156930741815197, 32'sd0.018726941183132683, 32'sd0.040820508721907255, 32'sd0.009107077618715605, 32'sd0.044180548496456, 32'sd-0.02701995544624001, 32'sd0.013919416123948009, 32'sd-0.043169177809362906, 32'sd-0.08964446020215276, 32'sd-0.04329652727721919, 32'sd-0.08559705179036012, 32'sd-0.052023761188895845, 32'sd0.07652633106020855, 32'sd-0.049433690492254136, 32'sd-0.04636585959690918, 32'sd0.02893947510725047, 32'sd-0.003270054484290504, 32'sd0.038731681123426814, 32'sd0.020858877345336268, 32'sd-0.014608951298566215, 32'sd-0.1002916494597801, 32'sd-0.05833225806773518, 32'sd-0.050470060210161184, 32'sd-0.2044199582306414, 32'sd-0.029777610135201957, 32'sd-0.003056916046900614, 32'sd0.010679944362692519, 32'sd-0.06968204823354804, 32'sd-0.01593677508019104, 32'sd0.11187096466038421, 32'sd0.043024315443268346, 32'sd0.13344514272332872, 32'sd0.057990596297998305, 32'sd-0.0650385241545288, 32'sd0.03371861892017677, 32'sd0.015377055262302847, 32'sd0.024328163985923062, 32'sd-0.08554726954084448, 32'sd-0.07370968716180981, 32'sd-0.10024594629111877, 32'sd0.029418370157490593, 32'sd-0.017491001770530586, 32'sd-0.0205439827151819, 32'sd0.0641279313286742, 32'sd-0.005434552366539367, 32'sd0.08423515091082177, 32'sd0.020476312241306135, 32'sd0.08507746011919728, 32'sd-0.04347033379116887, 32'sd-0.001088686328539042, 32'sd-0.051964524035351, 32'sd-0.10099690482245254, 32'sd-0.08743322802589264, 32'sd-0.02040083821828905, 32'sd-0.18069319768070227, 32'sd-0.10270871159034453, 32'sd-0.07342105018570141, 32'sd0.1309916893632028, 32'sd0.12512418505495862, 32'sd0.09905450319159238, 32'sd0.10042152853950817, 32'sd-0.008986588559890542, 32'sd-0.016892547739382667, 32'sd-0.04088557851514289, 32'sd-0.09170947405507222, 32'sd-0.03285537177136385, 32'sd-0.13230287841410726, 32'sd-0.1108594417239312, 32'sd-0.09210942913775233, 32'sd-0.0667976880676127, 32'sd0.10022647095051399, 32'sd0.11412615623552637, 32'sd0.005796978194628941, 32'sd-0.01664054198471837, 32'sd-0.07489712188252377, 32'sd-0.04062399735313101, 32'sd-0.08344205423005711, 32'sd-0.05073661448842499, 32'sd-0.04313016204822059, 32'sd-0.06534113665619849, 32'sd-0.04995170956232797, 32'sd-0.0075523924335195464, 32'sd-0.13078156718786207, 32'sd-0.06318176689771904, 32'sd0.1025394544022525, 32'sd0.21232281728580218, 32'sd0.16032506664751273, 32'sd0.13580676473596037, 32'sd0.13280401155777616, 32'sd0.0028885335250118807, 32'sd0.05077841649408998, 32'sd-0.14833475413490677, 32'sd-0.1694017232903505, 32'sd-0.027754397681163036, 32'sd-0.09004574576004053, 32'sd-0.054061912636744126, 32'sd-0.07830164851495403, 32'sd-0.05320227504087519, 32'sd0.04589419183696128, 32'sd0.012100302026368786, 32'sd0.07689253345404641, 32'sd0.07653452744394602, 32'sd-0.013627766405120787, 32'sd-0.10583183471398051, 32'sd-0.13232770494863977, 32'sd-0.04302438198719571, 32'sd-0.041145107224332594, 32'sd0.03720946177948038, 32'sd-0.017579205267182964, 32'sd0.01159477409289989, 32'sd-0.09684434590795285, 32'sd0.10166777273075328, 32'sd0.10573660617458763, 32'sd0.20063427819524518, 32'sd0.21390483943672967, 32'sd0.12906649865150963, 32'sd-0.023155311164350337, 32'sd-0.15195141734206516, 32'sd-0.08762122316851068, 32'sd-0.1452791189455832, 32'sd-0.09477520196975812, 32'sd0.036517180376491334, 32'sd-0.12939777130162824, 32'sd-0.07549767477133067, 32'sd0.01070359615777452, 32'sd0.039073835343294006, 32'sd-0.054994584471806725, 32'sd0.05069197100105369, 32'sd0.0027997613163192737, 32'sd0.14966643769773327, 32'sd0.026628191737131494, 32'sd-0.00828484975215431, 32'sd-0.13910872999305546, 32'sd0.018377724277424366, 32'sd0.012861178529441615, 32'sd0.0034791455520978465, 32'sd-0.037401695507925894, 32'sd0.0714754314420163, 32'sd-0.04921144772982988, 32'sd0.13598904045746033, 32'sd0.10790877157763776, 32'sd0.08963822412160344, 32'sd0.1302299571119493, 32'sd0.0793105298493755, 32'sd-0.059754441433111004, 32'sd-0.07600449886016654, 32'sd-0.09501166225424483, 32'sd-0.01817481154569018, 32'sd0.003275241026283438, 32'sd0.019910992744340654, 32'sd-0.017004323719999766, 32'sd-0.0777187468198332, 32'sd0.16612380741765967, 32'sd-0.04457222930866584, 32'sd0.03430294977847847, 32'sd0.04340577917992495, 32'sd0.14417258123336169, 32'sd0.1039134244688121, 32'sd0.008785512255070996, 32'sd-0.09043168681127431, 32'sd-0.1270462912775307, 32'sd0.053439148646635, 32'sd0.008017028613233808, 32'sd0.024258309292261172, 32'sd0.17749089064675283, 32'sd0.16502714335839785, 32'sd-0.051042448388058846, 32'sd0.056266389760566, 32'sd0.14438617250998267, 32'sd0.10957760683235311, 32'sd0.08212561969261384, 32'sd0.052424789288052075, 32'sd-0.04414032047009078, 32'sd-0.07844978025901103, 32'sd-0.15872360313736464, 32'sd-0.08436154606835759, 32'sd-0.11335198232800883, 32'sd-0.12553199078648572, 32'sd-0.015008270777550044, 32'sd-0.0013386617722862754, 32'sd-0.002923558343979369, 32'sd-0.04140914190950452, 32'sd-0.017921969567695106, 32'sd0.00796348278172722, 32'sd0.1476736401941391, 32'sd0.09930935966173145, 32'sd-0.057307553827781126, 32'sd0.05037250577014727, 32'sd-0.09283881996396692, 32'sd0.16511325945254549, 32'sd0.08511242090938216, 32'sd-0.14004713094718915, 32'sd0.01502638883950775, 32'sd0.08448813280981672, 32'sd-0.01836761833835397, 32'sd-0.017000249104254326, 32'sd0.06740522941132429, 32'sd0.14893808871112413, 32'sd0.16360105374906148, 32'sd0.01905008237818889, 32'sd-0.0029927560209935386, 32'sd-0.13355151631060774, 32'sd-0.17795194665382896, 32'sd-0.003040455151801845, 32'sd-0.09972449244569116, 32'sd-0.022071774775442716, 32'sd0.020453158979061952, 32'sd0.050319195814984154, 32'sd0.0336180487485857, 32'sd-0.012646673240970241, 32'sd0.011847017061743216, 32'sd-0.0023028655887890256, 32'sd0.0149686987078171, 32'sd0.07058091620692844, 32'sd-0.013059885955553982, 32'sd0.017284685411721203, 32'sd-0.03526481617732349, 32'sd-0.0034124091996138935, 32'sd-0.024869656351251438, 32'sd-0.10434323394444463, 32'sd-0.11293839908905952, 32'sd-0.13373743709022545, 32'sd-0.16745625826589758, 32'sd0.021658598574627836, 32'sd0.0565428656267214, 32'sd0.2005952335305556, 32'sd0.2082498824144038, 32'sd0.031127443224422027, 32'sd0.04159442537706006, 32'sd-0.11643684458446794, 32'sd-0.08707735884173319, 32'sd0.0513291101198862, 32'sd0.053939992772438196, 32'sd-0.010507560757711417, 32'sd0.1063498697904156, 32'sd0.02192579658888689, 32'sd0.06869561817924355, 32'sd-0.11302924377126353, 32'sd-0.027346919238745892, 32'sd-0.008503066403127271, 32'sd0.09123224104569723, 32'sd0.013535099383928616, 32'sd-0.10607629088731402, 32'sd0.12771422286071485, 32'sd-0.03555732576696909, 32'sd-0.04080391497539016, 32'sd0.0568250412412474, 32'sd-0.02311225693075707, 32'sd-0.03322544502832649, 32'sd-0.15247314683434782, 32'sd-0.12141312130407277, 32'sd-0.11064119123015678, 32'sd0.10178522204238352, 32'sd0.11732112890529024, 32'sd-0.025356766810117514, 32'sd0.07383601912655934, 32'sd-0.09278543022610267, 32'sd-0.10618815070254674, 32'sd-0.08069887766804315, 32'sd-0.06807025307150204, 32'sd-0.055532577001130845, 32'sd0.08257648248930508, 32'sd0.08684915249876617, 32'sd0.06901187204970705, 32'sd0.1175743913808759, 32'sd-0.09199246821762197, 32'sd0.053225079570484515, 32'sd0.024511312777907617, 32'sd0.059016681684003376, 32'sd0.11383275613669586, 32'sd-0.008581596983962788, 32'sd0.08963070147508312, 32'sd-0.0323179544492086, 32'sd0.027180803957793185, 32'sd0.028146064896063673, 32'sd-0.007096839780189167, 32'sd-0.08897550725831804, 32'sd-0.09217862138115293, 32'sd-0.005693611809124529, 32'sd-0.02979963097991496, 32'sd0.13972268486199602, 32'sd0.05012346825407065, 32'sd0.013006155980452055, 32'sd-0.05188811370846579, 32'sd-0.0980462248455565, 32'sd-0.11998682588412614, 32'sd-0.1562261750574609, 32'sd-0.07380409412607936, 32'sd0.01470228149103082, 32'sd-0.056292242322447734, 32'sd0.07835442364056364, 32'sd0.03492759388038397, 32'sd-0.08593096781715576, 32'sd-0.031407916521708296, 32'sd0.0055649765583630694, 32'sd2.052231994547534e-121, 32'sd0.04407483157432473, 32'sd-0.003069182828805907, 32'sd0.04096550288113707, 32'sd0.009237457321905588, 32'sd-0.07550351444284512, 32'sd-0.06073524969784232, 32'sd0.013972375039355243, 32'sd0.008536309898237029, 32'sd-0.012709527948532896, 32'sd-0.07052378737326863, 32'sd-0.020373846724026055, 32'sd-0.12655076110368868, 32'sd0.0810193566040024, 32'sd0.018030606342884194, 32'sd0.0732171370245566, 32'sd-0.09496371118747671, 32'sd-0.08911020925293565, 32'sd-0.0709990498297565, 32'sd-0.01176714562437252, 32'sd-0.028824972740978082, 32'sd0.0009825245135711915, 32'sd0.014194182402414508, 32'sd-0.005509077508867052, 32'sd0.10959235073011486, 32'sd-0.0040481817328829935, 32'sd0.0004895780605051594, 32'sd0.03908839619380231, 32'sd0.041316843309652705, 32'sd0.06536888461417166, 32'sd0.005103125268736083, 32'sd-0.010130418417979513, 32'sd-0.019137179212834574, 32'sd0.03430298944943121, 32'sd0.04905949906984915, 32'sd-0.02704303102637191, 32'sd0.09864347721889226, 32'sd-0.07650214721128776, 32'sd-0.008686583831650382, 32'sd-0.041744697191701166, 32'sd-0.15583112664305399, 32'sd0.02327236228804815, 32'sd0.04401576630823485, 32'sd-0.006889174934554064, 32'sd-0.055140601649637015, 32'sd-0.06605774757545976, 32'sd-0.09130600911462369, 32'sd-0.02197796668787819, 32'sd-9.981355150924478e-05, 32'sd-0.01712479705921353, 32'sd-0.04610963743814147, 32'sd0.09609363256180585, 32'sd0.026377719555082873, 32'sd0.07541385492407507, 32'sd0.05777819474486432, 32'sd0.08454290983494268, 32'sd0.029976136528027535, 32'sd0.010726836960191432, 32'sd0.037382632395034934, 32'sd-0.09534977087729349, 32'sd0.06347037294976211, 32'sd0.03411453203629904, 32'sd-0.059206136222476995, 32'sd0.08934994602916098, 32'sd-0.036561096817730024, 32'sd-0.07186421743921717, 32'sd-0.10138509619875576, 32'sd-0.1412336670213105, 32'sd-0.08636137982256635, 32'sd0.013417043021980091, 32'sd0.0491132680617682, 32'sd-0.02382746007520728, 32'sd-0.09151227841620944, 32'sd-0.05887643584237612, 32'sd-0.10005226035333888, 32'sd0.07210563477716142, 32'sd0.028201074494456274, 32'sd-0.10096770427907385, 32'sd-0.018654562749479617, 32'sd-0.04647273493767462, 32'sd-0.09757828826052606, 32'sd0.09762666305001268, 32'sd0.024700254125679506, 32'sd0.0855600518092656, 32'sd-5.548782960325235e-115, 32'sd-0.0031306531973804507, 32'sd0.019089916274630924, 32'sd-0.06617395463929183, 32'sd-0.039007849800190106, 32'sd-0.04482334658160689, 32'sd-0.09150000427882372, 32'sd-0.008851300982265591, 32'sd0.0416961779548877, 32'sd-0.00686744706423006, 32'sd-0.07868092885559111, 32'sd-0.05893483779155429, 32'sd0.08347242957278814, 32'sd-0.09402069173180932, 32'sd-0.012245430270266396, 32'sd-0.10227302508699106, 32'sd-0.03339391163199779, 32'sd0.01163917346729417, 32'sd-0.03355924681602915, 32'sd0.028145931684970052, 32'sd-0.07122112763162132, 32'sd-0.018493836000959187, 32'sd-0.0890256372493259, 32'sd0.09362759725921244, 32'sd0.04583911413307105, 32'sd0.11987613496377612, 32'sd0.05914289008626518, 32'sd0.09202022573236662, 32'sd0.08474815913205815, 32'sd0.04201517981169491, 32'sd0.06661958052182701, 32'sd0.04737774275635338, 32'sd-0.03490072537435832, 32'sd-0.1494376574089963, 32'sd-0.10471037373935493, 32'sd-0.042102622272094235, 32'sd0.0671165311973035, 32'sd0.0319054838498244, 32'sd0.034461323740938556, 32'sd-0.027748477673579207, 32'sd0.020015303521890626, 32'sd-0.029883648221222733, 32'sd-0.10604052975242732, 32'sd-0.032521117263011705, 32'sd-0.0856039205481272, 32'sd-0.12021428380378904, 32'sd-0.10179158190691348, 32'sd0.005105959291797165, 32'sd0.03781167968242879, 32'sd-0.007351036743853612, 32'sd0.012493879989018375, 32'sd-0.08836764936155057, 32'sd-0.0022585818766838557, 32'sd0.07410403970762228, 32'sd0.04518836184099516, 32'sd0.05022161658079717, 32'sd0.03808315758094835, 32'sd0.0739111595077792, 32'sd0.03424660305247824, 32'sd0.11549198722712319, 32'sd0.06911576732135812, 32'sd-0.07282723349701073, 32'sd0.008850416506880131, 32'sd0.017839027399486646, 32'sd-0.03222147110641266, 32'sd0.12701629066000944, 32'sd0.12976499905287406, 32'sd0.035728293648297334, 32'sd-0.13050651529071702, 32'sd-0.050022178151746734, 32'sd0.1380296768358412, 32'sd0.07166434376551639, 32'sd-0.0698770577958233, 32'sd0.05105972570541361, 32'sd0.09205618132435367, 32'sd0.08248161897084962, 32'sd0.10981579857663032, 32'sd-0.0031005993573938804, 32'sd-0.053020942352044347, 32'sd-0.08536893302463407, 32'sd-0.07395081201956025, 32'sd0.027179481296282147, 32'sd0.052466965051375825, 32'sd0.08874985387331688, 32'sd1.0445965819378089e-129, 32'sd0.044780323374417605, 32'sd-0.019910297912088024, 32'sd0.1061302358525461, 32'sd0.00663450025433212, 32'sd-0.0906648658690996, 32'sd-0.0980545575161843, 32'sd0.008192661353953707, 32'sd0.005217592110664277, 32'sd0.04924424352146451, 32'sd0.08024063440814105, 32'sd0.004678544661569605, 32'sd0.015127248207193973, 32'sd0.031907895515111556, 32'sd-0.009110302236184139, 32'sd0.12989761786214132, 32'sd-0.06845376158062576, 32'sd0.09246364629511765, 32'sd0.021936857546064725, 32'sd0.0364995456048951, 32'sd0.0711144789753559, 32'sd0.031963957119820065, 32'sd0.03395270944984306, 32'sd0.061344954938344035, 32'sd-0.09541362770633319, 32'sd-0.038434134882350146, 32'sd0.0011529514425070437, 32'sd-5.663240626414552e-115, 32'sd-4.274614403923456e-124, 32'sd-1.0888364313235557e-121, 32'sd-0.0013483026479624352, 32'sd0.13349705514409566, 32'sd0.0671705984700944, 32'sd-0.04051928618720217, 32'sd-0.09382515247795026, 32'sd-0.09154341472444306, 32'sd0.0605288649158765, 32'sd0.03347338348588816, 32'sd-0.02702173315591232, 32'sd-0.04873496919560861, 32'sd-0.06511509718832145, 32'sd-0.0926018035073845, 32'sd0.005326967950569084, 32'sd0.07619780818172024, 32'sd-0.02483796957225965, 32'sd0.006691768064586548, 32'sd0.0099585146780046, 32'sd0.08964570525530695, 32'sd0.02652446087137943, 32'sd0.0835502920376015, 32'sd0.06486556764644393, 32'sd-0.01832958690711997, 32'sd0.07235825469072357, 32'sd-0.05657055080993216, 32'sd0.05098959870838959, 32'sd-3.8394127335098425e-126, 32'sd9.972595092719248e-121, 32'sd5.662139740370278e-115, 32'sd0.04625669094068984, 32'sd-0.08490640511927346, 32'sd0.04245412126027835, 32'sd-0.000760668949523787, 32'sd-0.12294682036940219, 32'sd0.04753096812989359, 32'sd0.22215211826032122, 32'sd0.11557004223543564, 32'sd0.09888034213593358, 32'sd-0.053792593565039015, 32'sd-0.10859260461233647, 32'sd0.01239305955993248, 32'sd0.05169814255986389, 32'sd0.09150628868581907, 32'sd-0.0420269980741053, 32'sd0.05096308231116161, 32'sd-0.16317845798112293, 32'sd-0.06826161049057462, 32'sd0.12623071076735656, 32'sd-0.015841958333688937, 32'sd-0.046172755700135695, 32'sd0.014511645220515765, 32'sd0.02316409743874883, 32'sd-0.025108882894951858, 32'sd0.012461138556394335, 32'sd-5.112045251092539e-118, 32'sd-2.0580426482436628e-127, 32'sd-1.4538249911123424e-123, 32'sd3.446741214745486e-122, 32'sd0.045019616879836556, 32'sd-0.08284228619486493, 32'sd0.028813055113349726, 32'sd0.11452017148469043, 32'sd0.1643529983274812, 32'sd0.0946378482061372, 32'sd0.05566095149910141, 32'sd0.024884840544208624, 32'sd0.07568719398221607, 32'sd0.08254801973943064, 32'sd-0.13417098661003984, 32'sd-0.0006941374459623189, 32'sd-0.02942372598868464, 32'sd-0.03279253868843756, 32'sd0.006754307448008663, 32'sd-0.10050965202793147, 32'sd-0.006774558692683525, 32'sd0.03702987488498998, 32'sd0.07047803441278244, 32'sd-0.10745776344623356, 32'sd0.06361043196390612, 32'sd0.12069392845503302, 32'sd0.08581204511851598, 32'sd3.91547857396974e-118, 32'sd7.178803667556192e-125, 32'sd-4.799624338805072e-119, 32'sd1.6667749783386833e-123, 32'sd4.084009796729969e-120, 32'sd-1.1043672861938833e-123, 32'sd0.11662022342087133, 32'sd-0.039408540759028575, 32'sd0.06762284550391447, 32'sd-0.05806045812418366, 32'sd0.03200936284810424, 32'sd0.027153122326748397, 32'sd0.004619144611358237, 32'sd0.04605798770844695, 32'sd0.0967435062503442, 32'sd0.02177374611218349, 32'sd0.026459114297694517, 32'sd0.03420827511040459, 32'sd0.05563400610320767, 32'sd0.035494832161986525, 32'sd-0.0018831738350525375, 32'sd0.044866158377357634, 32'sd-0.03013019829169501, 32'sd0.15289661040929764, 32'sd0.10635094512791553, 32'sd0.1522722721104565, 32'sd8.402376880389533e-117, 32'sd6.588744592260437e-124, 32'sd-9.304818848197883e-118, 32'sd3.2174242387884416e-120},
        '{32'sd3.555791769714238e-119, 32'sd3.0740430831524685e-125, 32'sd-4.2132438443931075e-122, 32'sd3.7997981244083694e-120, 32'sd3.750438115274762e-124, 32'sd1.4125035958717733e-126, 32'sd-2.5035330132146845e-120, 32'sd2.06321475770467e-117, 32'sd5.594142120269132e-127, 32'sd-5.40223006376439e-117, 32'sd5.333253362521611e-127, 32'sd-1.319662473165756e-120, 32'sd0.011868580495614742, 32'sd-0.051532880157104985, 32'sd-0.025116209297410166, 32'sd-0.004083135967319939, 32'sd-1.0875440698829344e-121, 32'sd1.676203416222358e-122, 32'sd2.151181492788832e-122, 32'sd-1.2062263392286968e-123, 32'sd2.1253176076790695e-127, 32'sd1.4882680880023455e-125, 32'sd1.7584907529333476e-121, 32'sd1.335270284305947e-122, 32'sd1.7840552411535168e-125, 32'sd1.1394858225723744e-119, 32'sd3.4145556234649e-122, 32'sd-1.7729060688839785e-114, 32'sd-9.065206409431878e-123, 32'sd6.764474566282269e-126, 32'sd-2.2370870837344337e-124, 32'sd-5.742031424175371e-127, 32'sd-0.04292961916689301, 32'sd-0.011537209261404242, 32'sd0.02253566167089762, 32'sd0.000857437074530413, 32'sd0.052859704155336064, 32'sd-0.009497891745915268, 32'sd-0.04179123406626835, 32'sd-0.07275180345636914, 32'sd0.05546069873462204, 32'sd-0.035861270903376805, 32'sd0.026425076992110892, 32'sd-0.030739518920693553, 32'sd0.000947031037214523, 32'sd-0.04351826650145273, 32'sd-0.11711441070325629, 32'sd0.05567368391430973, 32'sd0.009072309860822357, 32'sd0.03223275828097471, 32'sd-0.045720249071418854, 32'sd0.03953516416564915, 32'sd2.5703189177400196e-119, 32'sd1.9663228555754785e-124, 32'sd7.228602434377275e-117, 32'sd6.609908495268483e-124, 32'sd3.924083031722547e-123, 32'sd6.6230578274698355e-115, 32'sd0.010398424765602562, 32'sd0.022445289675554245, 32'sd0.0433184118282286, 32'sd-0.0468411728887635, 32'sd-0.02228649466283892, 32'sd-0.04524496264396183, 32'sd-0.05429345660784408, 32'sd-0.001169971419636944, 32'sd-0.11521881507138557, 32'sd-0.12392781605361372, 32'sd-0.12578605677563073, 32'sd-0.0585752475704778, 32'sd-0.05750339732154134, 32'sd-0.011562451654739228, 32'sd-0.021413993882894392, 32'sd0.004596811631807837, 32'sd0.02637606028568678, 32'sd0.09324303694632811, 32'sd0.05139038148661407, 32'sd-0.07689067562456363, 32'sd-0.10173685974078009, 32'sd-0.06854917235492151, 32'sd0.029011223480278524, 32'sd-0.041400093780910883, 32'sd-1.2704418683780442e-118, 32'sd-3.1465359964799275e-114, 32'sd7.923221431264591e-120, 32'sd2.661799782076842e-116, 32'sd-0.020980143789510457, 32'sd-0.02804094668052451, 32'sd0.08995359029447843, 32'sd0.09992875709249137, 32'sd-0.05186975912167657, 32'sd0.041375356221477456, 32'sd-0.040696848037077356, 32'sd-0.10506232157533356, 32'sd0.008370754202994157, 32'sd0.00627401369772214, 32'sd0.012103602185389334, 32'sd-0.07555927221697134, 32'sd0.09358090019852766, 32'sd-0.039805154032873866, 32'sd0.10428816152842871, 32'sd0.04913861709940545, 32'sd0.03474527546644551, 32'sd0.005069513208025896, 32'sd0.09473089934148504, 32'sd0.002588565351797323, 32'sd0.03656986858994845, 32'sd0.00674251883521629, 32'sd0.0015515189962616682, 32'sd0.0828618282580751, 32'sd-0.003241506958793185, 32'sd-1.3194249276546505e-118, 32'sd1.055328553557875e-125, 32'sd-0.009875333557142537, 32'sd-0.04615640899155771, 32'sd0.0275647855511718, 32'sd0.02953902531528581, 32'sd0.00399041821282042, 32'sd0.01253383960972892, 32'sd-0.021810976362236927, 32'sd-0.026323424672357862, 32'sd-0.07973208595792708, 32'sd-0.101724732564091, 32'sd-0.06422272009962778, 32'sd0.046499660286865904, 32'sd0.08067183427738654, 32'sd0.05926911164992271, 32'sd-0.03869565723487928, 32'sd0.09862671026813333, 32'sd-0.045052940976292116, 32'sd-0.14668219518573883, 32'sd-0.054111620001961125, 32'sd-0.12815931878311745, 32'sd-0.13825791801689266, 32'sd0.002322236511222664, 32'sd0.042308655408831684, 32'sd0.0640366947622385, 32'sd0.07680911923969387, 32'sd0.019520199751194334, 32'sd0.04303831806170518, 32'sd8.046329079245526e-118, 32'sd0.010130026739051256, 32'sd0.1058265319441556, 32'sd0.15204819191843558, 32'sd0.0538145415588525, 32'sd-0.010172208689159532, 32'sd-0.03720140212041494, 32'sd-0.0381792924929454, 32'sd0.024684660647109672, 32'sd0.026589859441109094, 32'sd0.06009231512923731, 32'sd-0.1503387036790139, 32'sd-0.09905093144148647, 32'sd-0.00964945486440608, 32'sd0.026016608151052393, 32'sd0.08691684086643671, 32'sd-0.02514479876287559, 32'sd-0.022155582288801982, 32'sd-0.04910576805973096, 32'sd0.03495823722458818, 32'sd0.0034518223690865255, 32'sd-0.09894230196422113, 32'sd0.018036605591869512, 32'sd-0.04300808784111249, 32'sd-0.016046092990362006, 32'sd-0.020824677811256923, 32'sd0.048645611265611136, 32'sd-0.06003096841085123, 32'sd-1.372818030616228e-123, 32'sd0.019398953286150763, 32'sd0.0061035849250065085, 32'sd0.015952684501935176, 32'sd0.02850849548598751, 32'sd0.0038967042902770615, 32'sd-0.021690582344781124, 32'sd-0.029454662135230306, 32'sd-0.013915718650867418, 32'sd-0.02218002134243212, 32'sd-0.07524770032203747, 32'sd-0.13288393465530368, 32'sd-0.12236971707589349, 32'sd0.08888013235384094, 32'sd0.1320006021435245, 32'sd0.23288232139131274, 32'sd0.17582297223195917, 32'sd0.12855887152345238, 32'sd0.19374669373736905, 32'sd0.07213022494832379, 32'sd-0.027986623859609892, 32'sd0.13526586149648245, 32'sd-0.06526148120913357, 32'sd0.046641667207747185, 32'sd0.014954892314140659, 32'sd0.011585076174699864, 32'sd-0.017633372660292253, 32'sd0.04946080579115575, 32'sd0.01134801625991604, 32'sd-0.04126961217372459, 32'sd-0.022824213047462114, 32'sd-0.10054138422900996, 32'sd-0.05738965524745614, 32'sd-0.07551485818495192, 32'sd-0.004180550814148277, 32'sd0.07380546874832437, 32'sd0.005295141892821611, 32'sd-0.06837303239474465, 32'sd-0.10345557000368535, 32'sd0.020463283128184157, 32'sd0.08743151204701664, 32'sd-0.04670705176986481, 32'sd0.12462811766807834, 32'sd0.24087371244339895, 32'sd0.1385127251635278, 32'sd0.14597946119628996, 32'sd0.25477340735909115, 32'sd0.0714231604184982, 32'sd0.14463326169100454, 32'sd0.12476448133307651, 32'sd0.012166416744940673, 32'sd-0.15838180781041775, 32'sd0.08834272320744314, 32'sd0.1447497392417123, 32'sd0.059114158848429715, 32'sd-0.04809070667331112, 32'sd0.04881911389586497, 32'sd0.021641569832180522, 32'sd-0.024672909169227455, 32'sd-0.048923913435365, 32'sd-0.017822299564903613, 32'sd0.09759490503763496, 32'sd0.056041398261888836, 32'sd-0.05586593050400122, 32'sd-0.13024243207463682, 32'sd-0.005628893133100496, 32'sd0.02147300694809119, 32'sd0.07696846633526634, 32'sd-0.04730846275727071, 32'sd0.08735805496835711, 32'sd0.01841857399858747, 32'sd0.14466499603039565, 32'sd0.26636697149189015, 32'sd0.14097074940524226, 32'sd0.25460473488799784, 32'sd0.05805371420111152, 32'sd0.09096188903106803, 32'sd0.11682873130281542, 32'sd-0.06632430446587445, 32'sd0.030719478908777922, 32'sd0.13416575408238152, 32'sd0.12692439968662994, 32'sd0.0742317618268461, 32'sd0.04574637144714099, 32'sd-0.006823403642936886, 32'sd0.06698965841165086, 32'sd0.06982583724332035, 32'sd-0.007449449350094602, 32'sd0.04649424257683323, 32'sd-0.004217836203519396, 32'sd-0.09304151104411923, 32'sd-0.013857971739316403, 32'sd-0.007504495131371703, 32'sd0.09208295278307423, 32'sd0.043002298444466694, 32'sd0.047911650399267196, 32'sd0.0431285887353387, 32'sd0.0377289240559416, 32'sd0.19029325606589417, 32'sd0.14163586084319452, 32'sd0.028045176371516187, 32'sd0.21199594857765003, 32'sd0.09011879001445366, 32'sd0.13043290218791068, 32'sd0.13347850636460415, 32'sd0.006530335764267591, 32'sd-0.08762453855011708, 32'sd-0.029757582384892876, 32'sd0.10286799161836321, 32'sd0.09239653322209436, 32'sd0.027311874191932865, 32'sd0.07269328355053666, 32'sd-0.020593498623769895, 32'sd-0.005366132467098935, 32'sd0.0639910734053278, 32'sd0.012464549973074076, 32'sd0.04559300057991101, 32'sd-0.021177934303662098, 32'sd0.054599719319465764, 32'sd0.02190028614420389, 32'sd0.030294931220350617, 32'sd-0.05136101870526298, 32'sd-0.021309290395749688, 32'sd0.0017677914602339017, 32'sd-0.08890604133163763, 32'sd0.019252498936599707, 32'sd0.010126533487308248, 32'sd-0.06501221418468973, 32'sd-0.03526284902640986, 32'sd-0.08306864128503423, 32'sd0.008426098980831872, 32'sd0.04964216032427779, 32'sd0.01581979596778613, 32'sd-0.006878729103864508, 32'sd-0.01765406495024884, 32'sd-0.038191208148986265, 32'sd-0.0482377384564768, 32'sd0.049800559236675104, 32'sd0.04779705839078184, 32'sd-0.059470094211492984, 32'sd-0.006197271417858167, 32'sd0.06638237684744597, 32'sd0.09267702632357763, 32'sd0.08374861711021554, 32'sd0.012801510805544347, 32'sd-0.08244479956852957, 32'sd0.03037842505645969, 32'sd0.08420234048185711, 32'sd0.057561272565947876, 32'sd-0.07955643294793867, 32'sd-0.025938101401358975, 32'sd0.11407648112797666, 32'sd-0.16602951230000568, 32'sd0.018896047279638995, 32'sd0.15820010242972665, 32'sd0.011099753044678196, 32'sd-0.13256904848680973, 32'sd-0.02378669562886534, 32'sd-0.05561539009405838, 32'sd-0.08648185550470502, 32'sd0.07378579269466924, 32'sd-0.11418259700110839, 32'sd-0.12371198459432574, 32'sd-0.001962773519655873, 32'sd0.0204494531770925, 32'sd-0.027338846517286075, 32'sd-0.09389800360082629, 32'sd-0.10522019774926042, 32'sd0.018624739786759954, 32'sd0.012333821682870059, 32'sd-0.042609979177625275, 32'sd0.0441367671585647, 32'sd0.008574202624321925, 32'sd-0.09198414615763785, 32'sd-0.169394607588487, 32'sd-0.07311252247273808, 32'sd-0.0872970618574505, 32'sd-0.015849207451997745, 32'sd-0.03914127710991838, 32'sd-0.051285871399141085, 32'sd-0.1585318834679249, 32'sd-0.08316069272378528, 32'sd-0.0614169073891777, 32'sd0.13543434366817642, 32'sd-0.05841357589874848, 32'sd0.059287082972947824, 32'sd0.030251687098617152, 32'sd-0.012708674568069818, 32'sd0.009187182138055468, 32'sd-0.05669401920226947, 32'sd-0.06552738956213856, 32'sd-0.08659625925978423, 32'sd-0.06946093979993499, 32'sd-0.09926974230124723, 32'sd-0.14751971328808297, 32'sd-0.06379068268016774, 32'sd-0.02232453558425031, 32'sd-0.04916875616090373, 32'sd0.005115329533318108, 32'sd-0.07672850478341985, 32'sd0.050287582043473986, 32'sd-0.045530456857343, 32'sd-0.01579471382216711, 32'sd-0.0036277237525455777, 32'sd0.042260000667994804, 32'sd-0.034474437465195795, 32'sd-0.1748356354650822, 32'sd-0.12890524211540696, 32'sd-0.1179002869294005, 32'sd-0.14768391546470275, 32'sd0.04637218811601501, 32'sd-0.027148032542414085, 32'sd-0.10242731506595264, 32'sd-0.05499575746212083, 32'sd0.034676670920240536, 32'sd0.0057334347085503555, 32'sd-0.08726412747631755, 32'sd-0.019796600733067823, 32'sd-0.17531595771486483, 32'sd-0.13226933730664933, 32'sd-0.08291157451626234, 32'sd-0.0056497485283063835, 32'sd-0.002060413716443683, 32'sd-0.061347649670658554, 32'sd0.025029414757769475, 32'sd-0.00422757532849315, 32'sd-0.007440527630580854, 32'sd0.027590894677679514, 32'sd-0.07751828326880647, 32'sd-0.06302468268187682, 32'sd0.05786689967903663, 32'sd0.014587663171344502, 32'sd-0.12206708222921879, 32'sd-0.17120460946659594, 32'sd-0.12704308837165354, 32'sd-0.24493266241216796, 32'sd-0.15542483212665498, 32'sd-0.06952103830576914, 32'sd-0.04571688604143287, 32'sd0.06039519532897388, 32'sd0.012854291242638993, 32'sd-0.050146125150164776, 32'sd0.11666790567937935, 32'sd0.08283441151172109, 32'sd0.02875520724294507, 32'sd-0.1190464772208275, 32'sd-0.0924841146145734, 32'sd-0.23772002115358443, 32'sd-0.08130631594747705, 32'sd0.06267714339627957, 32'sd0.004405341429182203, 32'sd-0.007963405232869366, 32'sd0.052682561699058376, 32'sd0.000681035349879879, 32'sd0.06882956986480683, 32'sd-0.061191850772762686, 32'sd-0.07708700303982721, 32'sd0.06412913886097785, 32'sd-0.07764241287086522, 32'sd0.016250284219621033, 32'sd-0.07573663900153828, 32'sd-0.19850411053355366, 32'sd-0.03772263500652806, 32'sd-0.1651018526201541, 32'sd-0.05766818078017359, 32'sd-0.03660194071564757, 32'sd-0.06072860212685121, 32'sd0.10044874855915836, 32'sd-0.006645917267984223, 32'sd-0.1049937776201248, 32'sd0.0029533455048437987, 32'sd-0.06425540874500996, 32'sd-0.022728454946038392, 32'sd-0.1300445153864846, 32'sd-0.16111337682844862, 32'sd-0.14269401202674614, 32'sd-0.000187569866066305, 32'sd0.0072374512553865285, 32'sd-0.0492357584783765, 32'sd-0.027663387822099567, 32'sd0.0493771761640373, 32'sd-0.02920473488170687, 32'sd0.02115658896444258, 32'sd0.03547852385529565, 32'sd-0.08039554037510209, 32'sd-0.09758773155020391, 32'sd-0.0432530706883318, 32'sd-0.06252724106319366, 32'sd0.070906796984314, 32'sd0.0014478677788908885, 32'sd-0.06068300342462331, 32'sd-0.15188400098511168, 32'sd-0.04422853665204954, 32'sd-0.10929588732138393, 32'sd-0.1325434527360602, 32'sd-0.007752230442964667, 32'sd-0.03467729527875737, 32'sd-0.0347803186207346, 32'sd0.022093969776358562, 32'sd0.0006231059766259719, 32'sd-0.0771743495890399, 32'sd-0.2308847828317594, 32'sd-0.08833444593638316, 32'sd-0.07579813687831459, 32'sd0.10791304741666335, 32'sd0.06580157197430178, 32'sd-0.12601130672270755, 32'sd-0.06707076180989986, 32'sd2.723334027797227e-121, 32'sd0.03148435736428469, 32'sd0.0694413743901089, 32'sd0.057251142719055396, 32'sd-0.0748038985122674, 32'sd-0.12962650000979617, 32'sd-0.10739736840367364, 32'sd0.045516725880024554, 32'sd0.08188801419262375, 32'sd-0.044175661047711236, 32'sd-0.14108036191980536, 32'sd-0.08753170057066183, 32'sd-0.016525523367986655, 32'sd-0.026688870074771553, 32'sd-0.12895436409181082, 32'sd0.01827492696540117, 32'sd-0.05007524842683507, 32'sd0.10576954124814678, 32'sd0.09341720673406144, 32'sd0.03888648987840115, 32'sd-0.1238166298500017, 32'sd-0.2001305194088694, 32'sd-0.13808651596919339, 32'sd-0.13841781353507052, 32'sd0.031796242121428585, 32'sd0.11837990046820665, 32'sd-0.03540062032306978, 32'sd-0.020862062163626516, 32'sd-0.04776815687496392, 32'sd-0.05478229745429585, 32'sd-0.021513022208451166, 32'sd-0.10570095402486111, 32'sd-0.17684019869640977, 32'sd0.011837145715942209, 32'sd0.03541692912938583, 32'sd0.060722247489155445, 32'sd0.07851001409785098, 32'sd-0.00012889501717104396, 32'sd-0.02977039668401324, 32'sd-0.019695637869455877, 32'sd0.10203937857836645, 32'sd0.042087526624208796, 32'sd-0.05851877405395525, 32'sd0.03228469265184196, 32'sd0.11939066523993647, 32'sd0.23487534547432695, 32'sd0.025222008896530125, 32'sd-0.041910312551873, 32'sd-0.18307503889145404, 32'sd-0.06978706743455829, 32'sd-0.045039675582706586, 32'sd-0.039044496196011344, 32'sd0.06700215560034509, 32'sd-0.009504275592780538, 32'sd-0.018363393518100218, 32'sd-0.06096191084193688, 32'sd0.008623348332392585, 32'sd0.05495015591596471, 32'sd0.09946352207309354, 32'sd-0.1289319461920857, 32'sd0.03375071733426136, 32'sd0.08783368072877291, 32'sd0.11500216105745173, 32'sd-0.03246019144226684, 32'sd-0.09436383331936714, 32'sd-0.04958571910270557, 32'sd0.03844550965536875, 32'sd0.032749832293650166, 32'sd0.1574612227805347, 32'sd-0.06659784086870169, 32'sd0.029142455830350605, 32'sd-0.008990536365347801, 32'sd0.02085741352013257, 32'sd0.13388738520936247, 32'sd0.06225903819164632, 32'sd-0.07567837880285634, 32'sd-0.13535430177202767, 32'sd-0.11379189151414246, 32'sd-0.06329537559985521, 32'sd-0.12685216283239323, 32'sd0.10144173222136432, 32'sd0.06576607732405773, 32'sd-0.05271992488819308, 32'sd-0.04024835402614453, 32'sd-3.6326499696217525e-114, 32'sd-0.01883430544921067, 32'sd0.04937514832499897, 32'sd-0.02584081039205956, 32'sd0.022459010838221348, 32'sd0.014474510876589066, 32'sd0.10538005904455344, 32'sd0.062125390877330544, 32'sd-0.014269554232373624, 32'sd-0.12341935700753583, 32'sd0.03686307541736179, 32'sd0.027212023407849912, 32'sd-0.05127481348489925, 32'sd-0.08005140150679259, 32'sd0.027678817618053183, 32'sd-0.006789959290068134, 32'sd0.09464505339786265, 32'sd0.2292237620188292, 32'sd-0.00704795617904195, 32'sd-0.022316158633971708, 32'sd-0.17011547884827766, 32'sd-0.058094028905898216, 32'sd-0.03872815007935019, 32'sd0.01785155705493924, 32'sd0.025377022167637188, 32'sd-0.04405861037351795, 32'sd-0.03235788805102279, 32'sd0.019665433323720692, 32'sd-0.05870843294167215, 32'sd-0.05663632835737232, 32'sd0.007158281662765766, 32'sd-0.05562691928161918, 32'sd-0.06501761446868058, 32'sd-0.024061346369978098, 32'sd0.029932991931394752, 32'sd-0.04615296947053608, 32'sd-0.16002520718825428, 32'sd-0.13342873910515307, 32'sd-0.057962785371947975, 32'sd-0.059447062250898845, 32'sd-0.06561025941349992, 32'sd0.01969813232617128, 32'sd-0.01266835096198655, 32'sd-0.01178184221142428, 32'sd0.08203171033935197, 32'sd0.10348286035095036, 32'sd-0.13825755165156156, 32'sd-0.1242039251421786, 32'sd-0.13708948888783162, 32'sd-0.09955598278480011, 32'sd-0.13708380106245843, 32'sd-0.044306566458869115, 32'sd-0.0015891025288373003, 32'sd0.03894141561134764, 32'sd-0.041899948185044715, 32'sd0.03339281701916493, 32'sd-0.011153769379702382, 32'sd-0.046052636236964324, 32'sd-0.012232697246285118, 32'sd-0.018418373158102658, 32'sd-0.0371065323503395, 32'sd-0.13788159429337835, 32'sd0.09312614754696995, 32'sd-0.054470759301984854, 32'sd-0.09524173576632125, 32'sd-0.1307732207377492, 32'sd0.029654831824595242, 32'sd-0.0053759511693638115, 32'sd0.1600845373591889, 32'sd0.09471055141103307, 32'sd0.13813661606849584, 32'sd0.0237965453166152, 32'sd-0.07595692063990742, 32'sd0.020209972594880176, 32'sd-0.15907508295054884, 32'sd-0.19014397610366218, 32'sd-0.16759438698721074, 32'sd-0.16118300564386445, 32'sd-0.20256501960361656, 32'sd-0.0822710547285152, 32'sd-0.06034261970071009, 32'sd-0.03731701630673132, 32'sd0.001356882142026742, 32'sd0.011904126247257505, 32'sd-7.558541417208581e-121, 32'sd0.030177558442490496, 32'sd0.04079378528341985, 32'sd-0.10081633725813134, 32'sd-0.043150767945084254, 32'sd-0.09989618572333266, 32'sd-0.1453351190239663, 32'sd-0.07415704908766182, 32'sd-0.16723280697846357, 32'sd-0.13781444530631118, 32'sd-0.03871638503155079, 32'sd0.03433822396281524, 32'sd0.003082197040870837, 32'sd0.1374128766412564, 32'sd-0.04893956051648439, 32'sd-0.11450510271183395, 32'sd-0.043855570491681484, 32'sd-0.09023202561268406, 32'sd-0.11516697894687893, 32'sd-0.18581013454280196, 32'sd-0.08237700194772753, 32'sd-0.07864276262093096, 32'sd0.07570775582305682, 32'sd0.04396255086681555, 32'sd-0.03486651133043315, 32'sd0.03378913377448868, 32'sd-0.07762338143273015, 32'sd-3.6297771218438345e-124, 32'sd2.5389273430576484e-124, 32'sd-3.799269149713058e-118, 32'sd0.032023480819881094, 32'sd0.002227474845771968, 32'sd-0.038658516271488315, 32'sd0.1314390892459991, 32'sd0.05150069747776648, 32'sd-0.07256450762885466, 32'sd-0.022623321533374728, 32'sd-0.0594694009216602, 32'sd0.004090069471776259, 32'sd0.10033115377291882, 32'sd0.15529150478149342, 32'sd0.09901538350648935, 32'sd-0.0018981459624095559, 32'sd0.014235240758161027, 32'sd0.03652507706125738, 32'sd0.001720747359919234, 32'sd-0.2136876932559718, 32'sd-0.13216807384971277, 32'sd-0.021110949739433234, 32'sd-0.2654675610566142, 32'sd-0.09544469477937652, 32'sd-0.012141557488114104, 32'sd-0.10212112002480672, 32'sd0.02351739589765432, 32'sd-0.028598021449213983, 32'sd8.955928108086255e-128, 32'sd1.316706551365586e-125, 32'sd-5.012508370063209e-120, 32'sd0.05241679657559297, 32'sd-0.04397519802712273, 32'sd-0.09771304980769442, 32'sd0.04957000946164623, 32'sd-0.01725562742571542, 32'sd0.108884544660588, 32'sd0.10812645325435272, 32'sd-0.08200614022854597, 32'sd0.10671350911565154, 32'sd-0.018896178238371735, 32'sd0.1229315203017379, 32'sd0.04026898035892927, 32'sd0.08353432170507, 32'sd-0.02154504637915952, 32'sd-0.04310923266615223, 32'sd0.07518187392437585, 32'sd-0.08801388061041053, 32'sd-0.04075301575235283, 32'sd-0.1083878049710831, 32'sd-0.03959405260852228, 32'sd0.09611265853714636, 32'sd-0.07143351624648867, 32'sd0.011983642123523703, 32'sd0.04280908629875627, 32'sd0.016084267001992742, 32'sd-8.692138134330791e-130, 32'sd7.51512286094344e-125, 32'sd-3.949291475347575e-124, 32'sd2.079918535223711e-117, 32'sd-0.0047342925553401196, 32'sd-0.06838846715986532, 32'sd0.00617146077655876, 32'sd-0.08780799931155626, 32'sd0.08672382578825916, 32'sd0.06207602887710983, 32'sd0.1909175015281479, 32'sd0.09992786428913374, 32'sd0.025264576658458587, 32'sd0.03363624259448683, 32'sd0.008096619137244522, 32'sd-0.011275270186891758, 32'sd0.08190248644283835, 32'sd-0.023675437573627153, 32'sd0.04709093243754054, 32'sd0.08388758684100395, 32'sd0.03242736422692745, 32'sd-0.04836015707028755, 32'sd-0.05496769525392724, 32'sd0.0752871834198866, 32'sd0.009891743396299267, 32'sd-0.09324159481758947, 32'sd-0.026958197841649857, 32'sd3.47892600780937e-122, 32'sd-4.976547204527782e-124, 32'sd-1.0271767946787477e-120, 32'sd-7.544685003536896e-122, 32'sd2.88541884510506e-120, 32'sd-2.9984981353056717e-120, 32'sd0.0420923115894882, 32'sd0.005163778055370715, 32'sd-0.012219179995046788, 32'sd0.07913554188906213, 32'sd-0.05183374719437695, 32'sd0.06823735558432767, 32'sd0.07401248484453442, 32'sd0.046693369021198916, 32'sd-0.09257737885020137, 32'sd-0.05681167040724563, 32'sd0.035774430886029225, 32'sd0.03568984839325553, 32'sd0.09913525190403742, 32'sd0.12817482340464953, 32'sd0.02891182773588114, 32'sd-0.012509949448525586, 32'sd-0.03382787672564637, 32'sd-0.025378649460650094, 32'sd-0.036443226892338663, 32'sd-0.025971525309694033, 32'sd6.116237649872152e-124, 32'sd7.587422540977916e-127, 32'sd4.6787893695826705e-120, 32'sd-1.8919246978119444e-125},
        '{32'sd9.558672772776355e-117, 32'sd4.2119675076516605e-125, 32'sd-9.71926415461561e-121, 32'sd4.004853328025251e-118, 32'sd-3.2085127020511723e-121, 32'sd7.06578382872149e-121, 32'sd-3.309751353655941e-120, 32'sd8.030393221539229e-127, 32'sd-1.0807685425505812e-120, 32'sd-7.325454046097581e-115, 32'sd-7.302679988266296e-122, 32'sd3.6560277910306204e-116, 32'sd-0.051086611692993576, 32'sd0.04669513204375572, 32'sd-0.034542816853790397, 32'sd-0.08007553926900843, 32'sd2.656374557298732e-122, 32'sd-2.2622382629881715e-124, 32'sd-7.551812958640203e-115, 32'sd7.008969545977551e-127, 32'sd-8.831519210337365e-117, 32'sd-7.365781512638053e-119, 32'sd1.5098985743872943e-115, 32'sd3.1918501847116e-114, 32'sd1.4844772362297267e-125, 32'sd1.5777784152726005e-119, 32'sd1.5778589172916096e-125, 32'sd4.771182469125669e-123, 32'sd6.401021480483625e-126, 32'sd4.2148846400148217e-125, 32'sd2.2816639526385076e-117, 32'sd-2.7523444742030518e-121, 32'sd0.14434321169833805, 32'sd0.006150361156269715, 32'sd0.0754903654896103, 32'sd-0.014163739450512317, 32'sd0.08305801148251507, 32'sd0.004196896009418839, 32'sd0.04200062197562328, 32'sd0.01996855283483159, 32'sd0.0207388780523621, 32'sd0.07478226334832379, 32'sd0.08604357061090957, 32'sd0.049154130269617034, 32'sd0.007118395755198642, 32'sd0.061014085237802676, 32'sd0.02347554555310915, 32'sd-0.015327110914977628, 32'sd0.08182287127924814, 32'sd0.031182984157600267, 32'sd0.04633350035499602, 32'sd0.00543934806711916, 32'sd-1.7211552413520415e-124, 32'sd2.501575524680191e-120, 32'sd7.189568683028159e-125, 32'sd-4.4323792353727306e-120, 32'sd7.379806806918904e-115, 32'sd1.0709019935388055e-121, 32'sd0.06742589308050097, 32'sd0.005000067790087103, 32'sd0.022404777020680538, 32'sd0.06583332080667861, 32'sd-0.050259082707218655, 32'sd-0.027719387110898174, 32'sd-0.035382473471764556, 32'sd0.009367378163441313, 32'sd-0.11766115713840726, 32'sd-0.04549842854085068, 32'sd-0.025810827579208204, 32'sd0.10061661063857147, 32'sd0.09786651774711856, 32'sd0.022445291739241403, 32'sd-0.036288578503074403, 32'sd-0.11315269288710637, 32'sd0.11214980775583902, 32'sd0.01885734288824763, 32'sd0.11234198480350693, 32'sd0.09372468959375922, 32'sd0.1157446005613782, 32'sd-0.0054605841284138465, 32'sd-0.018213770018828252, 32'sd0.06561513794037181, 32'sd-5.583814025002054e-115, 32'sd-3.9645800113448326e-119, 32'sd6.984072664849211e-122, 32'sd-3.2927352533350317e-118, 32'sd0.07658615355929002, 32'sd0.07726227259681023, 32'sd0.0273155765515413, 32'sd-0.06435442540600785, 32'sd0.013832119996848115, 32'sd-0.08688583958163099, 32'sd0.18075738135790467, 32'sd0.08693109319428609, 32'sd0.09393088342384781, 32'sd-0.047917226707037575, 32'sd-0.027958580878668864, 32'sd-0.017863268477733507, 32'sd0.012028593596904096, 32'sd0.07666230181686476, 32'sd-0.003910601292713713, 32'sd-0.05822285985433677, 32'sd0.11700984831381131, 32'sd0.1391610789722428, 32'sd0.12324496791169706, 32'sd0.0014684294569009826, 32'sd-0.045601445921950014, 32'sd-0.10382406744155868, 32'sd-0.10466643609345277, 32'sd0.00048823296971262786, 32'sd0.07546027821591604, 32'sd1.76964152918953e-121, 32'sd-4.305817366475402e-118, 32'sd0.06239028770030627, 32'sd0.010213530061080575, 32'sd0.03660537583536563, 32'sd-0.07142883475338933, 32'sd0.034205267600241875, 32'sd-0.008128871157001744, 32'sd-0.07897637814374092, 32'sd0.06336133925906369, 32'sd0.0797403931812206, 32'sd0.055346248672649694, 32'sd0.10715593294653256, 32'sd0.0032987621819555346, 32'sd0.06365519088779018, 32'sd0.11668402779232305, 32'sd0.16045083174662852, 32'sd0.07945550622559674, 32'sd-0.05802456291395906, 32'sd0.08363367721889356, 32'sd-0.014146096665469246, 32'sd0.07835996384972617, 32'sd0.012734998100890975, 32'sd-0.1060938425015448, 32'sd0.026711217174313275, 32'sd-0.03703864957141828, 32'sd0.02747224307441656, 32'sd0.07765788468302338, 32'sd0.014583034863307722, 32'sd-5.888096672262801e-127, 32'sd0.00927738209228446, 32'sd0.034724863909101775, 32'sd0.009787899647185945, 32'sd0.0003300939769747547, 32'sd-0.04187062866100907, 32'sd-0.10617086527653695, 32'sd-0.02343823369235136, 32'sd-0.004622621436276187, 32'sd0.015473038661661295, 32'sd-0.0018547349467963065, 32'sd-0.012077163643155685, 32'sd-0.14987596117037735, 32'sd-0.11296796864751696, 32'sd-0.07468942871896128, 32'sd0.06613124072334801, 32'sd-0.0037064028716554593, 32'sd-0.0060014300691669294, 32'sd-0.01686496895515055, 32'sd0.048101010418967284, 32'sd0.0614013875272558, 32'sd-0.05605960500478164, 32'sd-0.09530292068723169, 32'sd-0.012902094629292126, 32'sd0.04984599346378947, 32'sd0.013753575840115882, 32'sd0.0632537080863697, 32'sd-0.05555137692511371, 32'sd-1.1278829237649843e-115, 32'sd0.0038174618544677304, 32'sd-0.02493715237984526, 32'sd0.09111374915122121, 32'sd0.05214857872175648, 32'sd0.08366932001451696, 32'sd0.11344217916415719, 32'sd-0.045508782470461334, 32'sd0.023279508608029482, 32'sd-0.12077341944533217, 32'sd-0.06682994688677361, 32'sd-0.05617136828392686, 32'sd-0.025501296125377895, 32'sd-0.061658252337655525, 32'sd0.0014694941274214245, 32'sd0.038410281733793614, 32'sd0.038629799945976324, 32'sd-0.09768625204494188, 32'sd-0.06322933132237263, 32'sd-0.02810764718138009, 32'sd-0.0058229891441821235, 32'sd-0.02566704453117332, 32'sd-0.10616224848667591, 32'sd0.02017232439040817, 32'sd0.0684157319524187, 32'sd0.017625933612200224, 32'sd0.04822031288919782, 32'sd0.052575389183411, 32'sd0.010579853382167692, 32'sd0.06279188764330867, 32'sd0.06707533994528715, 32'sd0.01114378362835391, 32'sd-0.07805464164041663, 32'sd-0.10363658137705975, 32'sd-0.07499503290179096, 32'sd-0.03838735780876338, 32'sd0.044191266448764505, 32'sd-0.10893163518939737, 32'sd-0.04985947759615256, 32'sd0.007705672225979916, 32'sd0.08526510413484216, 32'sd0.03799819375469084, 32'sd0.15851946227599942, 32'sd0.0462276892347814, 32'sd-0.0628485188398001, 32'sd0.013740372540427115, 32'sd-0.18000439724794712, 32'sd-0.21104971118850915, 32'sd-0.11465695647636238, 32'sd-0.0968638565180314, 32'sd-0.06437073126723564, 32'sd-0.16694779335361576, 32'sd-0.11882982058621103, 32'sd0.013438490527812147, 32'sd0.004628317654385156, 32'sd-0.078012711658724, 32'sd0.025735159315281073, 32'sd-0.04162592917331029, 32'sd0.05633845292892525, 32'sd0.08380265944992851, 32'sd-0.06966974158324217, 32'sd-0.09259162874314421, 32'sd-0.14431987912686367, 32'sd-0.10853060607973387, 32'sd-0.01352542121724644, 32'sd-0.04290567419136433, 32'sd-0.1316496956711237, 32'sd-0.014391683838695017, 32'sd0.021481530593405285, 32'sd-0.029868901735270768, 32'sd-0.028904501966554138, 32'sd-0.09388860234991765, 32'sd-0.1425518471256315, 32'sd-0.0761272451643661, 32'sd-0.17440813255601992, 32'sd-0.14159367069947307, 32'sd-0.12696037129069856, 32'sd0.014701146992662248, 32'sd-0.029612730545863962, 32'sd-0.02025953124710335, 32'sd-0.02172785376636223, 32'sd0.03994280358114079, 32'sd0.08767634554214601, 32'sd0.05590355908081327, 32'sd0.038596779077179115, 32'sd-0.12653093804640642, 32'sd-0.032133133384083856, 32'sd0.08667228853668066, 32'sd-0.01837590058972763, 32'sd-0.1708882159483519, 32'sd-0.014714571311249702, 32'sd-0.05024748263855859, 32'sd-0.0760878351230132, 32'sd-0.07259158916500741, 32'sd-0.050484938390091154, 32'sd-0.07078059814756203, 32'sd0.016485705395754002, 32'sd0.055787738240994825, 32'sd0.009574069345416332, 32'sd-0.04813902239170025, 32'sd0.07788165491604, 32'sd0.12225070209723411, 32'sd-0.0021833090203150045, 32'sd-0.01567067936077877, 32'sd-0.024671386500822116, 32'sd0.07117121758123504, 32'sd0.11985822536741808, 32'sd0.002885832571881038, 32'sd0.11973989846429757, 32'sd0.0895471893600362, 32'sd-0.02704044797516763, 32'sd-0.010878115386348523, 32'sd0.0118619371832423, 32'sd-0.09970589252129074, 32'sd-0.04712560618111317, 32'sd0.019838965387856712, 32'sd0.04881767267162739, 32'sd-0.02868416927907738, 32'sd-0.11423877809801591, 32'sd-0.05222263636023362, 32'sd-0.0682122747057423, 32'sd-0.11202043394636477, 32'sd-0.10870690943427234, 32'sd-0.06055558598929931, 32'sd0.09348488061604786, 32'sd0.1365615863422597, 32'sd0.13528465105840315, 32'sd0.06966916421640615, 32'sd0.06654259186511381, 32'sd0.15743998024256023, 32'sd0.09535754128181795, 32'sd0.0567451420314411, 32'sd0.020442506771480847, 32'sd-0.02216322441750088, 32'sd-0.05330072712676248, 32'sd0.14757067462638748, 32'sd0.12795046623019682, 32'sd-0.0467729534670277, 32'sd0.06957777797292776, 32'sd0.08374468593485701, 32'sd-0.05024404051158402, 32'sd0.03419174134406594, 32'sd0.06505498303613252, 32'sd0.019465286417419687, 32'sd0.02865629980329647, 32'sd-0.1193799425844099, 32'sd-0.08109068192132243, 32'sd-0.11822457004810738, 32'sd-0.053369721944917396, 32'sd0.005248694712894997, 32'sd0.0915164689595134, 32'sd-0.07028703015696122, 32'sd0.014444902421114916, 32'sd0.037642388137496485, 32'sd0.040813775859236935, 32'sd-0.05581647090034689, 32'sd0.0717386137164078, 32'sd0.26548631666107464, 32'sd0.05102715844639135, 32'sd0.08464249280404809, 32'sd0.0010848505267639513, 32'sd-0.022451055314984848, 32'sd-0.0374785680587207, 32'sd0.043562053308353256, 32'sd-0.05808420057386352, 32'sd-0.010715012893350842, 32'sd0.008656247343262546, 32'sd0.07012795327715719, 32'sd0.034735136605987704, 32'sd0.06094234241514732, 32'sd-0.0222388202038228, 32'sd0.10529563362959492, 32'sd0.002482217102288443, 32'sd-0.017581209613464526, 32'sd0.016081052850548637, 32'sd-0.020472304930073376, 32'sd-0.05315933011607109, 32'sd0.0035498428252715535, 32'sd-0.0692303111213446, 32'sd-0.11492981236102619, 32'sd-0.038682288976412106, 32'sd-0.021346472516683358, 32'sd0.05541847921740989, 32'sd-0.0774405023215935, 32'sd0.029312118893457993, 32'sd-0.0061946012281169655, 32'sd-0.09225518621999476, 32'sd-0.0010658442267060502, 32'sd-0.072427191040129, 32'sd-0.1003696118311261, 32'sd0.05970256973277916, 32'sd0.01887664634702625, 32'sd-0.1015082586295125, 32'sd-0.14031171292784395, 32'sd-0.04319144202299457, 32'sd0.002312896885959533, 32'sd0.08132816865096545, 32'sd0.020645852185474198, 32'sd-0.018322267470667754, 32'sd0.06807511372578816, 32'sd-0.00968492910534406, 32'sd-0.11641172355186856, 32'sd-0.06714739277390151, 32'sd0.013299902767048316, 32'sd-0.044761076459508685, 32'sd0.04165907637209252, 32'sd-0.012399375431463, 32'sd-0.037230430476010344, 32'sd-0.12280639417082338, 32'sd-0.06469286852824596, 32'sd0.011478218634014341, 32'sd0.04295127688951262, 32'sd0.026227302961287557, 32'sd-0.19401930962831995, 32'sd-0.14074347127690556, 32'sd-0.002911744892134576, 32'sd0.02323170107589225, 32'sd-0.04261746800149874, 32'sd0.028602734633800753, 32'sd0.12644959290907476, 32'sd-0.19326608811752288, 32'sd-0.07248732786836337, 32'sd-0.009647757438122713, 32'sd0.02384394698006913, 32'sd0.11396471110344973, 32'sd0.029094606246955843, 32'sd-0.058092271645968835, 32'sd0.08215732936605735, 32'sd0.08277244480792878, 32'sd-0.15474304789353127, 32'sd-0.1502847834801427, 32'sd-0.028059060549496227, 32'sd-0.06128862305346775, 32'sd0.13035415104506237, 32'sd-0.046244944954659604, 32'sd-0.16308094914750895, 32'sd-0.09619833240341012, 32'sd-0.05738384880505495, 32'sd-0.03583675284588794, 32'sd-0.04402023981755075, 32'sd-0.05585813712743697, 32'sd-0.24089727692735935, 32'sd-0.22940524400693807, 32'sd-0.07364711466973126, 32'sd-0.01122489770129102, 32'sd0.06154674453692797, 32'sd0.07436091677794301, 32'sd-0.0016870390941145252, 32'sd-0.03687340062506696, 32'sd-0.05802827152043819, 32'sd0.01739307841827637, 32'sd-0.041067097340635864, 32'sd0.04800842974972081, 32'sd0.053240416061167486, 32'sd0.09041566228992429, 32'sd0.04505808553588255, 32'sd0.09937831742827037, 32'sd-0.012512134066592228, 32'sd-0.030382348091569932, 32'sd-0.09140241904664945, 32'sd0.021958970898569026, 32'sd0.051730764881579926, 32'sd-0.07449105430480726, 32'sd0.03792985058880282, 32'sd-0.0375113161522097, 32'sd0.019720052583677383, 32'sd0.018329470599856283, 32'sd-0.16685158306414066, 32'sd-0.0824380227529182, 32'sd-0.1701890734338042, 32'sd-0.0824897615428886, 32'sd-0.05812714761625267, 32'sd0.03296121135405976, 32'sd0.040780840905307425, 32'sd-0.025399844581923896, 32'sd-0.008805468159772123, 32'sd-0.10902339231172246, 32'sd0.021487502172013204, 32'sd0.07719562479828412, 32'sd-0.016629859092208484, 32'sd0.005083820136808546, 32'sd0.06643810607435639, 32'sd0.06948678436909111, 32'sd-0.0044026371054715135, 32'sd-0.001099028006583659, 32'sd0.022202557258164397, 32'sd0.06095382836736007, 32'sd-0.09630109822652862, 32'sd-0.051089205610396884, 32'sd-0.053222671118038245, 32'sd0.004123332445425031, 32'sd-0.011855057779310259, 32'sd-0.03542093450576683, 32'sd-0.04382568870614102, 32'sd0.012293133192745253, 32'sd-0.1723260363046996, 32'sd-0.011374128256691943, 32'sd-0.2183066343963611, 32'sd-0.02732939087942501, 32'sd-0.1220471878070431, 32'sd-0.027101661473397327, 32'sd-0.024344894209288055, 32'sd0.0326519679821356, 32'sd0.010479741244775749, 32'sd-0.006899970213378301, 32'sd-0.010043434350553106, 32'sd0.06803922959326089, 32'sd0.05981667936840876, 32'sd-7.227466358737192e-120, 32'sd0.01803352762184248, 32'sd0.08429692928627879, 32'sd-0.003125556187134273, 32'sd-0.03444186915991601, 32'sd0.11472365288279865, 32'sd0.11182248382813716, 32'sd0.07601367486204273, 32'sd0.09026630811241888, 32'sd-0.06303638553415532, 32'sd0.038172901454903284, 32'sd-0.06467143546306568, 32'sd-0.12770252275893038, 32'sd-0.0013866331286278592, 32'sd-0.07382014448243536, 32'sd-0.04863118559243094, 32'sd-0.09814428675859195, 32'sd-0.13328095342432517, 32'sd-0.0683205789746912, 32'sd-0.13010327016531584, 32'sd-0.06623997799072616, 32'sd-0.02641448544842744, 32'sd0.003196889522560313, 32'sd0.08972448752451291, 32'sd-0.08063739305915205, 32'sd-0.13069413235577096, 32'sd-0.04669182656041754, 32'sd-0.0939966548699484, 32'sd-0.008529954978452848, 32'sd0.01870475396479924, 32'sd0.07577037747301986, 32'sd0.005787349645043531, 32'sd-0.008180872207861175, 32'sd0.04346928959404261, 32'sd0.1255402633973114, 32'sd0.04617079068369583, 32'sd0.09913334980545209, 32'sd-0.009953897822894948, 32'sd0.062086760405617385, 32'sd-0.07527145441133762, 32'sd-0.009191138725579485, 32'sd0.007542372174691181, 32'sd0.015467216680778795, 32'sd-0.04648042137557327, 32'sd-0.01965781865671683, 32'sd-0.10350960998301971, 32'sd-0.0948875674366665, 32'sd-0.15469682322358233, 32'sd-0.12961420484457783, 32'sd-0.042227435230693985, 32'sd-0.011814232369050465, 32'sd-0.03821662508591346, 32'sd0.0555348359744386, 32'sd0.027464638095622763, 32'sd-0.0482465255448549, 32'sd-0.03675169846575938, 32'sd0.01756548594324168, 32'sd-0.08073389019837313, 32'sd0.010627922095526897, 32'sd-0.029685934163600488, 32'sd-0.0010889681452216794, 32'sd-0.022829976760344428, 32'sd0.1380087792000484, 32'sd0.12816358676176778, 32'sd0.10541973397745572, 32'sd-0.032677276650477184, 32'sd-0.03387292062170881, 32'sd0.041647040742312354, 32'sd0.08230697936660256, 32'sd-0.021930117136554933, 32'sd0.07388879474479969, 32'sd0.07659546756464021, 32'sd-0.032046383304777507, 32'sd-0.08278300802371831, 32'sd-0.04112967438591653, 32'sd-0.0843274867604739, 32'sd0.011397855296500954, 32'sd-0.06596657477609219, 32'sd-0.15663719960070183, 32'sd0.015836521963737374, 32'sd-0.0235543966503851, 32'sd0.0643422718656114, 32'sd-0.05203343316299288, 32'sd-0.047051738431701094, 32'sd-1.9948513265547252e-126, 32'sd0.03850418235695336, 32'sd-0.004165434192623016, 32'sd-0.03701055951257604, 32'sd-0.03247176531076588, 32'sd0.12112187161180611, 32'sd0.15682698018732996, 32'sd0.009032701746938371, 32'sd0.044579565332915634, 32'sd0.16817208079092472, 32'sd0.04559838786110509, 32'sd-0.028215127106000985, 32'sd0.11520093793913515, 32'sd0.08405349116860059, 32'sd0.17159721139386983, 32'sd0.14148364375168704, 32'sd0.09937867779715052, 32'sd-0.051619408236686225, 32'sd-0.015511120791228489, 32'sd-0.08538639232351357, 32'sd0.0009651586321380834, 32'sd-0.021452457687517516, 32'sd0.02403358052527947, 32'sd-0.029907882839812924, 32'sd0.005624460318720995, 32'sd0.041140630442192315, 32'sd-0.0961027398263958, 32'sd0.11528681792326843, 32'sd-0.01689168119791558, 32'sd-0.043544557986586685, 32'sd-0.08189553273026134, 32'sd-0.12792573347489308, 32'sd-0.18201335135278804, 32'sd-0.0312761526659638, 32'sd0.0844181723513797, 32'sd-0.010963622280750259, 32'sd0.04410609131518577, 32'sd0.052332234135480576, 32'sd0.11643499069576027, 32'sd0.10854376572229806, 32'sd0.1548198450308135, 32'sd-0.006094275365005761, 32'sd0.17780465923750907, 32'sd0.039137255681738065, 32'sd0.0201278628261384, 32'sd0.09044886758858825, 32'sd0.08320176582565038, 32'sd-0.07661663211640583, 32'sd0.006992373337207877, 32'sd0.005782539476296487, 32'sd0.029419414055523736, 32'sd0.018909196089281675, 32'sd0.013464578357780806, 32'sd-0.04058970414048684, 32'sd-0.043474251324150726, 32'sd-0.007236602816592021, 32'sd0.11800840252129462, 32'sd0.11705889701610685, 32'sd0.08375384016712652, 32'sd0.08868788317305175, 32'sd-0.14530463936806362, 32'sd-0.11783522309543526, 32'sd-0.0713781422068463, 32'sd-0.1287228165484295, 32'sd-0.011401457562203135, 32'sd-0.046528115916117586, 32'sd0.15042561333765733, 32'sd0.08671575870368137, 32'sd-0.007738495987717448, 32'sd0.09294056270619815, 32'sd0.05145215602848736, 32'sd-0.014549206905128594, 32'sd-0.014551061500451311, 32'sd0.05129980565615578, 32'sd-0.0031994949407599897, 32'sd0.03968374733587042, 32'sd-0.009458782767248566, 32'sd0.1080734713065208, 32'sd-0.16536954072779697, 32'sd0.05327025944172166, 32'sd-0.03411659336218291, 32'sd0.012084561374326248, 32'sd-0.012709562756548998, 32'sd0.026256510860002684, 32'sd-9.300909585398142e-116, 32'sd0.011612556949408782, 32'sd-0.039730465979150364, 32'sd-0.043589740715529214, 32'sd-0.06133934664716307, 32'sd-0.023130993352844596, 32'sd-0.068658302478436, 32'sd-0.14235403370527638, 32'sd-0.03289693834661632, 32'sd0.013101473809937947, 32'sd0.009365928330602229, 32'sd-0.026696002295003667, 32'sd0.10467295454881569, 32'sd-0.019058256956012338, 32'sd-0.0593316084844476, 32'sd0.01521345072168765, 32'sd0.05660833034813502, 32'sd-0.01771441370017723, 32'sd-0.08753670197602535, 32'sd-0.004966312926643367, 32'sd0.02434110734145159, 32'sd-0.10217307131892128, 32'sd-0.07956660067744833, 32'sd0.054621042786598746, 32'sd0.009315803560525136, 32'sd-0.007738402152221587, 32'sd0.10802377968656289, 32'sd3.653428879626543e-126, 32'sd2.5568300123850668e-126, 32'sd-1.1283807090602498e-125, 32'sd0.0850233833150347, 32'sd0.006321664934759958, 32'sd-0.04043587802815659, 32'sd-0.03710548907276809, 32'sd0.012119451550684657, 32'sd0.028242792588838685, 32'sd-0.0678923570363721, 32'sd0.0538843988670526, 32'sd0.039964049817516265, 32'sd-0.1074258125815992, 32'sd0.024999531488476025, 32'sd-0.11467831317405182, 32'sd-0.07406011436034454, 32'sd-0.08269679723558825, 32'sd0.06735613099752058, 32'sd-0.07525294356466654, 32'sd-0.048970508840326735, 32'sd-0.043145974301788965, 32'sd-0.019197595701595734, 32'sd0.1832285458746144, 32'sd-0.05990310764493334, 32'sd-0.11072466593338064, 32'sd-0.0016995062478771322, 32'sd0.034910251314564246, 32'sd-0.035764602621444944, 32'sd-1.1767715342055358e-115, 32'sd-2.0986783814823955e-123, 32'sd-3.5760079511392323e-128, 32'sd0.04010808854156194, 32'sd-0.06292436065500491, 32'sd0.00494938079611182, 32'sd-0.06469454748197569, 32'sd-0.05423175914715899, 32'sd-0.029407629074560192, 32'sd-0.033959706260022274, 32'sd-0.03215462130803323, 32'sd-0.01302487041349211, 32'sd-0.05738915021164989, 32'sd-0.015470715667172794, 32'sd-0.04780793123483717, 32'sd0.0890002279654293, 32'sd-0.03777878259467905, 32'sd-0.009980708424705925, 32'sd-0.0819575746189231, 32'sd0.16950696184726827, 32'sd0.07291737205549696, 32'sd0.013060295014016439, 32'sd0.045896149870576566, 32'sd-0.016563882834671185, 32'sd-0.04183316048289884, 32'sd-0.03489429408135521, 32'sd0.02700564837015332, 32'sd0.016852039344603328, 32'sd1.3416205422984664e-122, 32'sd-2.4025296100162127e-120, 32'sd-3.994855883818666e-118, 32'sd1.1959931590679924e-125, 32'sd0.07216998653470669, 32'sd0.023550275187920654, 32'sd-0.03462179190314629, 32'sd-0.04467214975272887, 32'sd0.0013486598376399248, 32'sd-0.0919001346058581, 32'sd-0.05297553352245607, 32'sd-0.18464108738141827, 32'sd-0.06465424394347108, 32'sd-0.05813506504514257, 32'sd-0.03962167042903566, 32'sd-0.11314240690449792, 32'sd0.11713083861050545, 32'sd0.06772546499261886, 32'sd-0.13334165566152822, 32'sd-0.007085282740734696, 32'sd-0.0414072810716626, 32'sd0.058285873533463754, 32'sd0.06634378018112193, 32'sd0.024912684833844165, 32'sd-0.04300010061884341, 32'sd0.008179225553758827, 32'sd0.039676534342215596, 32'sd1.1194099396120874e-115, 32'sd-3.4021207462105826e-129, 32'sd7.490348492101574e-117, 32'sd-8.129732387224284e-123, 32'sd2.4415002259750088e-126, 32'sd-2.5962557732485944e-121, 32'sd0.06350587782052984, 32'sd0.04972450731263939, 32'sd0.01604499286763144, 32'sd-0.0178703147709238, 32'sd0.08464208693454128, 32'sd0.06862942308272839, 32'sd0.05171216387781084, 32'sd0.07844542722098018, 32'sd0.05763550504802586, 32'sd-0.08149821349322096, 32'sd-0.01755676817300803, 32'sd0.10608179504127815, 32'sd0.08946624573956205, 32'sd0.006676737074815416, 32'sd0.009977464210521479, 32'sd0.024213340326063263, 32'sd0.029298824299038632, 32'sd0.08831304979462366, 32'sd-0.04608115328979656, 32'sd0.050874349447479754, 32'sd1.663004954124585e-120, 32'sd-7.580791668168467e-123, 32'sd6.7738428260410796e-124, 32'sd-8.820260763147281e-127},
        '{32'sd6.946567124720819e-124, 32'sd2.1686735714672864e-127, 32'sd-4.615170805231431e-128, 32'sd7.345494507657487e-120, 32'sd-1.2687460213829739e-121, 32'sd1.827481557843685e-126, 32'sd3.0026000965198144e-126, 32'sd-5.3945401301739565e-118, 32'sd-9.34227479741028e-122, 32'sd9.668870543985718e-120, 32'sd2.4781198234164126e-116, 32'sd-9.532434087407331e-120, 32'sd-0.04461636245464157, 32'sd-0.024080605641253184, 32'sd-0.01651202998698632, 32'sd0.010217974842910815, 32'sd2.5614154634012917e-126, 32'sd-1.3246729702209987e-122, 32'sd3.3807142488071185e-115, 32'sd4.135169880651024e-118, 32'sd1.058728236440256e-124, 32'sd-8.60870897682777e-117, 32'sd-1.9794703354260873e-121, 32'sd8.286470043948026e-121, 32'sd9.028371446627426e-125, 32'sd-2.126128372212687e-115, 32'sd-2.6516240614475074e-122, 32'sd7.001232478163766e-122, 32'sd-3.3512978479840994e-120, 32'sd-2.1422751309005214e-124, 32'sd6.805980381280123e-126, 32'sd-1.5414236928932272e-114, 32'sd-0.043364480556262686, 32'sd0.006321761282893071, 32'sd-0.059168072200023736, 32'sd0.012432117402100241, 32'sd0.030912482437425556, 32'sd-0.07031672188351269, 32'sd0.0006100160003146056, 32'sd-0.08512431281158842, 32'sd-0.06370471704947303, 32'sd-0.021867735052903976, 32'sd-0.04249740622153214, 32'sd-0.01849179166763139, 32'sd-0.08729234885020555, 32'sd0.004597985552285383, 32'sd0.05443106791863175, 32'sd-0.12460323601999314, 32'sd-0.05592665259123753, 32'sd-0.08499170056688243, 32'sd-0.07140849120338208, 32'sd-0.0288412242582171, 32'sd2.4418817791883587e-125, 32'sd-1.5277835174192367e-117, 32'sd-8.30990299040733e-120, 32'sd-1.7713601423330976e-117, 32'sd7.107310727283588e-127, 32'sd-1.8586785205550877e-125, 32'sd-0.03615765464202755, 32'sd-0.0104197850627202, 32'sd0.00508437642818423, 32'sd0.011865665814372971, 32'sd-0.05845905510744624, 32'sd-0.09721427177556193, 32'sd-0.10382951616389621, 32'sd0.045082500098354426, 32'sd-0.06971428211216213, 32'sd-0.15118884581463424, 32'sd-0.04937644767795131, 32'sd-0.16701891871499536, 32'sd-0.14444776205138224, 32'sd-0.035819505429713454, 32'sd-0.15105503666878348, 32'sd0.03700379127320304, 32'sd0.16461555032630953, 32'sd-0.11843979079190768, 32'sd0.03494155845494544, 32'sd-0.014883673341189589, 32'sd0.11348044342385241, 32'sd-0.10677497941899622, 32'sd-0.049749616376089385, 32'sd-0.06790274892118167, 32'sd-1.964976722144205e-120, 32'sd-2.248688300743602e-124, 32'sd-7.532313287628582e-124, 32'sd1.3359192603598962e-117, 32'sd-0.06245174897722155, 32'sd-0.07766619056066217, 32'sd0.025385183181672183, 32'sd-3.660465273200678e-05, 32'sd-0.09113987592904114, 32'sd-0.10181714741293907, 32'sd-0.1011307911062076, 32'sd-0.027231922161546202, 32'sd-0.07740307163071969, 32'sd0.055788560632776645, 32'sd-0.12994639868041072, 32'sd-0.17456600969794211, 32'sd-0.07768045317523879, 32'sd-0.06930533998820655, 32'sd-0.14542777917325259, 32'sd0.00791426215907686, 32'sd0.09421922295567707, 32'sd-0.06253584655568341, 32'sd0.06061088707653933, 32'sd0.10065758383979977, 32'sd0.10209617800835387, 32'sd0.016000930447497775, 32'sd0.09475452138931013, 32'sd-0.10676672244919637, 32'sd-0.00020304382236981154, 32'sd-1.8843754946986617e-128, 32'sd-7.567285125044111e-115, 32'sd0.014677669682177027, 32'sd0.03928758873799227, 32'sd-0.06879626522285241, 32'sd-0.04982288425204711, 32'sd-0.012404655307134431, 32'sd0.0017748736864310621, 32'sd0.02813817037318708, 32'sd-0.023950713089717704, 32'sd-0.2605233917103129, 32'sd-0.19695719539073958, 32'sd-0.13758028875261255, 32'sd-0.0887574402892088, 32'sd-0.10380750309585299, 32'sd-0.14149013157585077, 32'sd0.01703247197802347, 32'sd0.022728161799001646, 32'sd0.0906630931128707, 32'sd0.0284928497126434, 32'sd-0.15055478461886046, 32'sd-0.09475368228610538, 32'sd-0.0015548529870656734, 32'sd0.0354557862424563, 32'sd0.08109292713153601, 32'sd0.003820712947075929, 32'sd-0.07278379222140577, 32'sd-0.07630491916707376, 32'sd-0.011590625762073153, 32'sd-2.221942304794302e-125, 32'sd-0.019177278016013006, 32'sd-0.04204154060931324, 32'sd-0.05873969396739706, 32'sd0.04697329440708517, 32'sd-0.033972752740442015, 32'sd-0.04991267507576271, 32'sd-0.06064391414401437, 32'sd-0.045148165632519645, 32'sd-0.0945065895713455, 32'sd-0.10467829882434841, 32'sd-0.001637010254625639, 32'sd0.07220327600541845, 32'sd0.05243315096910804, 32'sd0.026987494254730515, 32'sd-0.026457360560969367, 32'sd-0.03028955072293315, 32'sd-0.011732802900370574, 32'sd-0.014531526971762862, 32'sd0.07064645321514368, 32'sd0.057116952763299624, 32'sd-0.1156896640577484, 32'sd-0.11005224281049451, 32'sd-0.08807981218160545, 32'sd-0.061645221105055416, 32'sd0.02214337979182342, 32'sd0.054301319541630345, 32'sd-0.03489014047757432, 32'sd-2.0596798855179655e-124, 32'sd0.04937139746826472, 32'sd0.040921951964611215, 32'sd-0.0393114561814086, 32'sd-0.10627257991573337, 32'sd-0.16160622978428404, 32'sd0.016704501746448403, 32'sd-0.08231727629608532, 32'sd-0.031805067482341604, 32'sd0.038892442130753165, 32'sd0.0704602421047044, 32'sd0.028175968734403208, 32'sd0.07111283147692288, 32'sd0.00725709759845994, 32'sd0.09003921728824679, 32'sd0.02868519311660359, 32'sd0.030372392823163792, 32'sd0.0470044639195892, 32'sd-0.024250216130314323, 32'sd0.10111880639041688, 32'sd0.21353403809972427, 32'sd0.07210440346140064, 32'sd0.023707754133058152, 32'sd-0.07477631565061742, 32'sd-0.009894489869696349, 32'sd0.03244473983593865, 32'sd0.06983794471061112, 32'sd-0.06566536592381692, 32'sd-0.007447142053519033, 32'sd-0.08661472822173333, 32'sd0.019816552874179272, 32'sd0.009518862313538863, 32'sd-0.06260885028605293, 32'sd0.007304486482135066, 32'sd0.01621863809970439, 32'sd-0.07500944381953724, 32'sd-0.001484911723889564, 32'sd-0.06307072724901237, 32'sd0.028246995994248843, 32'sd0.004746844185659794, 32'sd0.06639689672501736, 32'sd0.044423807875485985, 32'sd-0.02055152960842869, 32'sd0.007215439712537639, 32'sd-0.006482042326581394, 32'sd0.10654252363843807, 32'sd0.15909518512240214, 32'sd0.13394777036107858, 32'sd0.150793422618828, 32'sd0.11488382530480441, 32'sd0.1159040194638522, 32'sd0.021960982095084017, 32'sd0.04566298295831001, 32'sd0.057247131499502425, 32'sd0.022181086472497096, 32'sd0.026939191530697456, 32'sd-0.023082989571903013, 32'sd0.005671577415623574, 32'sd-0.08979182152051171, 32'sd-0.05488744497846585, 32'sd-0.011969017629351712, 32'sd0.003242897728808683, 32'sd0.02222957225128934, 32'sd-0.03339459625033199, 32'sd-0.09191267272838796, 32'sd-0.09520907290097232, 32'sd-0.1357207108599254, 32'sd-0.15145626760344694, 32'sd-0.12775814920178355, 32'sd-0.06735826154797632, 32'sd-0.039370721209966146, 32'sd0.0068633553869991235, 32'sd0.050592003782426356, 32'sd0.16870518432015527, 32'sd0.21132791290280778, 32'sd0.03217437085277986, 32'sd0.10242291554111117, 32'sd0.07997824724107414, 32'sd0.04987651751227321, 32'sd0.07308376487548057, 32'sd0.15033935119620334, 32'sd0.08605638432434375, 32'sd-0.031175740775230488, 32'sd-0.013791268513953195, 32'sd-0.05199172344184532, 32'sd0.012650335677224102, 32'sd0.08297594027764892, 32'sd-0.06886567085506037, 32'sd-0.14241271170810946, 32'sd-0.002826416172917166, 32'sd-0.04645048429275967, 32'sd-0.07106386598095038, 32'sd0.02070287593099996, 32'sd-0.03366483835026861, 32'sd0.007043902483225036, 32'sd0.03867601649193185, 32'sd-0.02890246046774527, 32'sd0.00029122903386267156, 32'sd-0.041808417914913625, 32'sd0.05271109676350128, 32'sd0.12642563317706912, 32'sd0.07449424266405191, 32'sd0.10627730528882984, 32'sd0.08350530766111768, 32'sd0.09892686975172728, 32'sd0.08824931720147208, 32'sd0.03175509662185918, 32'sd0.05381006643338352, 32'sd-0.008603962775759533, 32'sd0.05591516464695092, 32'sd-0.0005809237500445972, 32'sd0.022270888649365085, 32'sd-0.00976762489834927, 32'sd0.010745768405711377, 32'sd-0.06198120839245458, 32'sd0.006564253582944349, 32'sd0.03220872938259746, 32'sd0.10005765422159243, 32'sd0.009029508431569891, 32'sd0.09945386054615839, 32'sd-0.10903265296021333, 32'sd0.06239338638091145, 32'sd0.0646698341658556, 32'sd-0.019443214727565588, 32'sd-0.052385200300027954, 32'sd-0.09819898921550463, 32'sd-0.05557356867216908, 32'sd-0.0006937865573399473, 32'sd-0.09044619998865563, 32'sd-0.21400270918810352, 32'sd-0.10069555102271406, 32'sd-0.018113369941910148, 32'sd-0.03895386534852695, 32'sd0.028035369569030806, 32'sd0.01433249857440125, 32'sd0.060019215181146876, 32'sd0.07019284244489428, 32'sd0.0860416186715569, 32'sd-0.033110150612522905, 32'sd-0.06013476942336891, 32'sd0.038223727280359505, 32'sd-0.004255523491212799, 32'sd-0.11577945188975021, 32'sd0.0032505688828564, 32'sd0.11470640529402522, 32'sd0.1155902570024286, 32'sd0.009084055815955974, 32'sd-0.029174432424605313, 32'sd0.050417535164033335, 32'sd0.15341426216408194, 32'sd-0.035784855140386915, 32'sd-0.1397247233422195, 32'sd-0.13607489349544336, 32'sd-0.14632433800540653, 32'sd-0.17097972692931246, 32'sd-0.028470617536956233, 32'sd-0.2466636933015504, 32'sd-0.23605005456790684, 32'sd-0.14898296325615246, 32'sd-0.08799325942391943, 32'sd-0.057241119576125286, 32'sd0.010445034890243184, 32'sd0.11634264249415167, 32'sd0.02703172625541313, 32'sd-0.1425636720154884, 32'sd0.06283158699457371, 32'sd0.0318687329425015, 32'sd-0.06585987533596648, 32'sd-0.04742278708003106, 32'sd-0.028699560086636437, 32'sd0.04440007964143649, 32'sd0.08841437125260083, 32'sd0.11372300177632802, 32'sd0.005847474074232393, 32'sd0.15537079592823455, 32'sd0.14684836446928837, 32'sd0.15724543724798468, 32'sd0.046755764249231724, 32'sd-0.07072557294178528, 32'sd-0.20201698008333385, 32'sd-0.028338574385140244, 32'sd-0.12299495092290116, 32'sd-0.23944771399781098, 32'sd-0.028441112165666887, 32'sd-0.15283974713728582, 32'sd-0.21784498759070048, 32'sd-0.06673863626304842, 32'sd-0.0431161232705106, 32'sd0.04937297830194493, 32'sd0.08021699237722403, 32'sd0.11035946381373325, 32'sd0.008216745840127335, 32'sd-0.09529629631187182, 32'sd0.006521577481565521, 32'sd-0.17896677028107255, 32'sd0.019473386096532465, 32'sd0.032379064954862195, 32'sd-0.013540257472009128, 32'sd0.023519162283573612, 32'sd0.06788612764446421, 32'sd0.08689285665095801, 32'sd0.04171102006742166, 32'sd0.018090483499577804, 32'sd0.18716864726116644, 32'sd0.1909124339921926, 32'sd0.08583956902443128, 32'sd0.08436725351375933, 32'sd-0.07060903075930183, 32'sd-0.062129005392268566, 32'sd-0.0037943739922359073, 32'sd-0.008690845651571164, 32'sd-0.11121800862176624, 32'sd-0.16080161015364847, 32'sd-0.15511118950173364, 32'sd-0.1602817691734508, 32'sd-0.035358070431111645, 32'sd0.08190497321327908, 32'sd0.0828977405792325, 32'sd-0.04984593188027101, 32'sd-0.082906173922147, 32'sd0.026333685991693858, 32'sd0.07545873782378995, 32'sd0.026990958594358464, 32'sd-0.014448238111094002, 32'sd-0.028344392643371377, 32'sd-0.014802273733223693, 32'sd-0.037852862974827775, 32'sd0.08675626340876684, 32'sd-0.0034942273619582797, 32'sd0.07386594140170431, 32'sd0.06815896008425869, 32'sd0.10167530168988281, 32'sd0.03199365395080853, 32'sd0.06087690812766535, 32'sd0.22478724167615083, 32'sd0.07662629128929074, 32'sd-0.09388785088570345, 32'sd0.0979300873317606, 32'sd0.12546641550373916, 32'sd0.10072697188110066, 32'sd-0.027392666716091488, 32'sd-0.016828992566550936, 32'sd-0.10969682473903937, 32'sd0.002487790065084975, 32'sd0.05148043779056561, 32'sd0.007303791865204632, 32'sd-0.018654545367514205, 32'sd-0.14565978109753447, 32'sd0.03564078837413121, 32'sd0.030667199663904497, 32'sd-0.06949727784488038, 32'sd-0.03042277591353132, 32'sd0.056904806159293976, 32'sd-0.07978454094921753, 32'sd0.0028347214893524736, 32'sd0.10817710482772788, 32'sd0.082512470228675, 32'sd0.039869724434087234, 32'sd0.1409947462649449, 32'sd-0.04655977990734266, 32'sd0.06462615497985308, 32'sd0.08182225689014057, 32'sd0.14203342679792758, 32'sd-0.009138083741135554, 32'sd0.10928609904206672, 32'sd0.0539695248052628, 32'sd0.01945993430185656, 32'sd0.06794338760354506, 32'sd0.01672656854699701, 32'sd-0.02637045122178566, 32'sd0.06287365904963539, 32'sd-0.07698031075349382, 32'sd0.022544926552577536, 32'sd-0.09572250240473529, 32'sd-0.06072643866512035, 32'sd0.0018645735027065262, 32'sd-0.06348504052455653, 32'sd-0.09944696386601107, 32'sd-0.012294223278694158, 32'sd-0.021164959295361423, 32'sd0.007244462891515441, 32'sd-0.11441256445062298, 32'sd0.008269369425527612, 32'sd-0.03055734628012569, 32'sd-0.05167438540952029, 32'sd0.08192708033225617, 32'sd-0.055569676689842556, 32'sd-0.028341996518954048, 32'sd-0.05647838315193418, 32'sd0.15107007716630544, 32'sd0.13418468873338635, 32'sd0.1356496214240457, 32'sd0.11581871400785768, 32'sd0.1370888517590685, 32'sd0.04250093519764369, 32'sd0.08274462202683862, 32'sd0.11192295075746325, 32'sd0.034745802239882585, 32'sd-0.02065936739330355, 32'sd0.006915552083634039, 32'sd0.02779988978676979, 32'sd-0.1292689752707482, 32'sd-0.10183578220891068, 32'sd-0.0571579356932593, 32'sd-0.17042704616514603, 32'sd-0.11639354206447618, 32'sd0.09601499567799328, 32'sd-0.0323363154394674, 32'sd1.1195583385756793e-116, 32'sd0.03139805742030711, 32'sd0.004518699574588471, 32'sd0.09254395056257309, 32'sd-0.07783146869303097, 32'sd-0.04919994983616087, 32'sd-0.0045636957586667175, 32'sd-0.10047861569593532, 32'sd0.0006588980016891877, 32'sd0.04284408607188038, 32'sd0.17276099489486998, 32'sd0.23136221488433983, 32'sd0.27491748064319566, 32'sd0.20173785240101322, 32'sd0.1448914192211653, 32'sd0.18769165283223332, 32'sd0.08446251573899469, 32'sd0.14354510837156953, 32'sd0.11120201745568879, 32'sd0.025256773657676028, 32'sd-0.03501783634118136, 32'sd0.006335984910344864, 32'sd-0.06110005325013922, 32'sd-0.1935295419228761, 32'sd-0.183255147412026, 32'sd-0.024754861447263295, 32'sd-0.009600685905486378, 32'sd-0.11963403591782841, 32'sd-0.017184898420637206, 32'sd0.024839676045549933, 32'sd0.08441117914438105, 32'sd0.08353643615858894, 32'sd-0.05698762090003181, 32'sd-0.08329915594908205, 32'sd-0.07473043608320055, 32'sd-0.04276930933805677, 32'sd-0.1641314898703954, 32'sd-0.12842613745801562, 32'sd0.05408028668746902, 32'sd0.18103186600166057, 32'sd0.0689784454604211, 32'sd0.11878496769617787, 32'sd0.07494330219445983, 32'sd0.07588947229795974, 32'sd0.18302860121470094, 32'sd0.11772843041110181, 32'sd0.015600250196050137, 32'sd0.11903909439618245, 32'sd0.013412329600578771, 32'sd-0.024615517240514483, 32'sd-0.04738834396723883, 32'sd-0.17597923083687378, 32'sd-0.07516931298981314, 32'sd0.1049897253406998, 32'sd0.03608068066409898, 32'sd-0.01843601153778632, 32'sd-0.045317358792140945, 32'sd-0.013925022648400317, 32'sd0.048954654576370826, 32'sd0.04939420183172777, 32'sd0.04735698784587637, 32'sd-0.14070146562662053, 32'sd-0.17347309233231212, 32'sd-0.18537603089935029, 32'sd-0.18436677493062173, 32'sd-0.26438738503328874, 32'sd-0.030336788699520775, 32'sd-0.03581440683856542, 32'sd-0.0825022705128301, 32'sd0.017738275954630078, 32'sd0.021294816077845228, 32'sd0.012569798604338033, 32'sd0.18172964566009045, 32'sd0.09978309111214911, 32'sd0.1347000134658197, 32'sd0.021003305461618445, 32'sd-0.0017904192598436725, 32'sd-0.039319115427272955, 32'sd-0.06742330224617568, 32'sd0.005327259301951846, 32'sd-0.025477290997901737, 32'sd-0.03661428633857157, 32'sd0.0265564696597531, 32'sd-0.06459258146321475, 32'sd-2.1976640660341743e-124, 32'sd-0.023087585156437943, 32'sd-0.024319126705259642, 32'sd-0.06782436896216373, 32'sd0.04815898034181692, 32'sd0.05951835928866408, 32'sd0.011427459457225723, 32'sd-0.1777837003647451, 32'sd-0.17992934813720696, 32'sd-0.19445466431578318, 32'sd-0.18403397667206478, 32'sd-0.12364596956271214, 32'sd-0.18124108442103037, 32'sd-0.081844240029478, 32'sd-0.04976138397304028, 32'sd0.09130867177716553, 32'sd0.16913705483009947, 32'sd0.16860539457774723, 32'sd0.1155133455088235, 32'sd-0.01524486743707255, 32'sd0.010271296740170332, 32'sd0.04476593311168523, 32'sd0.09240409229566698, 32'sd0.05309028577109105, 32'sd0.042813947103573266, 32'sd0.09497361435357868, 32'sd-0.061217991621214864, 32'sd0.05346614768431782, 32'sd0.020897934004125766, 32'sd-0.013104208372705482, 32'sd0.0778152525261799, 32'sd-0.015285686064784192, 32'sd0.024137070347489464, 32'sd0.0543923906698971, 32'sd-0.03354440827722641, 32'sd-0.013482465608282203, 32'sd-0.004131069223463483, 32'sd-0.11604373059358666, 32'sd-0.15291441325788996, 32'sd-0.1422748664930449, 32'sd-0.23606031471823272, 32'sd-0.15612157238854227, 32'sd0.038898244584600374, 32'sd0.09629604564949254, 32'sd0.2332494227314501, 32'sd0.11814858681467105, 32'sd0.07735133548647505, 32'sd-0.04282853810002378, 32'sd0.010198760600801045, 32'sd0.06746177163471478, 32'sd0.010281650801636403, 32'sd0.04815776302856582, 32'sd0.11236417962101061, 32'sd0.02746425686339745, 32'sd-0.05856716163800686, 32'sd-0.02506538982736801, 32'sd-0.03900901521574276, 32'sd0.04367808283159781, 32'sd0.05295735188671014, 32'sd-0.07501459373150919, 32'sd0.020033674025559195, 32'sd0.00824006076618907, 32'sd-0.02329845079541469, 32'sd-0.0649863437295937, 32'sd-0.05792820435842302, 32'sd0.10552396650138635, 32'sd0.04565062548473417, 32'sd-0.04678117863759595, 32'sd-0.035577537167860704, 32'sd-0.006929602058679873, 32'sd0.08923264259505921, 32'sd0.13885572267207183, 32'sd0.017322196207796597, 32'sd0.009358359464541827, 32'sd-0.04118360452629021, 32'sd-0.10946938541582137, 32'sd0.1017126260010908, 32'sd0.09228310022078705, 32'sd0.03751157906863437, 32'sd0.02765844573844632, 32'sd0.06656732256747437, 32'sd-0.19026333186787045, 32'sd-0.03834752036743753, 32'sd-0.016080020277783286, 32'sd-2.0118357772083207e-127, 32'sd-0.03395876029155809, 32'sd-0.054036174332437334, 32'sd0.04739892067676201, 32'sd0.07083911379049139, 32'sd0.06439188402728757, 32'sd-0.05015095216753151, 32'sd0.030783507919592088, 32'sd0.07880414795418034, 32'sd-0.027591154299406593, 32'sd0.07305074239743667, 32'sd0.037381265411358035, 32'sd0.0587509504726183, 32'sd0.17898876104637115, 32'sd-0.02060863488468673, 32'sd0.035638351018079495, 32'sd0.020211843251531508, 32'sd-0.16437197086959637, 32'sd-0.11837100885535838, 32'sd-0.03017168733600346, 32'sd-0.020091141676481527, 32'sd0.1587984489709837, 32'sd0.10855752186463648, 32'sd0.06996788888451835, 32'sd-0.07330323927409829, 32'sd-0.10027056727626898, 32'sd-0.035440025857281614, 32'sd-6.731508998485278e-123, 32'sd-1.43940138405255e-123, 32'sd-3.1966666369311884e-122, 32'sd-0.03644999187704794, 32'sd-0.0011171689276698404, 32'sd0.08642263110269893, 32'sd0.016675830589979585, 32'sd-0.008171045112625378, 32'sd0.071729576322301, 32'sd0.03921841679244224, 32'sd0.01340219310248119, 32'sd0.09441511107211725, 32'sd0.08348299900568974, 32'sd0.09343618433093961, 32'sd0.14091268753046793, 32'sd0.14443826702312373, 32'sd0.15325439333885507, 32'sd-0.047411131592366644, 32'sd-0.022779282724788533, 32'sd0.008260519591745095, 32'sd0.020362153156178127, 32'sd0.11311084055754024, 32'sd0.11878228017100252, 32'sd0.11092110127401371, 32'sd-0.03127566249299428, 32'sd-0.06542834305720896, 32'sd-0.09736740314418307, 32'sd-0.03293393160530294, 32'sd3.6251197336117786e-114, 32'sd8.311715665714732e-124, 32'sd-7.931894817839643e-120, 32'sd-0.07286954193138032, 32'sd-0.08685092896469768, 32'sd0.0632130242048025, 32'sd-0.0248270084801238, 32'sd0.09461016758503356, 32'sd-0.028008351038303136, 32'sd0.045554036309509126, 32'sd-0.004386404109515112, 32'sd0.06474274979134345, 32'sd0.13795611974245847, 32'sd0.0173506500430142, 32'sd0.05579158625135247, 32'sd-0.12018209044191817, 32'sd0.05253798748109174, 32'sd0.00859218474781092, 32'sd0.03015499163129666, 32'sd-0.02769876510093127, 32'sd0.03813463439441363, 32'sd0.04684026654469411, 32'sd-0.03151091012411145, 32'sd0.00896727549615583, 32'sd-0.011923413325235147, 32'sd-0.004341018554746139, 32'sd0.03671556497194084, 32'sd0.039725700871413513, 32'sd8.696309016717881e-127, 32'sd-4.516854353236148e-124, 32'sd-1.1119176866944013e-121, 32'sd7.093061709109423e-126, 32'sd-0.0411416572691332, 32'sd-0.027981329063751757, 32'sd-0.03306762678096514, 32'sd0.028728546598081023, 32'sd0.11672838365102789, 32'sd0.006714959706677693, 32'sd0.03290168886650027, 32'sd0.07894763393431754, 32'sd0.11077966578337312, 32'sd0.10372484739039513, 32'sd0.1799339704936705, 32'sd-0.016488238565342456, 32'sd0.001220718707291276, 32'sd0.012489253476062086, 32'sd-0.043434333285603255, 32'sd-0.09863402745006139, 32'sd-0.1603094472290477, 32'sd-0.021888297854228887, 32'sd0.09067856320040975, 32'sd-0.06068963523390316, 32'sd0.07435168624087851, 32'sd0.08421568672486734, 32'sd0.04332484021534311, 32'sd1.5614124239730235e-127, 32'sd4.68174356840144e-123, 32'sd1.109367921489778e-121, 32'sd2.6313001490532777e-122, 32'sd-1.501852382554876e-115, 32'sd-4.3270716499102425e-125, 32'sd0.017578180678492473, 32'sd0.05190993990782498, 32'sd-0.023845056684681128, 32'sd-0.046526634921447, 32'sd0.011381823864776241, 32'sd0.02120452185511458, 32'sd0.02857462260041057, 32'sd0.05499803118621645, 32'sd0.07316792448950928, 32'sd0.06803647213545438, 32'sd0.06777437404508428, 32'sd-0.021793787830797048, 32'sd-0.12300486487100859, 32'sd-0.10144685506272696, 32'sd0.0036346576964635035, 32'sd-0.10790033915911025, 32'sd-0.04341898443331713, 32'sd-0.08479404125658355, 32'sd0.02232166957435712, 32'sd-0.04647724437658561, 32'sd-5.490674276520945e-128, 32'sd5.922027682760834e-126, 32'sd9.006553913564673e-127, 32'sd-2.032598994168495e-119},
        '{32'sd-1.7842817477916678e-122, 32'sd2.4705881297309804e-125, 32'sd5.497431571555262e-121, 32'sd-1.1880274171727806e-118, 32'sd4.049170736759205e-123, 32'sd-5.152125139383337e-124, 32'sd-2.7693967638770906e-126, 32'sd-8.762853111424339e-122, 32'sd1.7059289551806698e-114, 32'sd-6.017882164189954e-120, 32'sd-2.507749244151397e-126, 32'sd2.9369470054901967e-116, 32'sd0.0466388938275438, 32'sd0.06570703090263211, 32'sd0.04257289551839914, 32'sd-0.07633210798713325, 32'sd1.5960782230517252e-117, 32'sd1.1553817170406894e-125, 32'sd-6.362446843247952e-125, 32'sd-2.486463680768974e-124, 32'sd-5.395480963808592e-120, 32'sd-2.81794671038896e-121, 32'sd3.342508494057024e-122, 32'sd1.052766324521804e-127, 32'sd5.3699615126289635e-118, 32'sd1.190947258642295e-127, 32'sd9.025269742463695e-121, 32'sd-1.2023194085045288e-122, 32'sd3.3875789802076214e-120, 32'sd2.651202427611083e-127, 32'sd1.0038613109301586e-124, 32'sd-5.148277019196826e-121, 32'sd0.05610907761282534, 32'sd0.0385990295109895, 32'sd-0.10791673413123085, 32'sd-0.02328443616111855, 32'sd-0.017556754733401257, 32'sd0.01317765456480483, 32'sd-0.03701531473747482, 32'sd0.08262418440310816, 32'sd-0.008690646198192991, 32'sd0.1202796930953503, 32'sd-0.05006714851793982, 32'sd0.04370478273875376, 32'sd-0.0700673704395723, 32'sd0.022546966231447287, 32'sd0.09742782722490637, 32'sd0.12083276080705596, 32'sd0.04736325588950462, 32'sd0.017988537058612773, 32'sd0.08625062223876626, 32'sd0.09890986184548232, 32'sd-6.53062750202622e-117, 32'sd4.356187597694829e-127, 32'sd2.207661240688798e-118, 32'sd-2.0923933486011577e-117, 32'sd-4.7441964343868206e-126, 32'sd-4.1337387390484286e-117, 32'sd0.10042422494329555, 32'sd0.03593613558628036, 32'sd0.08497734867681363, 32'sd0.02321232760888579, 32'sd-0.01980364298344, 32'sd-0.07796002377253751, 32'sd-0.0023854247031526725, 32'sd-0.09439544830667645, 32'sd-0.041144824351258, 32'sd-0.061493786713596475, 32'sd-0.05575385705783512, 32'sd-0.04039374132423464, 32'sd-0.1062971896045176, 32'sd-0.013034753763742971, 32'sd-0.015797466541515464, 32'sd-0.007610650270227092, 32'sd-0.00800198179865429, 32'sd-0.04562365909355941, 32'sd-0.02753570600131975, 32'sd0.09867198778934995, 32'sd0.12834996767184378, 32'sd-0.03129620812026182, 32'sd0.040713553674719814, 32'sd0.15219661649828123, 32'sd-2.023637689878248e-126, 32'sd-1.6637571331310385e-124, 32'sd3.949711270272022e-123, 32'sd3.2390741713771167e-121, 32'sd0.07103270559569849, 32'sd0.12763199751196846, 32'sd0.059582883920574765, 32'sd-0.046879118541544494, 32'sd-0.13099367495092085, 32'sd0.011001583913188966, 32'sd-0.02159932642904028, 32'sd-0.0585331965581916, 32'sd0.06761963132898127, 32'sd-0.08289841309677973, 32'sd-0.0067555922088895215, 32'sd0.024707987136521784, 32'sd-0.06992915305170834, 32'sd-0.04576576593826897, 32'sd-0.021965304477471564, 32'sd0.16010974608002973, 32'sd0.0680624958130162, 32'sd0.07895045974766349, 32'sd0.014262531870674212, 32'sd0.09580200245818996, 32'sd0.05693493423997983, 32'sd0.014992666885372683, 32'sd0.03637580621102713, 32'sd0.03934812041620693, 32'sd0.09618953173298143, 32'sd-6.572539791740419e-125, 32'sd-3.7956657155594696e-122, 32'sd0.06011924439010198, 32'sd-0.0021328980671612967, 32'sd0.07293857884454659, 32'sd0.03429689961203949, 32'sd0.015117596938087813, 32'sd-0.12390774698906738, 32'sd-0.05837643797016793, 32'sd0.02280972214926435, 32'sd-0.03531897761416512, 32'sd-0.1605906706042969, 32'sd-0.08191009185450941, 32'sd-0.07525649509759108, 32'sd-0.04456416319928774, 32'sd-0.05662957381060999, 32'sd-0.00988988812232282, 32'sd-0.03781363609593768, 32'sd0.026132014647765354, 32'sd-0.015741744181133163, 32'sd0.02273419633365358, 32'sd-0.07126829160229103, 32'sd0.007278394600311645, 32'sd0.027890906069664833, 32'sd0.08304447884157037, 32'sd-0.08369672853434504, 32'sd0.05027700395682606, 32'sd0.023812474558914724, 32'sd-0.025193042394091644, 32'sd2.7371732235942947e-122, 32'sd0.03892676865661495, 32'sd0.0014405138947760398, 32'sd-0.06508766946806874, 32'sd0.10143339125516036, 32'sd0.12476555923289752, 32'sd0.10023766667983337, 32'sd0.04124200431054713, 32'sd-0.024925143493796324, 32'sd-0.12855676413771083, 32'sd-0.15701502749777035, 32'sd-0.12474850116905756, 32'sd-0.02298469335130084, 32'sd-0.0808885982325963, 32'sd-0.02609520693839602, 32'sd-0.029248518016325355, 32'sd-0.0737070317045044, 32'sd-0.03722624994108601, 32'sd-0.034195716047941735, 32'sd-0.09813983463557585, 32'sd-0.006994374627891435, 32'sd-0.015005936001813647, 32'sd0.03815087167517828, 32'sd0.013214614669799863, 32'sd0.026362864962813343, 32'sd0.06752618052919239, 32'sd-0.003757996223147011, 32'sd0.06992528304020572, 32'sd-3.1020948965792e-127, 32'sd-0.01150296049850917, 32'sd0.026017460413347022, 32'sd-0.0874909726783835, 32'sd0.08152389756321869, 32'sd0.016034299978518737, 32'sd0.049315011501895406, 32'sd0.0953427990566306, 32'sd-0.019057567732006984, 32'sd-0.08154730162711668, 32'sd-0.19244907598803027, 32'sd-0.11745574222237501, 32'sd-0.015819018703087127, 32'sd0.0887085715995367, 32'sd0.028819981732023135, 32'sd-0.00851460198527334, 32'sd0.02683694908273525, 32'sd0.12441823955149853, 32'sd0.023516567365927037, 32'sd0.062377886076898884, 32'sd0.10454666697721929, 32'sd0.010885692617679755, 32'sd0.002131719228803041, 32'sd0.006744750837669101, 32'sd0.08678155078412338, 32'sd0.021243376318882137, 32'sd-0.0066594524013792065, 32'sd0.0026721252885390685, 32'sd0.11808964067518182, 32'sd0.07221740457588394, 32'sd-0.020874445661114873, 32'sd0.03347208288452899, 32'sd0.07869138741598142, 32'sd0.006008550732660854, 32'sd-0.05642999944636083, 32'sd-0.03025433520651679, 32'sd-0.1201225787971821, 32'sd-0.023834052618913273, 32'sd0.01899218293239158, 32'sd-0.0981959710065768, 32'sd0.019117762663752008, 32'sd-0.01915118836758181, 32'sd0.15176587828406707, 32'sd0.14929865758659677, 32'sd0.12444345696878938, 32'sd0.12265743462026972, 32'sd-0.06749558445912608, 32'sd-0.10459299812814565, 32'sd-0.013648101263413794, 32'sd0.0059337653816310685, 32'sd-0.005206330085417133, 32'sd0.10832407584236972, 32'sd0.012664670001055691, 32'sd0.07035385738596997, 32'sd0.06222843322087622, 32'sd-0.01630010992488663, 32'sd0.019876677802949688, 32'sd0.0017460648449875314, 32'sd-0.0076517038649831825, 32'sd0.07891310078587047, 32'sd0.06164180956944871, 32'sd-0.008205841561863247, 32'sd0.07663332402243113, 32'sd0.068822741388731, 32'sd0.08984540073709027, 32'sd-0.03699041057144288, 32'sd-0.05168920981174934, 32'sd-0.07843072062330435, 32'sd-0.05957969489727651, 32'sd0.09749440152108892, 32'sd0.21332798135996714, 32'sd0.14323499761716355, 32'sd-0.014689129479180035, 32'sd0.04223216990621659, 32'sd0.043252643770508234, 32'sd0.002274169883603689, 32'sd-0.04765138602369383, 32'sd-0.016625011305930158, 32'sd0.023096081389840473, 32'sd-0.03537094024142625, 32'sd0.09441110102450993, 32'sd0.03229131041557304, 32'sd-0.02817826282041193, 32'sd0.030449265118701496, 32'sd0.11632469207406779, 32'sd0.09019285052091881, 32'sd0.05683180212713877, 32'sd-0.028825824799696555, 32'sd-0.004536125690655779, 32'sd-0.002103308617551334, 32'sd0.03016042669965531, 32'sd0.08225733467745636, 32'sd0.08895949877444179, 32'sd0.005929837743241409, 32'sd-0.18569749317138298, 32'sd-0.2420419890061914, 32'sd-0.21734586355181795, 32'sd0.037001697991876144, 32'sd0.21651869681543365, 32'sd0.06282409172696708, 32'sd-0.08494593307778409, 32'sd-0.06160671289136609, 32'sd0.05265749794391703, 32'sd-0.031588657422376674, 32'sd-0.09489289284364776, 32'sd-0.02513951221762557, 32'sd-0.09733117434964957, 32'sd0.000495138488614205, 32'sd0.08956535029483358, 32'sd0.1005889670389981, 32'sd-0.06031683659327581, 32'sd0.06705982135455828, 32'sd0.08346378063676929, 32'sd-0.02949181481554578, 32'sd0.05403266025311451, 32'sd0.0069325276781674865, 32'sd-0.07585325128072246, 32'sd-0.15997764203843237, 32'sd-0.08685663653760162, 32'sd0.003496503405543912, 32'sd0.09133403559504566, 32'sd0.0034775878985163523, 32'sd-0.1763827847879272, 32'sd-0.23830887273491874, 32'sd-0.10550659451596442, 32'sd0.15051395436168327, 32'sd0.09194943453939115, 32'sd0.09115906907759376, 32'sd-0.027468858194439224, 32'sd-0.06996088052666355, 32'sd0.127017988572465, 32'sd0.08000223856595563, 32'sd-0.04062077455099156, 32'sd0.03064224714585001, 32'sd0.12212024203448107, 32'sd0.00472646140564764, 32'sd0.05544363452848155, 32'sd0.06790749316709518, 32'sd-0.008345882089232506, 32'sd0.027118655931414604, 32'sd0.07061637008523546, 32'sd-0.004511386665361094, 32'sd0.08379137692068903, 32'sd0.023301062092469463, 32'sd0.06881656944929365, 32'sd-0.16149986677590408, 32'sd-0.0018139325072597386, 32'sd0.04345191468199221, 32'sd0.03767233115411971, 32'sd-0.055969662193037194, 32'sd-0.039393265299112405, 32'sd-0.16070185155436487, 32'sd-0.11022759187435519, 32'sd0.21792624874493016, 32'sd0.16554040287848898, 32'sd-0.005761750957473103, 32'sd-0.013860215372070314, 32'sd0.07575899597194324, 32'sd0.017869901371334946, 32'sd0.009303793602890383, 32'sd-0.07709686714909057, 32'sd0.005741364033482211, 32'sd0.00965702807953598, 32'sd0.07671922793246483, 32'sd0.09138525573258702, 32'sd-0.0018896629203353091, 32'sd0.04664146899855572, 32'sd0.004439856771646484, 32'sd0.12573732562984372, 32'sd-0.04886005220788287, 32'sd-0.05003723480497717, 32'sd0.000438669812483034, 32'sd-0.06759519721782667, 32'sd-0.06489101478434559, 32'sd-0.0006952731456715639, 32'sd-0.012379071490404524, 32'sd0.07527635074625934, 32'sd0.03143794980816249, 32'sd-0.08481029422085315, 32'sd-0.09485826383099201, 32'sd-0.07445211319209981, 32'sd0.18667183268206636, 32'sd0.1304380590671983, 32'sd0.00762998085423692, 32'sd-0.022953768892623475, 32'sd-0.03913573685921842, 32'sd0.043222311775386386, 32'sd-0.02078263465137062, 32'sd0.0025467931821635406, 32'sd-0.10516032161290302, 32'sd0.016286591009469283, 32'sd-0.07791959850534262, 32'sd-0.12312051501094545, 32'sd0.027085601937182985, 32'sd0.02702487872014295, 32'sd0.09536587374480424, 32'sd0.07464735345509486, 32'sd-0.09036037814987309, 32'sd-0.003747483706382925, 32'sd-0.08186663200546994, 32'sd0.05774860011147564, 32'sd0.01436485377046545, 32'sd0.07204789554786202, 32'sd0.011578362175609237, 32'sd-0.08827406448434227, 32'sd0.08506198074914124, 32'sd0.07387668184303103, 32'sd-0.044184101918266876, 32'sd0.019870916461529484, 32'sd-0.027563392535150295, 32'sd0.14303591155971776, 32'sd0.08942860443319317, 32'sd-0.017797839461558534, 32'sd-0.04292430948411831, 32'sd-0.15691288894554872, 32'sd-0.034504892958242404, 32'sd-0.02111074884491246, 32'sd-0.038504833564742914, 32'sd-0.08277842435824055, 32'sd-0.12953671438910092, 32'sd-0.1269044610488151, 32'sd0.029391440570655823, 32'sd-0.01973139228136042, 32'sd-0.03693378469086917, 32'sd0.166201347585974, 32'sd0.020859997771879243, 32'sd0.06665396341661814, 32'sd0.06612776518280401, 32'sd0.007559155756871879, 32'sd-0.04571130809172724, 32'sd0.022649807815174422, 32'sd0.027274385560230437, 32'sd0.08687170687858455, 32'sd0.03260095360027299, 32'sd0.01906465478761654, 32'sd0.04659930267757227, 32'sd0.0033432084512992704, 32'sd0.01813696489802542, 32'sd0.09029163084240789, 32'sd0.05891879308055368, 32'sd-0.07684335563208569, 32'sd-0.04023150675101335, 32'sd-0.056478151255633956, 32'sd-0.04146856792448489, 32'sd0.08649495088090242, 32'sd0.08560578243821078, 32'sd-0.08160470437965534, 32'sd-0.2453820783866411, 32'sd-0.21925288791362263, 32'sd0.0035458697178337114, 32'sd0.01326243101818322, 32'sd0.007610646606567859, 32'sd0.07805535889969259, 32'sd0.024829380609429484, 32'sd0.08466945603647871, 32'sd-0.004803075780736839, 32'sd-0.06124205394720274, 32'sd0.053376148133437704, 32'sd0.06572201820764091, 32'sd0.15621668056559765, 32'sd0.10632246097291945, 32'sd0.0994176374051374, 32'sd-0.007735861521103687, 32'sd0.003701545736098013, 32'sd-0.06521597185591117, 32'sd-0.026818537122978704, 32'sd0.13821720283872305, 32'sd0.13385282748635066, 32'sd-0.07187609078845561, 32'sd0.0235513453329911, 32'sd-0.022489510063383813, 32'sd0.03146908263419671, 32'sd0.15901435243679318, 32'sd0.034766591296082276, 32'sd-0.09037170471358474, 32'sd-0.09540071774695902, 32'sd-0.09281524752796096, 32'sd0.05923518753769441, 32'sd-0.03247350357726263, 32'sd-0.013744082778866672, 32'sd0.06875589893410576, 32'sd-0.0540503882477277, 32'sd0.02630545755074627, 32'sd-0.07929621662758277, 32'sd0.03546050774117342, 32'sd0.09330699563663926, 32'sd-0.06851560320102594, 32'sd-0.025422495872124362, 32'sd0.07744263027980178, 32'sd0.0076611435772639324, 32'sd-0.03104387302741692, 32'sd-0.08086981349703684, 32'sd-0.0636933692011259, 32'sd0.10233963498559144, 32'sd0.17460084827907874, 32'sd-0.003359165036202955, 32'sd0.02836769499083967, 32'sd-0.06992085202185608, 32'sd-0.007841616589504212, 32'sd0.04599983956381987, 32'sd0.05930085506478026, 32'sd-0.05244454323535565, 32'sd-0.12950855427104124, 32'sd-0.027675730493040358, 32'sd-0.09897528331106936, 32'sd-0.05262469737674633, 32'sd-0.0071055183011824955, 32'sd-0.048107726849603925, 32'sd-2.626260537778754e-118, 32'sd0.005541584576993771, 32'sd0.06937991397097051, 32'sd0.00223962774366137, 32'sd0.003928632022413794, 32'sd-0.009884671960624333, 32'sd-0.12019587314940422, 32'sd-0.03393670440696905, 32'sd-0.034364452790595836, 32'sd0.09367694603953484, 32'sd-0.06539665079308181, 32'sd-0.060270932992788046, 32'sd-0.07103977182692726, 32'sd0.08538328568773147, 32'sd0.045182910353092305, 32'sd0.10499583734028144, 32'sd0.07411837658280516, 32'sd-0.009713439512047622, 32'sd-0.059469316740166984, 32'sd-0.05375223738252535, 32'sd0.03330831055186679, 32'sd-0.1859814695507301, 32'sd-0.07414462428685853, 32'sd-0.026675193464986847, 32'sd-0.058301327148388746, 32'sd0.023125727989253025, 32'sd0.012338787588230328, 32'sd0.03551725415672036, 32'sd-0.03276108578262679, 32'sd0.029082332284936323, 32'sd0.0979849466730354, 32'sd0.02073884004501753, 32'sd-0.12035685293659364, 32'sd-0.079172687383295, 32'sd-0.02320799853185484, 32'sd-0.016964064071704848, 32'sd0.07891548790642608, 32'sd-0.057365194763541724, 32'sd0.005982307216596693, 32'sd-0.05231253478995118, 32'sd0.09693439580221767, 32'sd0.1805477939168385, 32'sd0.08421725739315827, 32'sd0.09813524099658737, 32'sd-0.10370521637877231, 32'sd-0.0965751500154802, 32'sd-0.13142856222816168, 32'sd-0.09747407783530633, 32'sd-0.1803544597093962, 32'sd-0.12615368318190096, 32'sd-0.15312816710636512, 32'sd-0.01732357333178073, 32'sd-0.05438097397068681, 32'sd0.07342019752542492, 32'sd0.0073435433039726345, 32'sd0.042694733334610234, 32'sd0.06846233486374673, 32'sd-0.007183865454453333, 32'sd-0.05792237608696239, 32'sd-0.04815116544676663, 32'sd-0.009838845814990352, 32'sd-0.03112034105038421, 32'sd-0.0016577653047736049, 32'sd0.015349594269579112, 32'sd0.029638074239572893, 32'sd0.09121735230654962, 32'sd0.006061752042949884, 32'sd-0.045221849406914094, 32'sd0.18496913020439978, 32'sd0.19202166692508932, 32'sd0.11951271360513148, 32'sd-0.003438421483527676, 32'sd-0.08518096224658604, 32'sd-0.19197087374360208, 32'sd-0.20219575732999684, 32'sd-0.11550652030285258, 32'sd-0.12709979772265623, 32'sd-0.26753109926591884, 32'sd-0.19809352810203282, 32'sd-0.16547042904451256, 32'sd0.03340362306958829, 32'sd0.04577991624176015, 32'sd0.06260780724444943, 32'sd0.03666371630827116, 32'sd-2.209232632768596e-126, 32'sd-0.008152436224862551, 32'sd-0.11918883181392996, 32'sd-0.11019758682460021, 32'sd-0.09283917347889879, 32'sd0.06753108211691557, 32'sd-0.021701485586555724, 32'sd-0.08496865084362856, 32'sd-0.020581693516857832, 32'sd-0.07166742565000876, 32'sd0.044959082652579856, 32'sd0.032687043006506794, 32'sd0.06710859589513493, 32'sd0.14879906681736937, 32'sd0.0530002335065644, 32'sd-0.1255533534295686, 32'sd-0.17156923505779553, 32'sd-0.12528634802510494, 32'sd-0.07824037697733457, 32'sd0.007337908891475937, 32'sd-0.15762895808315533, 32'sd-0.13911337525910455, 32'sd-0.1622660346214274, 32'sd-0.11341288068338796, 32'sd-0.0032064760833888104, 32'sd-0.031234231875722853, 32'sd0.05045510458253292, 32'sd0.06133989846087161, 32'sd0.02147386171883721, 32'sd0.03622723980405154, 32'sd-0.10210589814821455, 32'sd-0.036801907000297465, 32'sd-0.052604843685946895, 32'sd0.025761559814849698, 32'sd-0.018406831977703576, 32'sd0.0738379677102153, 32'sd0.06086962299636383, 32'sd0.0427974238458003, 32'sd0.04968179186807571, 32'sd0.09559657715628968, 32'sd0.12306343193956154, 32'sd0.05290601599596365, 32'sd0.09698877180378383, 32'sd-0.12223104268042194, 32'sd-0.09205129532763977, 32'sd-0.04844172284208175, 32'sd-0.1233985244159759, 32'sd-0.10401744159770304, 32'sd-0.02492906368719034, 32'sd-0.03297038031710286, 32'sd-0.08924260754257904, 32'sd0.017648950244523003, 32'sd0.07463002038534586, 32'sd-0.04774428648887581, 32'sd-0.031166311607220283, 32'sd0.04879138577161311, 32'sd0.11428177185954908, 32'sd0.09625891423406183, 32'sd-0.09432843689649763, 32'sd-0.0038544209212592324, 32'sd-0.09500309690270105, 32'sd0.003496852666355169, 32'sd0.02438393239862297, 32'sd-0.004093421407949992, 32'sd0.06304343657354539, 32'sd0.09997326946099379, 32'sd0.09147240308840883, 32'sd0.049512879816812475, 32'sd0.057605687016958514, 32'sd0.15425668223854413, 32'sd-0.001002060128099629, 32'sd-0.061913242568316866, 32'sd-0.18435248125188466, 32'sd-0.10092910296729304, 32'sd-0.04854476961973224, 32'sd-0.07085514913336348, 32'sd-0.048877860241346605, 32'sd0.03111033607551109, 32'sd0.056435390699150045, 32'sd0.010506276656105809, 32'sd-0.0072386135114578185, 32'sd0.0002487323306826591, 32'sd0.018769845555706783, 32'sd0.07434170702515965, 32'sd-1.1687507888867274e-122, 32'sd0.08615936749617202, 32'sd-0.0322121841312765, 32'sd-0.13430953308083884, 32'sd-0.02017157017471895, 32'sd-0.014985540022621697, 32'sd-0.013115750989582125, 32'sd-0.04688110426508055, 32'sd-0.06954418784392778, 32'sd-0.019747070107634407, 32'sd0.010731823482356483, 32'sd0.00802151476336999, 32'sd0.059549536699014534, 32'sd-0.06528306039282607, 32'sd-0.11055040279184887, 32'sd-0.12392583151732327, 32'sd-0.14159151956787705, 32'sd-0.1339087317528531, 32'sd-0.12366211521660528, 32'sd-0.1182042651174091, 32'sd0.042455447341809956, 32'sd-0.10760532726188657, 32'sd-0.03847310771692925, 32'sd-0.05349089405878009, 32'sd0.0242059987012528, 32'sd0.07380504860547377, 32'sd0.0017938180767866523, 32'sd4.942360448898085e-118, 32'sd6.68772906165591e-122, 32'sd-8.117203838198642e-121, 32'sd-0.03992404731197002, 32'sd0.031217650823269737, 32'sd-0.008526787604430177, 32'sd0.04188095894704925, 32'sd0.059521772560132025, 32'sd-0.006054207001393125, 32'sd-0.012086187726825532, 32'sd0.025788704455375008, 32'sd-0.019417510786591985, 32'sd0.04693124190106233, 32'sd0.0280535850409639, 32'sd-0.1749047914763649, 32'sd-0.061210057307732706, 32'sd0.009299910431874968, 32'sd-0.07093801065916233, 32'sd-0.08421463329671167, 32'sd-0.1615740751766747, 32'sd-0.16666151611495597, 32'sd-0.0387812705813473, 32'sd-0.03245946706588668, 32'sd-0.022262849891968597, 32'sd-0.013442325953060023, 32'sd-0.023915315585783272, 32'sd-0.06684245658736009, 32'sd0.032413475628630964, 32'sd2.6930862525392837e-116, 32'sd-2.5838571685709903e-117, 32'sd2.2387149104645477e-124, 32'sd-0.022760612049022813, 32'sd0.03918843529343394, 32'sd-0.04588532059651108, 32'sd0.04785566577521594, 32'sd-0.048500361774919114, 32'sd0.057051802719679405, 32'sd0.04856116018027569, 32'sd0.08705668067948828, 32'sd0.05123303736382474, 32'sd0.0010896837292881036, 32'sd-0.04979900523948376, 32'sd-0.09600298478502117, 32'sd0.0467375969364655, 32'sd0.13498458894972215, 32'sd-0.009842178330543083, 32'sd-0.02552850277278155, 32'sd-0.11552702409005848, 32'sd-0.11732257278887678, 32'sd-0.006127530991627108, 32'sd-0.03868973491896021, 32'sd0.040833268591163735, 32'sd0.05689526601544686, 32'sd-0.05338889412596711, 32'sd-0.02303777786646724, 32'sd0.0133204217609093, 32'sd5.831503288718107e-122, 32'sd3.0854178090375254e-129, 32'sd3.196399643670589e-122, 32'sd-5.087602893179534e-124, 32'sd0.12960237522726417, 32'sd-0.10430505178611017, 32'sd-0.06697176894733681, 32'sd-0.009109857303242807, 32'sd0.06871803548994991, 32'sd0.0018416561687512466, 32'sd-0.005185957851995338, 32'sd0.02156205580984296, 32'sd0.09116646145413863, 32'sd-0.014079071675506321, 32'sd0.07516673728799668, 32'sd-0.028587949774019246, 32'sd-0.007996428826316054, 32'sd-0.018166198748998982, 32'sd0.11907576812369776, 32'sd0.06671148970253066, 32'sd-0.03380349742245673, 32'sd0.07180143865209115, 32'sd-0.044986146503187524, 32'sd0.06469057634179814, 32'sd-0.0008416089051896817, 32'sd0.10964455600618331, 32'sd0.07998878449386747, 32'sd-3.7171782174218667e-118, 32'sd-2.4331104557156575e-121, 32'sd9.680366856857106e-129, 32'sd-3.6202872538695285e-120, 32'sd-1.9686744127566442e-117, 32'sd2.0675746269336544e-118, 32'sd0.06180763871869473, 32'sd-0.048038689129495445, 32'sd0.07520376879904503, 32'sd0.019799310693745627, 32'sd-0.07762061022549802, 32'sd0.007375285550991771, 32'sd0.06042417959648282, 32'sd-0.01012973318539873, 32'sd0.09570175373726837, 32'sd0.09130470606120308, 32'sd0.057422768721267184, 32'sd0.004515193743727296, 32'sd0.09002351550872732, 32'sd0.01173058509857688, 32'sd-0.038210512976330144, 32'sd0.01749309588042752, 32'sd0.08493482490429176, 32'sd-0.024851440737796802, 32'sd-0.002952182612347003, 32'sd0.10756360272932648, 32'sd-4.597135349040434e-115, 32'sd-1.4231398098466445e-118, 32'sd-3.2229678705468966e-120, 32'sd2.61684718194673e-126},
        '{32'sd-3.680645934372999e-122, 32'sd-2.4192601656838826e-126, 32'sd-7.308043781791256e-115, 32'sd-4.6720756724052454e-122, 32'sd1.5432478468842584e-122, 32'sd1.9267156098796475e-118, 32'sd-1.3255918982322644e-118, 32'sd3.6426348791025785e-122, 32'sd-1.757125166593357e-123, 32'sd-4.3939351132173514e-123, 32'sd-3.188377110810069e-120, 32'sd3.549392397955086e-116, 32'sd-0.0725939889910267, 32'sd0.023471938215388177, 32'sd0.053083124955158684, 32'sd0.1035179396453052, 32'sd-4.039800365361871e-118, 32'sd-5.5214458667159645e-121, 32'sd6.588071854858927e-125, 32'sd-3.3119136026003745e-121, 32'sd-8.842423459389303e-127, 32'sd-1.5351524492940738e-127, 32'sd9.068067891801043e-121, 32'sd2.849953041478145e-120, 32'sd6.8152455631615e-127, 32'sd-1.4811407147875736e-115, 32'sd-1.3175284924692184e-122, 32'sd-1.3246633802902327e-126, 32'sd-2.0215232174003742e-117, 32'sd1.073661736460248e-119, 32'sd-8.79394841933316e-122, 32'sd-1.7356870346232147e-120, 32'sd0.028463016055892652, 32'sd-0.0027117504001971304, 32'sd-0.02411398881217488, 32'sd-0.017491804916671124, 32'sd0.07493728005079915, 32'sd-0.08133018349939651, 32'sd0.03323693411700166, 32'sd-0.08752645904107136, 32'sd0.04187414030740971, 32'sd-0.0785076994673189, 32'sd0.11041110570771524, 32'sd0.034734033964762163, 32'sd-0.004955045149200142, 32'sd0.08112282668493125, 32'sd-0.060079263836253026, 32'sd-0.010663101591807854, 32'sd-0.00011833975052088545, 32'sd0.0028014476574873244, 32'sd0.012464121829015176, 32'sd0.06259297019429762, 32'sd1.6517181455303457e-121, 32'sd-1.850248265342111e-122, 32'sd-2.462942048859107e-124, 32'sd-4.351081866331739e-126, 32'sd-1.296041527214297e-125, 32'sd-1.1491388580978908e-125, 32'sd0.04431490717942538, 32'sd-0.05463464401608574, 32'sd0.022364773848823113, 32'sd-0.025279173287249754, 32'sd-0.05193818184140129, 32'sd-0.06020987474172419, 32'sd-0.07365528166460113, 32'sd-0.03424239095618862, 32'sd0.1038569296860312, 32'sd0.04539728917461952, 32'sd0.0014115122241238481, 32'sd0.03268672057051598, 32'sd0.05230773547433312, 32'sd-0.08225294450993392, 32'sd0.033163704738313884, 32'sd0.022461282574542735, 32'sd-0.023542985822501142, 32'sd0.1486376801091382, 32'sd0.0925897536052746, 32'sd-0.027286233299327733, 32'sd0.08676223475717078, 32'sd-0.065796817904268, 32'sd0.07242994827707223, 32'sd0.08986291675406927, 32'sd3.4664935674684363e-122, 32'sd2.1724380889459054e-126, 32'sd-5.151643006542765e-116, 32'sd3.239608653590663e-115, 32'sd0.06862682797310099, 32'sd0.0587511885112907, 32'sd-0.042744314015046185, 32'sd0.019232942631143418, 32'sd0.04480451533946008, 32'sd-0.0496366834696899, 32'sd0.09830192506109856, 32'sd0.0564305480745071, 32'sd-0.08974607248139928, 32'sd0.06459926388877472, 32'sd-0.14055704080876427, 32'sd-0.1659623781689404, 32'sd-0.016519915201901388, 32'sd-0.046659992453869994, 32'sd-0.0032473129751718448, 32'sd0.0998671185044918, 32'sd0.048994998459795, 32'sd0.04351105828541196, 32'sd0.09542195853136651, 32'sd0.03039465011902044, 32'sd0.02818250625674663, 32'sd-0.028131531130462333, 32'sd-0.08145930613914378, 32'sd-0.052639716332622655, 32'sd0.03784639572228236, 32'sd5.15018709462407e-124, 32'sd4.838907959316874e-123, 32'sd0.1006935555737055, 32'sd-0.007172395057880745, 32'sd0.03785674274902104, 32'sd0.0470639769184368, 32'sd0.0032746497361386844, 32'sd0.003834291186645071, 32'sd0.0034548268539120017, 32'sd-0.0604869351386028, 32'sd-0.06078119538331984, 32'sd-0.017274617374219377, 32'sd-0.021268997892119876, 32'sd-0.07298165267074887, 32'sd-0.03212386770911395, 32'sd-0.009582080795118726, 32'sd0.05317562713474906, 32'sd0.07745088389376986, 32'sd0.041032966793050976, 32'sd0.06242525669161196, 32'sd0.06676017001236245, 32'sd0.05802666172282738, 32'sd0.10207910180903616, 32'sd0.06097714195491449, 32'sd-0.022395414067414993, 32'sd-0.039467922433773686, 32'sd-0.006064889295694174, 32'sd-0.0599943382695309, 32'sd0.08039835540057251, 32'sd1.9486540737414315e-126, 32'sd0.102600441462927, 32'sd-0.061313584608427486, 32'sd0.08675701765014474, 32'sd0.033269592110709754, 32'sd-0.056334071540869037, 32'sd0.020923593539122484, 32'sd-0.008012054404558029, 32'sd0.008195070735632838, 32'sd0.04734586625521679, 32'sd0.05494742051340673, 32'sd0.0023275548960354654, 32'sd0.12555117285059594, 32'sd0.05366060102912175, 32'sd-0.08140601106165518, 32'sd-0.07076646848354597, 32'sd0.08469211206231726, 32'sd0.14624513066017514, 32'sd0.03985053616836902, 32'sd-0.025197152958262505, 32'sd0.003843485144374853, 32'sd0.01209939740832132, 32'sd-0.12422940904408344, 32'sd-0.05166832466672733, 32'sd-0.021285522822883495, 32'sd-0.007771657524600894, 32'sd0.014575198956250037, 32'sd-0.08059517939192835, 32'sd-8.063313218751297e-126, 32'sd0.04516527482322174, 32'sd0.08794558228465713, 32'sd-0.06109700415471549, 32'sd0.040086721282441555, 32'sd0.04830467519928358, 32'sd0.05327948517835776, 32'sd0.08766652780045663, 32'sd0.005553335851547478, 32'sd0.003536033792977909, 32'sd-0.06743126861134491, 32'sd-0.08143077655614424, 32'sd0.0826895461217271, 32'sd-0.10336703382226993, 32'sd-0.04282033765476297, 32'sd-0.10314649872216673, 32'sd0.10157867310139788, 32'sd0.1234679407384605, 32'sd0.10951304814440307, 32'sd0.14755458878153313, 32'sd-0.016979350373425395, 32'sd-0.07973982148095053, 32'sd-0.06590887256729669, 32'sd0.020323960026545303, 32'sd-0.05942824601498855, 32'sd0.00904629811562161, 32'sd-0.027155229958350596, 32'sd0.036744253425367426, 32'sd0.051017069086423644, 32'sd0.03680706295857111, 32'sd-0.05418381223458231, 32'sd-0.03524842024336896, 32'sd0.0804321502897702, 32'sd0.04594431079416248, 32'sd0.13058111189755447, 32'sd0.21413067875912464, 32'sd0.09691819880836076, 32'sd0.005377656673565235, 32'sd0.026582196566916915, 32'sd-0.10622403220779357, 32'sd-0.10419851875725407, 32'sd-0.15274224290209415, 32'sd-0.2666480973957614, 32'sd-0.10784624154322016, 32'sd-0.010199046423243867, 32'sd0.17437985974520953, 32'sd0.185083164591224, 32'sd0.08545809158985386, 32'sd-0.11320072577136886, 32'sd-0.09924794076954634, 32'sd-0.06768411358927284, 32'sd-0.14877067818583756, 32'sd-0.03389931708251792, 32'sd0.11446661616961776, 32'sd-0.0382453768305078, 32'sd0.03128143873538974, 32'sd0.004136700970164897, 32'sd0.052295316654836214, 32'sd0.05169687252563798, 32'sd0.06982646672825853, 32'sd-0.027180136506290857, 32'sd0.0331464147191457, 32'sd0.004217219968116369, 32'sd0.135152775963449, 32'sd0.050725026935627714, 32'sd0.13597388976084215, 32'sd0.012855959933487173, 32'sd-0.09585587679618915, 32'sd-0.03743232493347323, 32'sd-0.133668362812765, 32'sd-0.2654923218947089, 32'sd-0.11011847179826713, 32'sd0.12207395628800746, 32'sd0.2134902134715274, 32'sd0.07506993426845757, 32'sd-0.0939075955141506, 32'sd-0.20897918155130396, 32'sd-0.2778832921275319, 32'sd-0.12295605295956934, 32'sd-0.017903274847000307, 32'sd0.07505832167924781, 32'sd0.12374094638918264, 32'sd0.09604525201416558, 32'sd0.013691507211556198, 32'sd-0.019928528808046703, 32'sd0.059327543748615374, 32'sd0.013555240208289989, 32'sd-0.026276288845953163, 32'sd0.054370742939462355, 32'sd0.08814557331195282, 32'sd0.06377797649182532, 32'sd0.07846052670459817, 32'sd0.08539958120994666, 32'sd-0.036571755118397005, 32'sd-0.024888062082075134, 32'sd0.06237864000445128, 32'sd0.04966499605059518, 32'sd-0.09205805760247882, 32'sd-0.020062721132082875, 32'sd0.13422920069328453, 32'sd0.32510173246562346, 32'sd0.2538454489236342, 32'sd0.07002370273522604, 32'sd-0.2133873375955567, 32'sd-0.23559479865583832, 32'sd-0.19454799754011362, 32'sd0.009345113370681288, 32'sd0.06027393951890806, 32'sd-0.0032492743413624426, 32'sd0.06129878615060669, 32'sd-0.060332968857504, 32'sd0.003504372056696265, 32'sd0.09363681670538589, 32'sd0.061291582132367475, 32'sd-0.021799223279624906, 32'sd-0.026373404975126743, 32'sd0.0743628102269735, 32'sd-0.09480198289423526, 32'sd0.05402526471656251, 32'sd0.08645387666112209, 32'sd0.09516481001812906, 32'sd-0.00443483037076472, 32'sd-0.039110691887063675, 32'sd0.08182596197103546, 32'sd0.025096318987189514, 32'sd0.012650995978686708, 32'sd0.05640898724253461, 32'sd0.142333582064828, 32'sd0.25180897663671886, 32'sd0.10013163381746222, 32'sd-0.15404007163811734, 32'sd-0.25775881686334046, 32'sd-0.13275236896214268, 32'sd-0.12037856139033572, 32'sd0.02190556056714742, 32'sd0.1587783642419583, 32'sd-0.13968566051293607, 32'sd0.06772729039590164, 32'sd0.06270719508325945, 32'sd0.019588396457072516, 32'sd0.11297075548850817, 32'sd0.009257245100149834, 32'sd-0.06955931669974702, 32'sd0.01206992389653486, 32'sd0.0816515799078107, 32'sd0.06663259445168382, 32'sd-0.03738106948120362, 32'sd-0.04037936589564802, 32'sd0.12017469793063898, 32'sd0.07591194239996926, 32'sd0.05620378180765421, 32'sd0.10771494674341674, 32'sd0.08788282974706313, 32'sd0.06877967946677904, 32'sd0.1613975510654218, 32'sd0.21283201406763083, 32'sd0.10541106002042028, 32'sd-0.13628191481061402, 32'sd-0.24881958178881405, 32'sd-0.17928201561011556, 32'sd-0.07073052254257117, 32'sd-0.016330770574073613, 32'sd-0.001437677324838711, 32'sd0.025377803768192972, 32'sd-0.16439865631604247, 32'sd0.006407284868308436, 32'sd-0.06974703734579915, 32'sd-0.023760941914488402, 32'sd0.03457068158602725, 32'sd0.0202710210765715, 32'sd0.08949577501296849, 32'sd-0.025639724773280085, 32'sd0.021425286430351728, 32'sd0.0725527524039998, 32'sd0.06711191308477366, 32'sd0.037846738004832264, 32'sd0.05567994720159233, 32'sd0.06535146014151741, 32'sd0.30409833043362733, 32'sd0.16133242776345083, 32'sd0.0947956039349589, 32'sd0.021214000067524722, 32'sd0.03614249617082022, 32'sd0.10393605402402878, 32'sd0.07337943418612985, 32'sd-0.11372129690186807, 32'sd-0.14498854999953673, 32'sd-0.03182933676135404, 32'sd0.002019342367652047, 32'sd0.020484396421140885, 32'sd-0.002624941673381775, 32'sd0.04787242437468172, 32'sd-0.017791605116034077, 32'sd0.014621526920930888, 32'sd-0.10574341505122965, 32'sd-0.009569535636759587, 32'sd0.052548327585641694, 32'sd-0.022265830862935536, 32'sd0.10224482619888663, 32'sd-0.07749177208507531, 32'sd-0.10319106053870782, 32'sd0.012653232224505226, 32'sd-0.030113117485996484, 32'sd0.018542574253699446, 32'sd0.07847102497977165, 32'sd0.12144476661568988, 32'sd0.029052554262908935, 32'sd0.08680493072889223, 32'sd0.011951850764502791, 32'sd0.02964904007379539, 32'sd0.03253200821115301, 32'sd0.06437703080969645, 32'sd0.008687047679800936, 32'sd-0.04672821757570873, 32'sd0.08863804425432886, 32'sd-0.03774953779696755, 32'sd0.11671560350555255, 32'sd0.033092977670598815, 32'sd-0.06122327007036262, 32'sd0.02208352623038291, 32'sd0.07803393106102754, 32'sd0.14299296361844308, 32'sd0.042567206447148204, 32'sd-0.02110845796669315, 32'sd-0.009780264429293865, 32'sd0.049873966466264866, 32'sd0.021435829499393586, 32'sd-0.00771532163690864, 32'sd-0.027657272279156455, 32'sd0.022827547562495148, 32'sd-0.027240638255271413, 32'sd-0.09390827386135901, 32'sd0.004155857708580359, 32'sd-0.06015121654883272, 32'sd-0.07530500891325748, 32'sd0.022804977161293687, 32'sd0.01268898248874421, 32'sd0.1699876186870432, 32'sd0.11487350805162355, 32'sd0.10604421924544026, 32'sd-0.04294225151760842, 32'sd-0.15016178141687983, 32'sd-0.0007831898215903877, 32'sd0.11626659608750713, 32'sd-0.05970592002998117, 32'sd0.027638035508620585, 32'sd0.07132911102337999, 32'sd-0.014724323147368674, 32'sd-0.0575452363416723, 32'sd-0.021148840520444266, 32'sd0.047721693079396825, 32'sd0.04280933039968513, 32'sd0.05696574251867198, 32'sd0.07959660627547469, 32'sd0.03104069025992529, 32'sd0.029891924055008498, 32'sd-0.06740218096013924, 32'sd-0.05710168774354185, 32'sd0.07074004601563358, 32'sd-0.03146331191651169, 32'sd-0.160290420718354, 32'sd-0.142035647961079, 32'sd-0.09990264264300214, 32'sd0.0072650414083164335, 32'sd-0.08558644835525811, 32'sd-0.020020502204912145, 32'sd0.08529424284051673, 32'sd0.22401947378795392, 32'sd0.03694934266461647, 32'sd-0.04874796977416817, 32'sd-0.017260011433281215, 32'sd-0.05989405147434525, 32'sd0.07193977267421692, 32'sd-0.025156920341417532, 32'sd0.10532572865845605, 32'sd-0.01985387991096868, 32'sd-0.033939661168648175, 32'sd-0.10577914626757992, 32'sd0.045820634060746185, 32'sd-0.004805943467964421, 32'sd0.07662229369885126, 32'sd0.07289555868518244, 32'sd-0.04326721552233698, 32'sd-0.06134345862062269, 32'sd-0.12596196164250545, 32'sd0.032357370060714506, 32'sd0.12170424667089366, 32'sd0.08320855953585665, 32'sd-0.0899755631451792, 32'sd-0.07332736513663782, 32'sd0.06335608722304197, 32'sd0.03940566649889573, 32'sd0.028229761233433175, 32'sd-0.0024297931061455823, 32'sd-0.02861358695775956, 32'sd0.19518373129479025, 32'sd-0.11280158982051025, 32'sd-0.002454791071895001, 32'sd0.028185600325560677, 32'sd-0.05287184394553775, 32'sd-0.02397126278001506, 32'sd0.05643493675442371, 32'sd0.010029616282883479, 32'sd-0.009102161901995559, 32'sd-0.023671567447524265, 32'sd-0.10506208016692867, 32'sd0.0015589545828166313, 32'sd-0.04131297445173881, 32'sd-1.5668623615822834e-123, 32'sd-0.03711285782073747, 32'sd0.0037873585833320617, 32'sd-0.09341656107807068, 32'sd0.05952306915502329, 32'sd0.07080575011800827, 32'sd-0.10126012292928513, 32'sd0.03807859769492146, 32'sd-0.030027282357287268, 32'sd0.03813744382597404, 32'sd-0.03795961856499812, 32'sd-0.08997204306959192, 32'sd-0.06526128140569072, 32'sd0.07415483723242076, 32'sd0.0021830443733294467, 32'sd0.02286686271036259, 32'sd-0.01629981938993848, 32'sd0.0806029657788623, 32'sd-0.08855520509103956, 32'sd-0.0018597515298829025, 32'sd-0.05358143053085661, 32'sd0.12034652245931833, 32'sd0.11652595131699688, 32'sd0.00947117753761832, 32'sd0.11267204967410589, 32'sd-0.12194257973956801, 32'sd0.02902785480200253, 32'sd0.05314676782441744, 32'sd0.0722584766851085, 32'sd0.07696530670209537, 32'sd-0.10960726011367974, 32'sd-0.07854770191003246, 32'sd0.061531497396638345, 32'sd0.02364951897881128, 32'sd-0.014049230064317983, 32'sd-0.085434750903013, 32'sd0.048707296266445536, 32'sd-0.04100263952291798, 32'sd-0.04356190724463249, 32'sd-0.09258364475585135, 32'sd-0.08339343048930607, 32'sd-0.09259196994260664, 32'sd0.007768716361075981, 32'sd-0.08916308319698081, 32'sd-0.12782354842721708, 32'sd0.02585788617093864, 32'sd0.03675012112889228, 32'sd0.06084976765652247, 32'sd0.11396125179805312, 32'sd0.11616492523951136, 32'sd0.01962453762317296, 32'sd0.015728640931407703, 32'sd0.11235409310435292, 32'sd-0.06872199488011549, 32'sd-0.02412538799830895, 32'sd0.011543953996600737, 32'sd0.019602061701811113, 32'sd0.06742330377293203, 32'sd-0.05801544526682443, 32'sd0.12022915547023766, 32'sd0.059860691668746094, 32'sd-0.026000453484550164, 32'sd-0.027595465699118596, 32'sd-0.0038944570157412968, 32'sd0.03726215611456873, 32'sd0.07199784210322704, 32'sd0.008225086391219159, 32'sd-0.028393073149962464, 32'sd-0.1400492260174072, 32'sd-0.1213231098985117, 32'sd-0.08371490204342821, 32'sd-0.22199334081120878, 32'sd-0.03463119218006872, 32'sd-0.03091914587701901, 32'sd0.07357821885208245, 32'sd0.02156585746746666, 32'sd0.04006365368084306, 32'sd0.1075822166208295, 32'sd-0.0028465157667235523, 32'sd-0.052861724908030275, 32'sd0.09651442093468575, 32'sd0.033703047935144434, 32'sd-0.09539100609382535, 32'sd-0.06158711224257343, 32'sd8.023012853387228e-120, 32'sd-0.02250553264891869, 32'sd-0.02549811693250724, 32'sd0.0981994069019147, 32'sd-0.05259932407735718, 32'sd-0.1120408126836354, 32'sd0.06354382201586062, 32'sd0.05501784744855737, 32'sd-0.01351745524075084, 32'sd-0.05550295362663794, 32'sd0.01323330938184828, 32'sd0.013083147279243913, 32'sd-0.04875722984429853, 32'sd-0.03915605172218322, 32'sd0.024191507225215937, 32'sd-0.012897537180530997, 32'sd-0.022159484599111604, 32'sd0.006220436980078913, 32'sd0.07033207731752918, 32'sd0.01818567283042255, 32'sd-0.0531642051903821, 32'sd-0.03391349955171753, 32'sd-0.05461270065125836, 32'sd0.044679561561814095, 32'sd0.06923008097986066, 32'sd-0.023115177584058434, 32'sd0.027945276687407993, 32'sd0.029939728380654094, 32'sd0.10964757222497078, 32'sd0.017763768262879998, 32'sd0.014760768424943373, 32'sd-0.00551243906846041, 32'sd-0.14404384038890067, 32'sd-0.11631454567786396, 32'sd-0.09701758180859654, 32'sd-0.025738823886136197, 32'sd-0.10178723301360788, 32'sd-0.028205022647004203, 32'sd-0.0068253272058828775, 32'sd0.03558166707127169, 32'sd-0.07039792218563597, 32'sd0.013733594807461487, 32'sd-0.040302773488741166, 32'sd-0.003847264041954057, 32'sd0.017806308217695112, 32'sd-0.07055197749495279, 32'sd0.07332474920097969, 32'sd-0.06701941866939443, 32'sd0.039603912615430774, 32'sd-0.062306278343389976, 32'sd0.01908610945763199, 32'sd-0.03611474831527255, 32'sd-0.03157250419255895, 32'sd0.0771463586681776, 32'sd-0.07759811935153756, 32'sd-0.0322599711057171, 32'sd-0.0062242795060857255, 32'sd0.1242128017006386, 32'sd-0.05409686052427519, 32'sd-0.014913140700071468, 32'sd0.0005592470094620248, 32'sd-0.021216185120214108, 32'sd-0.05659796955935361, 32'sd-0.09503320183887669, 32'sd-0.021936557412119043, 32'sd0.03133162281797507, 32'sd0.03861365163305581, 32'sd-0.07022983305255527, 32'sd-0.018535468584078608, 32'sd-0.05690110932977197, 32'sd-0.07631567689317184, 32'sd-0.004351199772441689, 32'sd0.023956835705747304, 32'sd-0.003231757789830523, 32'sd-3.590811813345023e-05, 32'sd0.10788149802816056, 32'sd0.07744594338519746, 32'sd-0.0646757486650606, 32'sd0.014790908439843257, 32'sd-0.04776542615678333, 32'sd0.10410250319271751, 32'sd0.06355038123519562, 32'sd0.012713799333576695, 32'sd0.04048410413049217, 32'sd2.3989908619714055e-125, 32'sd-0.022585944025925526, 32'sd0.05671148336365255, 32'sd0.06796662976556417, 32'sd-0.014149851855361936, 32'sd0.003264775811532458, 32'sd-0.041709697061859376, 32'sd0.07328915416537518, 32'sd0.09898152208892938, 32'sd0.057860574242292524, 32'sd0.13526075273052496, 32'sd-0.05946668879015078, 32'sd-0.1433900097405783, 32'sd-0.012605418334287029, 32'sd-0.06613078777806257, 32'sd0.010219668437517423, 32'sd-0.011119443179592544, 32'sd-0.06893426877205754, 32'sd0.07780790423024937, 32'sd0.07668763157092044, 32'sd-0.05835976594633175, 32'sd-0.027844788091206368, 32'sd0.0573588138019606, 32'sd0.10383656782419795, 32'sd-0.008177074017661089, 32'sd-0.042911832613353566, 32'sd-0.025703610619969588, 32'sd5.783064983818818e-119, 32'sd2.352460545330624e-120, 32'sd-1.9133396512794714e-126, 32'sd0.010127386268024147, 32'sd0.050972492663840255, 32'sd0.05052818143370817, 32'sd-0.0849876576254581, 32'sd-0.0027168119846423043, 32'sd0.04984633307925561, 32'sd-0.0418985234616354, 32'sd0.048454851482607086, 32'sd-0.02346586736047226, 32'sd0.05806258074955395, 32'sd-0.05189527187256973, 32'sd0.004986993846176302, 32'sd0.09486672666643056, 32'sd-0.08116910699206786, 32'sd-0.07603359279958455, 32'sd-0.0723251691373672, 32'sd-0.0061772033202778945, 32'sd0.04559169775459848, 32'sd-0.053438353369961264, 32'sd-0.01568508585686799, 32'sd0.06911277224680507, 32'sd0.0033778305846879964, 32'sd0.024299617943936664, 32'sd0.01184306221627935, 32'sd0.014808038833259944, 32'sd-3.7470464824125794e-122, 32'sd3.0525766594479214e-119, 32'sd-1.416751612358028e-127, 32'sd0.013988270738010934, 32'sd-0.002060553001846279, 32'sd-0.037697279975964906, 32'sd-0.11575429026487544, 32'sd0.09821360622236085, 32'sd0.016069101019723152, 32'sd-0.01717524256463651, 32'sd-0.0026875001104448, 32'sd-0.021403808947345223, 32'sd-0.015437686495931236, 32'sd0.036324104786301784, 32'sd0.023310132890488486, 32'sd-0.07534878945344667, 32'sd-0.00660683558810454, 32'sd-0.010444000260921908, 32'sd-0.024371251265149555, 32'sd0.06559274634587194, 32'sd-0.013664300416989699, 32'sd-0.06355519646701152, 32'sd0.03880983437251949, 32'sd-0.01984736630595264, 32'sd-0.014962765744167703, 32'sd0.05908088958560397, 32'sd0.0210648154674399, 32'sd0.061023799467551224, 32'sd-6.734148812855605e-124, 32'sd1.2464116903185513e-114, 32'sd-8.885581220254278e-127, 32'sd6.15645269369444e-123, 32'sd0.017592875004571865, 32'sd-0.03082547605185195, 32'sd-0.002576571883903134, 32'sd0.04991743254190567, 32'sd0.054885539866074896, 32'sd-0.03643283194749983, 32'sd-0.16258632732129585, 32'sd0.06700643415627508, 32'sd0.024438446438329518, 32'sd0.009594716946892684, 32'sd0.036497252607757706, 32'sd0.11428923233548913, 32'sd-0.04236010969560328, 32'sd-0.045664389281595615, 32'sd-0.1761250918128987, 32'sd-0.09053822431827255, 32'sd0.043781365140027846, 32'sd-0.08214558943000931, 32'sd0.04203292004922413, 32'sd-0.0424498416833081, 32'sd0.0038879387167629004, 32'sd0.02354321901849888, 32'sd0.06875333081035202, 32'sd-1.2678006399127925e-119, 32'sd-2.8308852727218216e-121, 32'sd3.3453398261024517e-122, 32'sd1.076497973964867e-124, 32'sd1.952067913280788e-126, 32'sd4.463344391912334e-118, 32'sd0.04008353910406047, 32'sd0.06266146457395123, 32'sd0.0854474774821785, 32'sd0.04174877109153132, 32'sd-0.04761501783078293, 32'sd0.0021560647829689545, 32'sd-0.02451962925686552, 32'sd0.0038557949058738764, 32'sd-0.009287714069053142, 32'sd-0.04326831577681453, 32'sd0.07097074480153706, 32'sd0.033549067017706186, 32'sd-0.001919905411799906, 32'sd-0.028117696937344148, 32'sd0.060736096726108954, 32'sd-0.04224138150119986, 32'sd0.0032830929085479917, 32'sd-0.015709051602907725, 32'sd0.05543910267782303, 32'sd0.10885966090957759, 32'sd-4.136986301486286e-116, 32'sd3.457176510479951e-121, 32'sd1.0161327995334252e-119, 32'sd-6.802481524832318e-124},
        '{32'sd-1.0395107965503844e-118, 32'sd5.258781404700007e-117, 32'sd-8.534916024215049e-124, 32'sd1.123676188259247e-119, 32'sd1.0704969294599718e-121, 32'sd-6.249022744267372e-126, 32'sd-1.374464016790699e-127, 32'sd-1.7663306398281935e-123, 32'sd-8.574413559437695e-117, 32'sd2.2926174732982097e-124, 32'sd-6.057090190112619e-124, 32'sd1.1690359974495381e-122, 32'sd0.047484941226729444, 32'sd0.12087666584825082, 32'sd0.043437438382863944, 32'sd0.06107759194334618, 32'sd1.3279710577350035e-122, 32'sd1.9291760837574897e-123, 32'sd-5.045501391216145e-115, 32'sd3.574929221240849e-119, 32'sd-3.138617936347068e-119, 32'sd2.5556409711084496e-126, 32'sd1.9053490635733343e-127, 32'sd-2.2908772262606285e-122, 32'sd1.3714042984561976e-121, 32'sd1.643255002153652e-117, 32'sd-7.18246477582648e-126, 32'sd-2.4682934557957246e-124, 32'sd1.0598324160475968e-124, 32'sd-6.2085706157686285e-124, 32'sd2.5022522052977288e-124, 32'sd-2.7424262853014177e-120, 32'sd0.06796760246199712, 32'sd0.0876670497755693, 32'sd-0.022737169136250054, 32'sd-0.03273849915110156, 32'sd-0.01739521221353131, 32'sd-0.1487569682972703, 32'sd-0.04945744271163366, 32'sd-0.013975256380148054, 32'sd0.08582641313373832, 32'sd0.12661261460361548, 32'sd-0.03988029856228843, 32'sd0.025025090891148107, 32'sd-0.007910866731104119, 32'sd0.029138734125208413, 32'sd0.07726448475578815, 32'sd0.05391972573359876, 32'sd0.02122519215827899, 32'sd0.12398921140666234, 32'sd-0.02061285541946961, 32'sd0.07226669303755123, 32'sd-3.355427127604455e-119, 32'sd-2.207006979543644e-118, 32'sd2.990579334479568e-119, 32'sd-4.538938712202444e-123, 32'sd1.9897093024484758e-120, 32'sd-3.494958478170528e-122, 32'sd0.07144884357357136, 32'sd0.06758726712376405, 32'sd0.05885159300782389, 32'sd-0.022816453161839344, 32'sd0.029092059579700905, 32'sd-0.0851414206137923, 32'sd-0.021718372192124615, 32'sd-0.09486466798265156, 32'sd-0.12222908180058625, 32'sd0.05361155613878372, 32'sd0.05077371791305481, 32'sd0.06931485651336475, 32'sd0.08866667233886337, 32'sd-0.013736859933820704, 32'sd0.01036129133819325, 32'sd0.08739470763955072, 32'sd-0.01912382847090221, 32'sd0.011880425460606761, 32'sd0.06888190816573998, 32'sd0.11881265778883277, 32'sd0.1379125145714912, 32'sd0.07756779724624298, 32'sd0.08070048423896917, 32'sd0.0517154540262457, 32'sd1.389418829046508e-120, 32'sd-1.5594661505162914e-116, 32'sd-4.346709676522964e-126, 32'sd-1.0785380977165803e-121, 32'sd-0.016455301893848095, 32'sd0.04186907753120919, 32'sd0.005954559313090512, 32'sd0.051328081051214954, 32'sd-0.016018614854408166, 32'sd0.034441141822543556, 32'sd-0.11105553613728111, 32'sd-0.11579370828499744, 32'sd-0.002553104882315363, 32'sd0.05907954493719257, 32'sd0.014234627453526567, 32'sd-0.0012472348818398172, 32'sd0.09406873431182369, 32'sd0.127725117090855, 32'sd0.08849322412087063, 32'sd-0.09324174109130653, 32'sd0.02373981000822884, 32'sd0.0377917537843893, 32'sd-0.0005767386176377713, 32'sd0.03916718900656955, 32'sd-0.04677778961950388, 32'sd0.030162687690386568, 32'sd-0.14812271543581093, 32'sd0.0409183075698658, 32'sd0.0025988343210962407, 32'sd3.207836283709616e-116, 32'sd2.7625816611553117e-121, 32'sd-0.001815638329503769, 32'sd0.008651598561892498, 32'sd0.0004236308977848514, 32'sd0.03979499077467887, 32'sd0.04509503926793073, 32'sd0.025709404084448953, 32'sd-0.011287488898746098, 32'sd-0.06272991673827247, 32'sd-0.03754788581505553, 32'sd-0.09045923542889699, 32'sd0.07075199112659471, 32'sd0.03403922184989424, 32'sd0.12061598360148364, 32'sd0.03378588986766792, 32'sd0.04075307823815166, 32'sd-0.007260978339998969, 32'sd-0.04011844241826603, 32'sd-0.0055626180621791855, 32'sd0.07142991131024694, 32'sd0.08379231892197758, 32'sd0.01901397001183099, 32'sd-0.06764022373241786, 32'sd-0.15589931418273437, 32'sd-0.14208055021988023, 32'sd-0.08111538908748175, 32'sd-0.04675877135467265, 32'sd0.08078362113723439, 32'sd2.5769778228667016e-114, 32'sd-0.0004892955890161547, 32'sd0.039988777370627754, 32'sd0.04829255609629693, 32'sd-0.047126102506935295, 32'sd0.03154537994216913, 32'sd-0.04616209887462148, 32'sd-0.09245390313211303, 32'sd-0.07794717935374718, 32'sd-0.14531028074808258, 32'sd-0.1843634771116766, 32'sd-0.04657086106273916, 32'sd-0.05018653759869345, 32'sd0.01647049530494371, 32'sd0.06905051862757669, 32'sd0.11790148789000778, 32'sd0.020556319118319545, 32'sd0.10884473833152955, 32'sd0.06584934125222672, 32'sd0.10133746977352062, 32'sd0.014092716664570888, 32'sd-0.10036791708105376, 32'sd-0.06019930289758816, 32'sd-0.1688287028218149, 32'sd-0.07828039518458836, 32'sd0.07918600399877357, 32'sd0.09052343308831629, 32'sd0.03560768120178167, 32'sd-1.3686196611666729e-123, 32'sd0.05005888616294534, 32'sd0.07640765998528182, 32'sd-0.03958442710342827, 32'sd0.06715968461385931, 32'sd-0.03333418631887485, 32'sd0.002994520979057826, 32'sd-0.11907651359054265, 32'sd-0.10848876497556742, 32'sd-0.1306919373086775, 32'sd-0.12378477230195285, 32'sd-0.19422568666539822, 32'sd-0.18634536145982328, 32'sd0.028969951651146016, 32'sd0.02310842833978169, 32'sd0.22071630470781448, 32'sd0.1531999143860794, 32'sd-0.0009346929257984112, 32'sd-0.024301724567485788, 32'sd-0.14475850136506654, 32'sd-0.13512258811410777, 32'sd-0.04767543001088601, 32'sd-0.052531206654108174, 32'sd0.01962852217303643, 32'sd-0.00015298178721263533, 32'sd-0.04882181883637574, 32'sd0.008971565830440424, 32'sd0.08968608714234866, 32'sd0.043058282292348024, 32'sd0.019152866215973334, 32'sd0.012079488187854967, 32'sd0.12269324235261936, 32'sd0.09635144899765019, 32'sd-0.053604109559427286, 32'sd-0.1287654890747886, 32'sd-0.08467661541562883, 32'sd-0.13436906307453056, 32'sd-0.2081179794118449, 32'sd-0.1522721923401614, 32'sd-0.11575490850668452, 32'sd-0.10203107172424258, 32'sd-0.06822297257966131, 32'sd0.17006818323160433, 32'sd0.11988075451958091, 32'sd0.007749964968142289, 32'sd-0.10995565185941371, 32'sd-0.00563850683140977, 32'sd-0.08196902525639939, 32'sd-0.041468873498173464, 32'sd0.07176564254115603, 32'sd-0.04594952107413125, 32'sd0.03735081330616807, 32'sd0.013528540469993293, 32'sd-0.011835557809685038, 32'sd-0.046353792266594335, 32'sd0.009875690235238451, 32'sd0.06425528619872894, 32'sd-0.027977008831658202, 32'sd0.06817074256487639, 32'sd-0.04323742780682021, 32'sd-0.01166452474299802, 32'sd0.03842877191954863, 32'sd-0.0695969005913298, 32'sd-0.12218925239523175, 32'sd-0.18209252067388432, 32'sd-0.13062007038768184, 32'sd-0.10196313035871385, 32'sd-0.05353809965846214, 32'sd-0.06094074589290978, 32'sd0.1325891828947048, 32'sd0.2228398507574266, 32'sd0.09795462745005167, 32'sd0.032568561773287555, 32'sd-0.22249568169446676, 32'sd-0.1255210695956047, 32'sd0.07738283363836237, 32'sd-0.02099723820712561, 32'sd0.018365350365532683, 32'sd-0.042603118908687086, 32'sd-0.0036153719148159444, 32'sd0.05463567829771117, 32'sd-0.08235007727233558, 32'sd0.004522578722344431, 32'sd0.009789394203538337, 32'sd0.02388879656227988, 32'sd0.036569082035221356, 32'sd0.024803035298900017, 32'sd0.00930556241548684, 32'sd-0.037874355306937765, 32'sd-0.061178940258543445, 32'sd-0.09527844020175819, 32'sd-0.1200333239932023, 32'sd-0.1848078555166581, 32'sd-0.07563856755943585, 32'sd-0.027935364338428314, 32'sd-0.0027816637602548, 32'sd0.02110983235798242, 32'sd0.1206269278539527, 32'sd0.17121704250421632, 32'sd-0.005630474761484413, 32'sd-0.23022279811483573, 32'sd-0.2703217116732523, 32'sd-0.02706017918223714, 32'sd0.01168418838715755, 32'sd0.04694139810737114, 32'sd-0.029296062912029106, 32'sd-0.11639617109301093, 32'sd0.10777357214513889, 32'sd-0.0417652208676982, 32'sd-0.12991919463661586, 32'sd0.03465848749255426, 32'sd-0.009063892319266884, 32'sd0.01900361663964919, 32'sd-0.0096959937911439, 32'sd-0.021996638148027957, 32'sd0.13511119440031497, 32'sd-0.062237480638314004, 32'sd0.07614430457401682, 32'sd-0.04303669086763793, 32'sd-0.08656766724097699, 32'sd-0.16886187596792496, 32'sd-0.05939117740858174, 32'sd0.04335038405663328, 32'sd0.022700151826250552, 32'sd0.09496239949125805, 32'sd0.17071453641466655, 32'sd0.10392196129946629, 32'sd-0.1643116798393144, 32'sd-0.2329063179360268, 32'sd-0.06960344147964068, 32'sd0.039419556952157465, 32'sd0.07810151459211559, 32'sd-0.0017484573643295894, 32'sd-0.06789562039002424, 32'sd-0.05782529953676936, 32'sd-0.01720211465217294, 32'sd0.0030261181166682367, 32'sd-0.010071291271732665, 32'sd-0.06723184991558513, 32'sd-0.03682937246405471, 32'sd-0.04644939552645401, 32'sd0.08406126175659971, 32'sd-0.11017665425314623, 32'sd-0.041364375152022, 32'sd0.006344490145583589, 32'sd-0.025936276050346426, 32'sd-0.007978230415792063, 32'sd-0.15663700143425893, 32'sd-0.13122538834782774, 32'sd0.07373535907997014, 32'sd0.08035146559613375, 32'sd0.05799535973794269, 32'sd0.03627199615092221, 32'sd0.0838881084652846, 32'sd-0.062238481459647506, 32'sd-0.10214221884261551, 32'sd-0.021049153162729387, 32'sd0.10564264221138976, 32'sd0.02042450058050596, 32'sd0.0449420237413849, 32'sd0.03350797637649806, 32'sd0.025108664249458897, 32'sd-0.021324799319343248, 32'sd-0.04632260914241599, 32'sd-0.10544031820486409, 32'sd0.034424597418108244, 32'sd-0.12930295431870803, 32'sd0.007423406882814042, 32'sd0.0866669389703205, 32'sd0.02321648328312303, 32'sd-0.08375536332044499, 32'sd-0.06102285130201622, 32'sd-0.019215634285157226, 32'sd-0.04657721687114082, 32'sd-0.0062364779620103445, 32'sd-0.09846409926877701, 32'sd-0.1627587912933219, 32'sd0.049215109821939766, 32'sd0.03207413589707948, 32'sd-0.04178778580775291, 32'sd0.03254039443365291, 32'sd0.04257680531004794, 32'sd0.03093145942058034, 32'sd-0.047170774417380296, 32'sd-0.02537647331211729, 32'sd-0.07287275269211628, 32'sd0.06206313362267792, 32'sd0.01975567308247677, 32'sd-0.0550320173068443, 32'sd-0.01228595892883887, 32'sd0.07957045319471948, 32'sd-0.044139472915679955, 32'sd-0.035701377187270025, 32'sd-0.058244186763400166, 32'sd-0.010769192125100371, 32'sd0.008723428276125605, 32'sd0.017705231236011424, 32'sd-0.031856502818118033, 32'sd-0.11508888419487348, 32'sd-0.109898040662492, 32'sd0.11794370259533826, 32'sd-0.025413831136210374, 32'sd-0.10022872527725304, 32'sd0.01676338754583918, 32'sd-0.045080686280849526, 32'sd0.058198347473351786, 32'sd0.006705158013692499, 32'sd-0.1698875363734729, 32'sd-0.05748330663049239, 32'sd-0.07185164774296542, 32'sd-0.061561939727369556, 32'sd-0.12785020166057914, 32'sd0.032463720999455416, 32'sd0.01713715426757979, 32'sd0.041283859521970064, 32'sd0.14883307179281158, 32'sd0.04076688126258905, 32'sd0.10790008958653395, 32'sd0.07760396150166818, 32'sd0.013849527730773591, 32'sd-0.05527411544073588, 32'sd0.022224943949655546, 32'sd0.015087559593342724, 32'sd0.006512837801747875, 32'sd0.0044110350040555005, 32'sd0.037790064035298956, 32'sd-0.06584357571691829, 32'sd-0.06062534629717784, 32'sd0.10276039888498144, 32'sd-0.03754761298761566, 32'sd0.02726116084111254, 32'sd0.01623641393222944, 32'sd0.05930382101074763, 32'sd0.10132603355106755, 32'sd0.09891282955015744, 32'sd0.005365504211302107, 32'sd-0.05894538517366518, 32'sd-0.1587568059186168, 32'sd0.035190899419123275, 32'sd-0.09087111301333436, 32'sd-0.006385008177583957, 32'sd-0.07716918218149225, 32'sd0.03408585973556401, 32'sd-0.03017476086794521, 32'sd0.0418462983054741, 32'sd0.13827491281214027, 32'sd0.1613327209808044, 32'sd0.09098394643301737, 32'sd-0.013932085649511025, 32'sd-0.03881541627857439, 32'sd-0.008527164872470776, 32'sd-0.06619082492013702, 32'sd0.0330487080643637, 32'sd0.04776331732115372, 32'sd-0.07143773633589037, 32'sd0.00584362739392664, 32'sd0.058679375115497874, 32'sd-0.05993755638250487, 32'sd0.05516785196710357, 32'sd-0.08394197440950776, 32'sd-0.05694540697007706, 32'sd-0.04749641943697514, 32'sd-0.02311312151727315, 32'sd-0.05698796344571337, 32'sd-0.007918971506702689, 32'sd-0.09144932397571606, 32'sd-0.09204646662557399, 32'sd-0.11718781050874615, 32'sd-0.09158413271968571, 32'sd0.027904854504177203, 32'sd-0.037303475397568286, 32'sd0.029482160077960486, 32'sd0.12476959407512105, 32'sd0.039655404729880314, 32'sd0.07579118180641431, 32'sd0.1586205893269527, 32'sd0.0803354246226998, 32'sd0.03410406477439406, 32'sd-0.0004661449751592383, 32'sd-0.03421778740973365, 32'sd0.035409126618744284, 32'sd-0.05122558169765512, 32'sd0.028922991790290346, 32'sd-0.148551500377098, 32'sd0.08170967897444921, 32'sd-0.04688183802284608, 32'sd0.027711748881577934, 32'sd0.1285563453990296, 32'sd-0.05359139535321231, 32'sd0.043652584664916526, 32'sd-0.05961511927780035, 32'sd0.11854866413501437, 32'sd0.029207860315574034, 32'sd-0.035556144822760094, 32'sd0.164709233036127, 32'sd0.020141107670369703, 32'sd0.006287898724819511, 32'sd0.02278855558145908, 32'sd0.11168128442143123, 32'sd0.028666532408595912, 32'sd0.0635249786675842, 32'sd-0.03697005437544252, 32'sd0.03897362960637519, 32'sd0.009905772647509565, 32'sd-3.618899418508825e-05, 32'sd0.077298477138877, 32'sd0.027236060267929924, 32'sd0.06477492863515995, 32'sd3.889812385870669e-129, 32'sd0.006878161808030853, 32'sd-0.03369561277143912, 32'sd-0.0815523108211662, 32'sd-0.001551131745364938, 32'sd0.05193422946422151, 32'sd-0.02887768151029492, 32'sd-0.04980050791119018, 32'sd0.08051841649448731, 32'sd0.056578514189815236, 32'sd0.08306913628856605, 32'sd0.2149801907766217, 32'sd0.16529553636127722, 32'sd-0.0049633884307846285, 32'sd0.13888168003154455, 32'sd0.10091040702039342, 32'sd0.12210864125976781, 32'sd0.11154062394451096, 32'sd-0.004366244368315151, 32'sd0.04808965634483597, 32'sd-0.007141805858720645, 32'sd0.02341566157505759, 32'sd0.011166796976413852, 32'sd0.08097340729939584, 32'sd0.024387466495159597, 32'sd-0.019622290437810466, 32'sd0.007245834450769948, 32'sd0.030549764928492727, 32'sd0.06378842902436697, 32'sd0.04797911317326482, 32'sd-0.05169578582931918, 32'sd-0.08670871802434975, 32'sd0.1039177680686844, 32'sd-0.056091918879020056, 32'sd-0.08132243256543747, 32'sd-0.065475264118447, 32'sd0.014651213979329992, 32'sd0.17703365880406188, 32'sd0.10106212710175398, 32'sd0.1324812639506444, 32'sd0.013469816334351785, 32'sd0.026478917420853187, 32'sd-0.008930899752488883, 32'sd0.07719783616354625, 32'sd0.005975228618178515, 32'sd-0.02308836002077531, 32'sd0.07570874723344402, 32'sd-0.006033734588595852, 32'sd-0.12256585201460357, 32'sd0.017303154443423754, 32'sd0.02332728026423949, 32'sd0.12856860758962835, 32'sd0.05316875977716494, 32'sd-0.024837058632104454, 32'sd0.048177141876800014, 32'sd0.053135172494050954, 32'sd0.05972544998367891, 32'sd0.04572872883262772, 32'sd-0.09152316329061878, 32'sd0.0798927194318595, 32'sd0.046822017518967717, 32'sd0.0745702314684434, 32'sd-0.07650190312610324, 32'sd-0.12049717898513024, 32'sd-0.030566784646738836, 32'sd0.10552104926748414, 32'sd0.050628245917400644, 32'sd0.10634049039005687, 32'sd-0.0596632503431086, 32'sd-0.054536043230791025, 32'sd0.011315995403906763, 32'sd0.09954967690386729, 32'sd0.018569979294632017, 32'sd-0.09735648927381756, 32'sd0.06569118712260995, 32'sd0.11397652788042162, 32'sd0.08728884005971488, 32'sd-0.03022628403122576, 32'sd0.03610002676573502, 32'sd0.08113574101218489, 32'sd0.03418848826174606, 32'sd-0.01693415129403417, 32'sd-0.0329604354202811, 32'sd0.04833303189542708, 32'sd-1.963394424289753e-117, 32'sd0.06946438499585887, 32'sd-0.09133710440906007, 32'sd-0.038640209023862594, 32'sd0.0011278396269938586, 32'sd0.005028138950839504, 32'sd0.016776927423469166, 32'sd0.03506980044628214, 32'sd-0.10645317077503097, 32'sd0.03839312183065678, 32'sd0.009401651072341723, 32'sd0.012897840764689224, 32'sd-0.07772564624850734, 32'sd0.042888888818199175, 32'sd0.0825686649346649, 32'sd-0.03169601585367404, 32'sd-0.02707795770742084, 32'sd-0.07876992366873327, 32'sd-0.14164285154839176, 32'sd0.06706538391701829, 32'sd0.0699303566095548, 32'sd0.024945972004975336, 32'sd0.007777637766399147, 32'sd0.00314601584659166, 32'sd-0.03204395146846318, 32'sd0.009481651837945776, 32'sd-0.12868565881597663, 32'sd-0.013697604031182713, 32'sd-0.006556481117553507, 32'sd-0.031344621577429295, 32'sd-0.1157855815088409, 32'sd0.07473837442730191, 32'sd0.128215416612385, 32'sd-0.033291932402026735, 32'sd0.012125630390552417, 32'sd0.10043268007860874, 32'sd-0.03251430439083625, 32'sd-0.05310330382873493, 32'sd-0.026186487458663296, 32'sd-0.00546498775192757, 32'sd0.11061967079865477, 32'sd0.016510996161483212, 32'sd0.1220016328525297, 32'sd0.08922295081147882, 32'sd-0.04116608195467917, 32'sd0.05615687412583307, 32'sd0.06499891689033598, 32'sd-0.07855294916384971, 32'sd0.007217480498364087, 32'sd-0.006226502752511544, 32'sd-0.04088360747498924, 32'sd0.03020552938494363, 32'sd-0.09796879437633609, 32'sd0.022068176344704437, 32'sd0.025346254612245503, 32'sd0.00851570488307825, 32'sd0.03591717504768037, 32'sd-0.0026699880702050114, 32'sd0.08748559017345164, 32'sd0.05609108213415042, 32'sd0.07372425167608276, 32'sd0.07709356720488676, 32'sd0.07039153703480042, 32'sd0.06809068895737337, 32'sd-0.04762640221924475, 32'sd-0.017944811855938263, 32'sd0.05620791184628719, 32'sd-0.1459011657884974, 32'sd0.1615274234314988, 32'sd0.025282948282170915, 32'sd-0.021691276670424444, 32'sd0.11606585527124408, 32'sd0.10302080891431803, 32'sd0.06123088629695687, 32'sd-0.02498553423708557, 32'sd0.0021285862861189554, 32'sd0.0336537159495954, 32'sd0.002426284041356712, 32'sd-0.07821142656980334, 32'sd-0.017255622302918393, 32'sd-0.06563031486702323, 32'sd0.0015874489254682118, 32'sd0.0066418963685629705, 32'sd0.05543388861255793, 32'sd1.3195566719858613e-118, 32'sd0.075095915322288, 32'sd-0.027009811758741065, 32'sd0.049889163314932816, 32'sd-0.0734889514841639, 32'sd-0.016908468126620356, 32'sd0.03718439776766913, 32'sd0.08685387581206143, 32'sd0.129225028831344, 32'sd0.10157206043575982, 32'sd0.00535046354749796, 32'sd-0.028488508565551865, 32'sd-0.07866386204264801, 32'sd-0.04828408316529936, 32'sd0.047335804971864404, 32'sd0.108788427851898, 32'sd0.021890198087513985, 32'sd-0.09137996402652931, 32'sd-0.04313385921360991, 32'sd0.06959185492818605, 32'sd-0.023704376703296597, 32'sd0.03259968240502566, 32'sd-0.03198846906763768, 32'sd-0.033342027556389195, 32'sd0.018051962377335407, 32'sd-0.04038033848634857, 32'sd0.007107949575064048, 32'sd1.194872584350887e-123, 32'sd-5.635644107906408e-125, 32'sd2.4984539840581506e-126, 32'sd-0.025242168771885818, 32'sd-0.017440672554723074, 32'sd-0.016908024319224686, 32'sd0.0008368354251595632, 32'sd0.033896984618174426, 32'sd0.15819586193478352, 32'sd0.1001561028273267, 32'sd0.020720067477709866, 32'sd-0.11352081274508614, 32'sd0.0042811243775866085, 32'sd0.09579234126217613, 32'sd-0.029035776599971842, 32'sd-0.06997577643851821, 32'sd0.13834498836411713, 32'sd0.046802311420923316, 32'sd0.024698523784023044, 32'sd-0.05207565911222931, 32'sd-0.07491467314459958, 32'sd-0.028200404222874165, 32'sd0.044358752677012614, 32'sd0.06298471899607948, 32'sd0.0505221273772534, 32'sd0.05100491523326313, 32'sd0.07708988100002248, 32'sd0.07973959016612267, 32'sd-4.4331563910251885e-118, 32'sd-4.696706468205164e-127, 32'sd3.1644496493038755e-115, 32'sd0.10402179649589834, 32'sd0.04420640119398252, 32'sd0.03219901784566784, 32'sd0.03791006017792756, 32'sd-0.001576755293799964, 32'sd-0.01603540332261353, 32'sd0.08375051926102482, 32'sd-0.06433644851178688, 32'sd-0.007353694534206793, 32'sd0.09019673793934936, 32'sd0.028332249451856494, 32'sd0.03840327304026143, 32'sd-0.037181619167455465, 32'sd-0.07616219690608157, 32'sd0.05863754684624827, 32'sd0.0007351597065911739, 32'sd-0.04421408372818832, 32'sd0.08205532093904272, 32'sd-0.05739643828124938, 32'sd-0.008020925717971873, 32'sd0.016355789146763704, 32'sd0.057129396749361204, 32'sd0.03384632132231464, 32'sd0.024842439269894313, 32'sd-0.012195486511181719, 32'sd-4.9152734514931627e-116, 32'sd-1.3794622353881658e-121, 32'sd6.24914919344933e-125, 32'sd-4.281133248864022e-115, 32'sd0.027538370193028294, 32'sd0.06193066368376364, 32'sd0.0320078126882235, 32'sd0.08220426655637136, 32'sd0.053490829359545716, 32'sd0.020733254666800524, 32'sd-0.09659185131679794, 32'sd-0.08881820207048399, 32'sd-0.01587812350917088, 32'sd-0.0552224359321833, 32'sd-0.13387061447611007, 32'sd0.005386784176523064, 32'sd-0.1459881461691854, 32'sd-0.17461793337402615, 32'sd-0.0619059439555427, 32'sd0.10965495417164342, 32'sd0.10125375479171356, 32'sd0.003986342884352869, 32'sd0.01698099297872669, 32'sd0.025100274326575286, 32'sd-0.011828339238994744, 32'sd0.08492174965910762, 32'sd0.017560659635227207, 32'sd3.248920628018137e-120, 32'sd-8.63795388720739e-122, 32'sd1.292803697527093e-122, 32'sd3.540455722343929e-126, 32'sd-7.723547093369051e-122, 32'sd-1.046281500803773e-119, 32'sd0.08087538797709318, 32'sd0.033360595865772835, 32'sd0.041323164928239176, 32'sd0.03394101165905414, 32'sd0.009539938524740037, 32'sd0.03490716986688725, 32'sd-0.015560066061219052, 32'sd-0.04632493422159953, 32'sd-0.05201096541658119, 32'sd0.06540499108557064, 32'sd-0.004409049556425292, 32'sd0.08272608948414072, 32'sd-0.05613996871886213, 32'sd0.0329591371390863, 32'sd0.09272182932300628, 32'sd0.1209359849660012, 32'sd0.06200316434990409, 32'sd0.016158468042001738, 32'sd0.0595709711489536, 32'sd0.05880783544765369, 32'sd-1.0847567576757552e-119, 32'sd-1.1097216532046988e-122, 32'sd8.53252702333064e-117, 32'sd1.0461560824930438e-117},
        '{32'sd-1.892337908434894e-125, 32'sd-8.177167145744672e-117, 32'sd-4.481940099458558e-118, 32'sd4.772893998939898e-123, 32'sd-1.0088191361111416e-120, 32'sd-4.1031748244385835e-117, 32'sd-1.1266858798208275e-122, 32'sd-2.6169217166004522e-126, 32'sd-4.187897587017713e-126, 32'sd5.548293764588426e-115, 32'sd2.3693336823639324e-116, 32'sd3.768925157953638e-122, 32'sd-0.05804394268281986, 32'sd-0.0930760536212465, 32'sd-0.02592150131772974, 32'sd-0.0077220478967430384, 32'sd8.147253809005459e-126, 32'sd5.2334392872602515e-118, 32'sd4.445570026265794e-125, 32'sd2.132134632525407e-124, 32'sd-2.0015192971099742e-119, 32'sd-9.73011101986536e-118, 32'sd2.555753169906604e-123, 32'sd3.8006243360455776e-123, 32'sd-1.6649213537172185e-121, 32'sd-3.2804533822936064e-116, 32'sd-3.8549978594358324e-123, 32'sd1.4887859157181083e-120, 32'sd-6.656355564678625e-117, 32'sd-1.2398140881141981e-116, 32'sd-7.734822176551829e-120, 32'sd-4.1665593246116005e-118, 32'sd-0.03529643943743521, 32'sd-0.04851732696422242, 32'sd-0.07561063965337932, 32'sd-0.07384431726205742, 32'sd-0.13266505196026354, 32'sd-0.013385070823613003, 32'sd-0.007152050337835748, 32'sd0.01989774505780774, 32'sd0.020246298347451352, 32'sd0.06662565494853445, 32'sd0.028550455404242975, 32'sd-0.03404575734178399, 32'sd0.0021521501840693377, 32'sd-0.0785212863435761, 32'sd-0.0010592042304463705, 32'sd-0.07195160823855377, 32'sd-0.11065895363038414, 32'sd-0.10091158278558929, 32'sd0.006828573678052936, 32'sd0.014223801785938614, 32'sd6.687782523774645e-124, 32'sd1.3105317053918676e-115, 32'sd3.329055981008575e-123, 32'sd-1.4265270478752636e-118, 32'sd-1.7336162863924968e-125, 32'sd1.0405727571689214e-127, 32'sd-0.04176514339517757, 32'sd0.017693390570676877, 32'sd-0.06662994836478969, 32'sd-0.04184782531340687, 32'sd0.001592609642740658, 32'sd-0.026181883383085428, 32'sd0.034752929882282034, 32'sd0.037952177798969304, 32'sd0.11606433339618889, 32'sd0.02041146694106899, 32'sd0.0559139075947245, 32'sd0.05673441796373222, 32'sd0.05561941993715279, 32'sd-0.09554616518035526, 32'sd-0.08882241516698272, 32'sd0.013683078128961308, 32'sd-0.10759059502641982, 32'sd-0.04974564137264518, 32'sd-0.033934736279822485, 32'sd-0.07706093448261514, 32'sd0.04056765025284111, 32'sd-0.051317736174555754, 32'sd0.0014251512746304236, 32'sd-0.05616874312222837, 32'sd8.760047412539571e-123, 32'sd3.944687313135657e-120, 32'sd3.7762623657080655e-126, 32'sd-1.0244139274483457e-125, 32'sd-0.01180299161848485, 32'sd-0.01094361440163879, 32'sd-0.05377132729259376, 32'sd0.05525337848433231, 32'sd-0.03834849339348447, 32'sd0.0845438270127048, 32'sd-0.00030357747514680593, 32'sd0.028147592935744165, 32'sd0.07845085575547867, 32'sd0.06075486380543604, 32'sd0.05017944292263193, 32'sd0.10189508887412393, 32'sd0.07521176039210503, 32'sd-0.1172961686370545, 32'sd-0.06714277959961064, 32'sd-0.07457401428379515, 32'sd-0.011308097666105733, 32'sd0.0009667878640641393, 32'sd-0.065732282838858, 32'sd-0.06908600093340862, 32'sd-0.002595734046879225, 32'sd-0.012855748564229337, 32'sd0.10712077099135901, 32'sd0.040831177438760365, 32'sd-0.022066510250555952, 32'sd-2.461162875662949e-120, 32'sd-1.039801325034137e-120, 32'sd-0.066239396671067, 32'sd-0.00425756647661376, 32'sd0.009760724186802601, 32'sd-0.045372808102851055, 32'sd-0.04924576823186041, 32'sd0.1321799445577981, 32'sd0.21054056519202008, 32'sd0.1672533189974596, 32'sd-0.05144247817248176, 32'sd0.060525423912591275, 32'sd0.13979077213947064, 32'sd0.10922123712695433, 32'sd0.06033431294505041, 32'sd0.08382454151125682, 32'sd0.033009983366588946, 32'sd0.0006720672678925334, 32'sd-0.06654145299604175, 32'sd0.01766416913133697, 32'sd-0.0035906529871914004, 32'sd-0.009744327656609944, 32'sd-0.03693716035743907, 32'sd0.0476107213444446, 32'sd-0.0017908592380376637, 32'sd0.037428700059946765, 32'sd-0.0722301081307413, 32'sd-0.021267387287639612, 32'sd-0.0878758230033271, 32'sd1.9730483052560883e-121, 32'sd0.050174100936099246, 32'sd0.00937939825903424, 32'sd0.13796148877759112, 32'sd0.08191912502386749, 32'sd-0.00743693172357894, 32'sd-0.05102988006313168, 32'sd-0.008081217595001255, 32'sd-0.04341723004041886, 32'sd0.0011335931639482992, 32'sd0.006664842160407745, 32'sd-0.015577652635427408, 32'sd0.04205885538001862, 32'sd0.15320580488749785, 32'sd0.0758138878716525, 32'sd0.03669657247088101, 32'sd0.13496262654800142, 32'sd0.09639392321271706, 32'sd0.14345661807874877, 32'sd0.12025680586524058, 32'sd-0.08168903926593772, 32'sd-0.047207936728585656, 32'sd-0.09091686778037815, 32'sd-0.07614620470271485, 32'sd-0.03441885041061436, 32'sd0.05638001904939429, 32'sd0.06518409430961718, 32'sd0.01010379414092843, 32'sd1.3692963571029903e-121, 32'sd-0.09130106846483865, 32'sd-0.07908475647420675, 32'sd0.09122963381142651, 32'sd0.09295323760977359, 32'sd-0.004618747670079157, 32'sd-0.1559737552388506, 32'sd-0.14605888016807433, 32'sd-0.08126565594148018, 32'sd-0.15258992710378347, 32'sd0.019645392726018732, 32'sd-0.027443064448280853, 32'sd0.07016631524948962, 32'sd0.05125512264085991, 32'sd0.09518615689271058, 32'sd0.10569709675696222, 32'sd0.20507736232303211, 32'sd-0.036618918133401894, 32'sd0.16169872913219377, 32'sd-0.002550027357158884, 32'sd-0.06847677869465363, 32'sd-0.20583405385302267, 32'sd-0.1729379297828, 32'sd-0.15272177248417895, 32'sd-0.08362390278289707, 32'sd0.06585321211162105, 32'sd-0.06770817581332478, 32'sd-0.010079549420938432, 32'sd-0.014201585912968323, 32'sd0.03596494407491644, 32'sd-0.08261756139605785, 32'sd-0.027825952487855743, 32'sd-0.016945028937559337, 32'sd-0.058777238525804444, 32'sd-0.09759907161696858, 32'sd-0.05061099058942409, 32'sd-0.016588144079638892, 32'sd-0.12070110628782023, 32'sd-0.05667176002271876, 32'sd-0.07335650395551387, 32'sd-0.032947783074721564, 32'sd-0.06069001544592382, 32'sd0.034545053289036814, 32'sd0.14859511872188708, 32'sd0.056258694531695984, 32'sd0.0014120649096016269, 32'sd0.09768457895000177, 32'sd-0.026910951886543185, 32'sd0.029085051373736456, 32'sd-0.08415948519938758, 32'sd-0.04748730218987635, 32'sd-0.046580509782068374, 32'sd-0.11317193175845279, 32'sd-0.012990227964529186, 32'sd-0.11049906036129144, 32'sd0.004941120617818432, 32'sd-0.08910048108745787, 32'sd0.04638545232238718, 32'sd-0.059949420849918264, 32'sd-0.0034939806871576574, 32'sd0.018949551663746525, 32'sd-0.07198583728974856, 32'sd-0.07112198079976847, 32'sd-0.055181684237876734, 32'sd0.04899275280212839, 32'sd-0.08573168466264179, 32'sd-0.04881019962019438, 32'sd-0.14710181333648034, 32'sd-0.1341963821217603, 32'sd-0.11680152257934816, 32'sd-0.0069199374312866975, 32'sd-0.09786630589993525, 32'sd0.01003482199891014, 32'sd0.09207220201722889, 32'sd0.1247542226589189, 32'sd0.05868722798758191, 32'sd-0.03760567944336212, 32'sd-0.1114836480307358, 32'sd-0.06088929299475406, 32'sd-0.07661681287469853, 32'sd-0.09144813248800587, 32'sd-0.13040967601280862, 32'sd-0.019471558584664424, 32'sd-0.10733316922026562, 32'sd-0.10413134551450984, 32'sd-0.05787943272179884, 32'sd-0.049770911880763116, 32'sd0.0652814412570802, 32'sd-0.07482387303884507, 32'sd0.03358225514473597, 32'sd0.014036473361505401, 32'sd0.012422631673675785, 32'sd0.07091110307405027, 32'sd-0.022951512551022037, 32'sd-0.14918765758427097, 32'sd-0.04343258121466118, 32'sd-0.14989678728004366, 32'sd-0.14620728254707088, 32'sd-0.1736210773727516, 32'sd-0.04174827770854562, 32'sd-0.02262733522489511, 32'sd0.07477744834490427, 32'sd0.16781747129562677, 32'sd0.11723833820624631, 32'sd0.08569927373657578, 32'sd-0.0728779375323261, 32'sd-0.11017072582673407, 32'sd-0.11796666877570457, 32'sd-0.1881139798340474, 32'sd-0.07622211683624784, 32'sd-0.017252503703863595, 32'sd0.022969447621999785, 32'sd-0.058303856144540506, 32'sd0.004551637031560149, 32'sd0.04758699365086422, 32'sd-0.0004589533783549484, 32'sd0.044226268062205774, 32'sd0.07079911987933288, 32'sd0.10798239760087841, 32'sd0.046155571056389386, 32'sd-0.007719318365743172, 32'sd-0.09750169380650817, 32'sd-0.11984871025282677, 32'sd-0.20114504529204066, 32'sd-0.11430855185221798, 32'sd-0.08154095712186134, 32'sd0.010971239474893292, 32'sd-0.05899694448054734, 32'sd-0.06014142322636153, 32'sd0.08938286852050113, 32'sd0.10737403465867817, 32'sd0.04266667338613027, 32'sd0.026871429767171114, 32'sd0.07334780952386304, 32'sd-0.06155171933492216, 32'sd-0.04502686656275023, 32'sd-0.10058798419024004, 32'sd0.04317273875030035, 32'sd-0.07508279672059051, 32'sd-0.073501603500061, 32'sd-0.0732034936829663, 32'sd-0.044976409591928904, 32'sd-0.11403532892070532, 32'sd-0.0065576571130335996, 32'sd-0.04717389213618651, 32'sd0.060278195598343756, 32'sd0.0033714766433287874, 32'sd-0.02170106447390511, 32'sd-0.21699922916523368, 32'sd-0.11791888895575492, 32'sd-0.0806054555220777, 32'sd-0.0015170009968473498, 32'sd-0.02253743189837863, 32'sd0.05636171363235037, 32'sd-0.020310832406708754, 32'sd-0.062178092633942285, 32'sd-0.043641132512908, 32'sd0.08352546050916144, 32'sd0.01745450244625121, 32'sd-0.031226704384093154, 32'sd0.00782208461675241, 32'sd-0.03689467865648152, 32'sd-0.08080492363409424, 32'sd-0.07759983552649476, 32'sd-0.16572233395654754, 32'sd0.02084013563107093, 32'sd0.017713536790081814, 32'sd-0.10369363131735222, 32'sd-0.05324130884296856, 32'sd-0.07363359676713362, 32'sd0.005664094682539403, 32'sd-0.1136679097569372, 32'sd0.03503468740192251, 32'sd-0.16804458537453387, 32'sd-0.05043219191845006, 32'sd-0.08962132870130514, 32'sd-0.18382373857110165, 32'sd-0.034225864696149556, 32'sd-0.04120915795269648, 32'sd-0.10305876377771736, 32'sd-0.09422194891167877, 32'sd-0.07706509686068463, 32'sd0.06916388833087306, 32'sd-0.08304913779981343, 32'sd-0.014427883696168878, 32'sd0.05095078557130036, 32'sd-0.18814187430282756, 32'sd0.017180640023150083, 32'sd0.002928973080720795, 32'sd-0.11434450696261177, 32'sd-0.1412821254765251, 32'sd-0.09723689496862797, 32'sd-0.07896209843845682, 32'sd0.04514178613406128, 32'sd-0.1212044897790603, 32'sd-0.08411344362783693, 32'sd-0.0349166403693689, 32'sd-0.021838565986274146, 32'sd-0.04850864829660653, 32'sd0.05153466618804955, 32'sd-0.06499783490087091, 32'sd-0.09163661674116508, 32'sd-0.13775675478644592, 32'sd-0.02414057094494983, 32'sd0.09647900683190133, 32'sd0.05323813773954671, 32'sd-0.12207065820676431, 32'sd-0.14199568839290522, 32'sd-0.0984068788665877, 32'sd-0.0939219409335898, 32'sd0.10148248152009996, 32'sd-0.11731841235058589, 32'sd-0.037396788188256334, 32'sd0.06690533260081297, 32'sd-0.0628309924674042, 32'sd0.13268617441411198, 32'sd0.10403685458124017, 32'sd-0.04587503193828363, 32'sd-0.062110687990673014, 32'sd-0.05066653286870991, 32'sd-0.0034958464205015133, 32'sd0.09905212224584903, 32'sd-0.040529893871258584, 32'sd-0.030682954669902725, 32'sd-0.07364692741456776, 32'sd-0.10537998644242304, 32'sd-0.09418100107052832, 32'sd-0.004678641373834197, 32'sd0.04123227206491657, 32'sd-0.08777888102806063, 32'sd-0.09332253412839199, 32'sd-0.05006879542824863, 32'sd-0.03976380738374522, 32'sd-0.0660003528895798, 32'sd-0.09488596141128458, 32'sd-0.10940163346067591, 32'sd-0.09208825269327982, 32'sd-0.044124983007555935, 32'sd0.10332804416050058, 32'sd-0.07738047703136217, 32'sd-0.04343879383013798, 32'sd-0.0454117227413044, 32'sd0.03182391195243958, 32'sd0.009226354324898088, 32'sd0.041646641063371764, 32'sd-0.058956957958677385, 32'sd-0.09562290954531748, 32'sd-0.08256872440742993, 32'sd-0.12567790565854242, 32'sd0.04154988999282393, 32'sd0.0739802555381146, 32'sd0.003656833118307358, 32'sd-0.012934955398804154, 32'sd-0.005981162697289002, 32'sd-0.023641351186034328, 32'sd0.1200366934302881, 32'sd-0.05442191096474799, 32'sd0.021352657224036037, 32'sd-0.0674546059345351, 32'sd-0.07121042435872672, 32'sd-0.11554521109306716, 32'sd0.03172688313384092, 32'sd-0.0923994623500308, 32'sd0.010887829555489236, 32'sd-0.03827314492216792, 32'sd0.07663420535829892, 32'sd0.1333677930378003, 32'sd-0.030669687387954826, 32'sd0.04886812411010244, 32'sd-0.02814466371241687, 32'sd0.045385202980163006, 32'sd-0.10855636548767772, 32'sd-0.09825927365778472, 32'sd0.003478053290203916, 32'sd0.10392231889631162, 32'sd0.08540675295496832, 32'sd-0.0022133677360035484, 32'sd0.02909285200701758, 32'sd-0.013325998771871076, 32'sd0.029855197441832536, 32'sd-0.05142278550242606, 32'sd-0.08168498606696063, 32'sd-0.1718539610845101, 32'sd0.0033154198957574925, 32'sd-0.010180604743525395, 32'sd-0.09518211440321067, 32'sd-0.04681427307937961, 32'sd-0.13921605941219978, 32'sd-0.02903248161553306, 32'sd-0.04213339281675553, 32'sd-0.057052565307030234, 32'sd-0.1039068684760888, 32'sd0.02301203610472465, 32'sd0.04261557405702679, 32'sd-0.04422822405976921, 32'sd-0.1342703926138197, 32'sd-0.08446343909073453, 32'sd0.020862120436108997, 32'sd-0.007454046919285511, 32'sd0.035837212426263705, 32'sd-0.05124858201248867, 32'sd-0.00549193834193349, 32'sd0.03839160484710731, 32'sd0.007828725423262664, 32'sd-0.0032421328445593573, 32'sd0.01784457481572981, 32'sd-0.0020097965270661935, 32'sd-0.104818454726347, 32'sd6.702566278197424e-115, 32'sd-0.1089082502107888, 32'sd-0.13607068840557526, 32'sd-0.00019881074725848954, 32'sd-0.03592030770671053, 32'sd-0.013452009179167546, 32'sd-0.03278702155211084, 32'sd0.011467179900861818, 32'sd-0.02679661745501517, 32'sd-0.07251182761753314, 32'sd-0.021869343031622194, 32'sd-0.02698601777408933, 32'sd-0.06503181710110724, 32'sd-0.0740241591142442, 32'sd-0.09721737989023467, 32'sd-0.01174011206567049, 32'sd0.029630806431408408, 32'sd-0.012685781291285928, 32'sd-0.007882434070257517, 32'sd0.020286224057015852, 32'sd-0.12087869720909823, 32'sd-0.002567382001415922, 32'sd0.03703020563272661, 32'sd-0.062368942792398054, 32'sd0.10128273613964574, 32'sd0.09201097757820173, 32'sd-0.05727180794307687, 32'sd-0.09528134327132762, 32'sd-0.036873989692166244, 32'sd-0.0734133706620223, 32'sd-0.0575654647247643, 32'sd-0.003408446599179281, 32'sd0.05664237162758035, 32'sd-0.033809008942304174, 32'sd0.023087645229642205, 32'sd-0.14222552125992746, 32'sd0.06119209297001074, 32'sd0.08832977514939865, 32'sd0.08749477060139757, 32'sd-0.030256405237791988, 32'sd-0.1508096823598619, 32'sd-0.06995988413080666, 32'sd-0.062452653536412564, 32'sd0.02671157881164144, 32'sd0.04467973509200006, 32'sd0.04559684843382094, 32'sd0.0514283248485109, 32'sd-0.037293980723669545, 32'sd0.01131174512034714, 32'sd-0.028128681579238608, 32'sd-0.08281205632843776, 32'sd-0.02193678504790565, 32'sd0.025634992871380324, 32'sd0.07394664653374029, 32'sd-0.018270602882337634, 32'sd-0.09200845687549156, 32'sd-0.030300322759860013, 32'sd-0.04827719988754153, 32'sd-0.05645566379165686, 32'sd-0.0009211793949846597, 32'sd-0.045590232007277735, 32'sd-0.02272994113989495, 32'sd-0.04245448306402882, 32'sd-0.010604230941713987, 32'sd-0.09437911334929146, 32'sd0.08713949298963226, 32'sd0.04058301371419648, 32'sd-0.10048071817379294, 32'sd-0.07575820129984055, 32'sd-0.01794873551821668, 32'sd-0.034353067446445305, 32'sd0.08795671837600381, 32'sd0.10353387925338967, 32'sd0.09978430328472768, 32'sd0.05177694776627975, 32'sd0.009646413481118358, 32'sd-0.07885252055162531, 32'sd-0.006198576340678217, 32'sd-0.060622056422271406, 32'sd-0.08855139311348076, 32'sd-0.06277753706752698, 32'sd-0.08767729954854528, 32'sd0.0713859735921764, 32'sd-0.031460050933916975, 32'sd8.108057663925457e-117, 32'sd0.022177242612748026, 32'sd-0.023181653461470626, 32'sd0.06621325980396407, 32'sd-0.06233523550341152, 32'sd0.009800267353368235, 32'sd-0.02339260120839273, 32'sd-0.03027620556012319, 32'sd0.005808237945192975, 32'sd0.11263829996904083, 32'sd0.06077654328948835, 32'sd0.029816471456539484, 32'sd0.033288394208671516, 32'sd0.07835332763563553, 32'sd0.053270149168150684, 32'sd0.11935123304435585, 32'sd0.08438167898260458, 32'sd-0.0023912246723898243, 32'sd0.10224139046931784, 32'sd-0.025941913485571774, 32'sd0.024609585608771068, 32'sd-0.0857665357063225, 32'sd-0.0826365716856505, 32'sd-0.014045789511890781, 32'sd-0.04488828124552077, 32'sd-0.05225664778092067, 32'sd-0.061760345706308416, 32'sd-0.07785068856550788, 32'sd-0.024497362816446967, 32'sd0.09398896317792789, 32'sd-0.0006184922752838251, 32'sd0.07231341047555534, 32'sd0.020189182528736707, 32'sd-0.08661318315978998, 32'sd-0.04656273214566429, 32'sd0.08504999350741618, 32'sd-0.03565217055764543, 32'sd0.005802518951538786, 32'sd0.10887927104350288, 32'sd0.010755043398589799, 32'sd0.06254419421962358, 32'sd0.20564576172386506, 32'sd0.14365478357075445, 32'sd0.023527212134629806, 32'sd-0.005481046030413605, 32'sd0.024085517058295095, 32'sd0.024686176254662136, 32'sd0.06837387622925314, 32'sd-0.06721200298915947, 32'sd-0.07311191058474478, 32'sd-0.019725724924019826, 32'sd0.0010812664286876962, 32'sd0.019112891579314357, 32'sd0.0011361884812072388, 32'sd0.017950921358690707, 32'sd-0.02353958615439917, 32'sd-0.03919253365053385, 32'sd0.03120393596875522, 32'sd-0.041936643658186036, 32'sd-0.12030800787641782, 32'sd0.010785040283535146, 32'sd-0.02662907528949772, 32'sd-0.10445121151358648, 32'sd-0.08789085363037992, 32'sd-0.030615371865676408, 32'sd0.07897550957434647, 32'sd-0.03601889623526616, 32'sd0.09827765738377213, 32'sd0.03615563293461879, 32'sd0.12856038028289862, 32'sd0.05079386620108339, 32'sd0.11732704084843244, 32'sd0.022100873239834323, 32'sd0.021347749953061573, 32'sd-0.0919053733146775, 32'sd0.09428912941407881, 32'sd0.03412182571024911, 32'sd0.10461570131595548, 32'sd0.009874707336255562, 32'sd0.04768565450480322, 32'sd0.08848482842169829, 32'sd0.011474436614719304, 32'sd-0.037208355887499746, 32'sd-0.040973041000871256, 32'sd-1.0420848859677345e-120, 32'sd0.0037077538790715524, 32'sd0.00509690223223497, 32'sd-0.0075094929755139955, 32'sd-0.07397177818634362, 32'sd0.06887152764866433, 32'sd-0.09252643892607304, 32'sd0.030929400619320088, 32'sd0.10794656430352155, 32'sd0.08117310591592627, 32'sd0.024768500427564774, 32'sd0.19037854459168732, 32'sd0.011072147750987284, 32'sd0.0740518143310374, 32'sd-0.018325165639987245, 32'sd0.15494712168757305, 32'sd0.11109308260342453, 32'sd0.0030121782131881975, 32'sd0.01730051034083242, 32'sd-0.09933984699601925, 32'sd0.10714049637806894, 32'sd0.025728124866235345, 32'sd0.032274977797079364, 32'sd-0.016615576458999193, 32'sd-0.01958924270820494, 32'sd0.04371192325454519, 32'sd-0.12138450247147403, 32'sd6.530787946187916e-126, 32'sd1.463717571667711e-115, 32'sd6.675360669501131e-124, 32'sd0.012101904930543427, 32'sd-0.017417127558877678, 32'sd-0.11224067247777632, 32'sd0.07510137397594684, 32'sd0.07536307050733104, 32'sd0.011656493767248716, 32'sd0.004841138639614748, 32'sd0.1275092552412135, 32'sd0.1673601394310462, 32'sd0.14511605018059923, 32'sd0.12253423558945317, 32'sd0.03876315246946197, 32'sd0.04515624634690169, 32'sd0.06607329119739369, 32'sd0.00520883177663593, 32'sd0.15613893822929895, 32'sd0.010981569325310183, 32'sd-0.00655073172270591, 32'sd0.07263461096604201, 32'sd0.03005589650340662, 32'sd-0.18789629641754182, 32'sd-0.11367475454502492, 32'sd0.044961169913376335, 32'sd0.06310850090619366, 32'sd-0.08266186082232505, 32'sd-1.4014091921551504e-123, 32'sd6.160250953520556e-124, 32'sd-2.7098803522133765e-123, 32'sd0.0658121331181852, 32'sd-0.035624644281939254, 32'sd0.013862717751769733, 32'sd0.0007377828316516065, 32'sd0.13037072631660057, 32'sd0.11471157893226214, 32'sd0.07443881439381894, 32'sd0.02152895265038443, 32'sd0.11343702656055163, 32'sd-0.03584881485117571, 32'sd0.0722729098262469, 32'sd0.06637571000985241, 32'sd0.01166379355160911, 32'sd-0.10716462201914718, 32'sd0.05480226154215524, 32'sd0.008318974008345257, 32'sd0.077565527089166, 32'sd-0.012934189511831722, 32'sd0.03845489612491804, 32'sd0.017471556913006118, 32'sd0.0552577105175345, 32'sd-0.041124284087228374, 32'sd-0.023805509863452406, 32'sd-0.07242989673081593, 32'sd-0.07293349367574752, 32'sd-2.7677394144217025e-121, 32'sd-1.556969132425232e-124, 32'sd-3.277636339175754e-119, 32'sd-2.586412111414413e-129, 32'sd-0.030556246308013527, 32'sd0.03550378047068631, 32'sd0.03207675556351479, 32'sd-0.1275397536520454, 32'sd-0.10927172700985013, 32'sd-0.08848337656290443, 32'sd-0.14972411229259938, 32'sd-0.04545028857636722, 32'sd-0.13770166675030052, 32'sd-0.03812681531800915, 32'sd-0.0692889027372627, 32'sd-0.16940666839428065, 32'sd-0.1218134928849916, 32'sd-0.06314895004185397, 32'sd-0.03919397410163912, 32'sd-0.03784667200195428, 32'sd-0.02272681349224467, 32'sd-0.09368407661899869, 32'sd-0.1339713570715115, 32'sd-0.08671465990042476, 32'sd-0.08958296042888189, 32'sd-0.019149935919397672, 32'sd0.0327297172507092, 32'sd3.9652968586858585e-119, 32'sd9.444360147222837e-123, 32'sd-9.540247753309037e-123, 32'sd6.53843814835999e-117, 32'sd-1.0988459426918805e-121, 32'sd1.032337053321939e-119, 32'sd-0.09359714921617535, 32'sd-0.11027269793952527, 32'sd-0.06625315152080377, 32'sd-0.042163567136503204, 32'sd-0.09935857448751884, 32'sd-0.03855303368535041, 32'sd0.017239609138969637, 32'sd0.02550464277278528, 32'sd-0.08532369738252117, 32'sd-0.0928298867969954, 32'sd-0.025960569672579557, 32'sd-0.11403890019119906, 32'sd-0.03968566083476146, 32'sd0.0054390443719446215, 32'sd0.0005281849270416404, 32'sd-0.01762643997056523, 32'sd-0.11210039404247975, 32'sd-0.03183256613046512, 32'sd-0.054731193398373, 32'sd-0.07584489580586415, 32'sd-5.867720260479855e-118, 32'sd-2.6015294125277254e-119, 32'sd6.124698866973333e-122, 32'sd2.382678659387524e-124},
        '{32'sd-2.2146575385222224e-122, 32'sd-1.7603969875503787e-125, 32'sd-4.9124586177581925e-121, 32'sd6.446701762001924e-115, 32'sd-4.209150578273593e-121, 32'sd1.417600965859739e-125, 32'sd1.2580643160451523e-118, 32'sd-1.0474158640678532e-120, 32'sd1.375912355136918e-118, 32'sd5.379345588680573e-118, 32'sd-2.5811342574244265e-117, 32'sd-1.8278110795916528e-126, 32'sd-0.042062640256573025, 32'sd0.00861891510856285, 32'sd-0.025768736279601585, 32'sd-0.0007941659101343513, 32'sd1.1290987403902304e-119, 32'sd-9.991435846632694e-116, 32'sd2.615988517694231e-126, 32'sd-4.930402562121646e-121, 32'sd-8.531442050293155e-120, 32'sd2.115493612682419e-123, 32'sd4.4678745912967674e-123, 32'sd-3.035440676641366e-119, 32'sd1.119101628829941e-123, 32'sd-4.426833143992529e-118, 32'sd-3.404607079171624e-114, 32'sd7.520963579627123e-115, 32'sd-9.227733442957975e-122, 32'sd-5.21988081983911e-118, 32'sd2.4027758042527315e-124, 32'sd4.389392425800094e-123, 32'sd0.02524772040824068, 32'sd-0.01483533197135916, 32'sd0.07427488478018253, 32'sd0.017240309757030513, 32'sd-0.0170878870589047, 32'sd0.02446758832181063, 32'sd-0.013447012066703765, 32'sd0.08070558093887276, 32'sd-0.07233361781563291, 32'sd-0.029118757059447862, 32'sd-0.011539478070496862, 32'sd-0.05004797031210393, 32'sd0.0034851155037951952, 32'sd0.011944790897956513, 32'sd-0.031167790202344614, 32'sd0.061910627852492114, 32'sd0.04188837864453725, 32'sd0.03566814445202052, 32'sd0.003760041918818527, 32'sd0.02704753607012976, 32'sd5.41142018121014e-124, 32'sd2.1048219710820816e-117, 32'sd-4.865212222885017e-123, 32'sd2.3866806638664612e-116, 32'sd3.9234703823380835e-118, 32'sd-6.811126734338398e-126, 32'sd0.02690778942777269, 32'sd-0.016093870651518745, 32'sd0.030106840103957765, 32'sd-0.03616549794490815, 32'sd0.008169794477320323, 32'sd0.025292060868174607, 32'sd-0.07997267765534087, 32'sd0.0054695121130634156, 32'sd0.034459677227683026, 32'sd0.04537928275109039, 32'sd0.01386102316288649, 32'sd0.03473195566477814, 32'sd-0.007205897799739785, 32'sd0.03503537360730678, 32'sd-0.03436531404758907, 32'sd0.052056430116782224, 32'sd0.10652465926568863, 32'sd0.09065158183022225, 32'sd0.10647784643932595, 32'sd0.1173820131622145, 32'sd-0.049985521500734695, 32'sd-0.007932936090167268, 32'sd0.027405634417043172, 32'sd0.13028626704546445, 32'sd-7.475781333528968e-125, 32'sd2.7011824553885115e-123, 32'sd-6.33515778978182e-123, 32'sd-8.226137142823412e-127, 32'sd0.11082049900314503, 32'sd0.02589726105671741, 32'sd0.01565057960635347, 32'sd0.03404393617637624, 32'sd-0.03928341262968946, 32'sd-0.04009295550213328, 32'sd-0.09198697874770301, 32'sd0.04838035742271617, 32'sd0.0433323727321156, 32'sd0.028299684390367574, 32'sd-0.012243675351479437, 32'sd0.047679868223264, 32'sd-0.056465586660233436, 32'sd0.038190724852941074, 32'sd0.03393443572261084, 32'sd-0.09009960821866866, 32'sd-0.013374632126450785, 32'sd0.013130152302941275, 32'sd0.043702892768857846, 32'sd-0.019857824874473698, 32'sd0.09825446684929166, 32'sd0.06345618130796511, 32'sd0.05274408762826266, 32'sd0.04090044145448793, 32'sd0.056750898184524695, 32'sd-2.2011441790574748e-116, 32'sd9.924573937318873e-120, 32'sd0.025428362704673874, 32'sd0.06954351386409807, 32'sd0.03189149478477069, 32'sd-0.06782787400172767, 32'sd0.08418283138002844, 32'sd0.004813589762553832, 32'sd0.00907888875607715, 32'sd-0.05244701847533081, 32'sd-0.1435433105719091, 32'sd-0.00017550411631205612, 32'sd-0.15250518727492152, 32'sd-0.004447117057807022, 32'sd-0.07296992341764834, 32'sd-0.009189061812891364, 32'sd-0.09762207901254198, 32'sd0.04140550539710756, 32'sd0.1148522888628356, 32'sd0.07792777512623247, 32'sd0.053735580754619344, 32'sd0.047627727519011204, 32'sd-0.07209035209683617, 32'sd0.1363393029342935, 32'sd-0.00451966947277244, 32'sd-0.05562672637671937, 32'sd-0.15118900593783896, 32'sd0.010956930505126623, 32'sd0.05441757944949419, 32'sd6.348298687503541e-125, 32'sd0.05860434433285021, 32'sd0.023853091646763053, 32'sd-0.05230912037903534, 32'sd0.042265184432115986, 32'sd-0.0035448224363888547, 32'sd-0.03617121001096223, 32'sd0.059062729103208464, 32'sd-0.022847363177711622, 32'sd-0.08514462058147733, 32'sd-0.18293737154261552, 32'sd-0.18570158101806397, 32'sd-0.09964789027858817, 32'sd0.047674595606089006, 32'sd0.027964780675863332, 32'sd0.10064673147824589, 32'sd-0.049487071130857416, 32'sd0.09430908650001592, 32'sd-0.016026506672393123, 32'sd0.010568790391368375, 32'sd0.015552891647217883, 32'sd0.026286550865036788, 32'sd0.06340389318018715, 32'sd-0.01110596128548924, 32'sd0.027007479419118855, 32'sd-0.0381237751762039, 32'sd-0.0058106960709133825, 32'sd-0.0697922317517589, 32'sd-2.773907381148774e-115, 32'sd0.052479293652692265, 32'sd0.05069589030652371, 32'sd-0.019305478419096495, 32'sd0.07487468680469517, 32'sd0.0742083755925363, 32'sd-0.12388993392419201, 32'sd-0.052226871744482053, 32'sd-0.04776632935246306, 32'sd-0.13204336169485073, 32'sd-0.058691204102286065, 32'sd-0.032942948019531126, 32'sd-0.010207677584188444, 32'sd-0.09696526373281009, 32'sd-0.07019523589311576, 32'sd-0.08595463185122383, 32'sd0.03263039404271636, 32'sd-0.04554864084768008, 32'sd0.08931678560422744, 32'sd0.07806017541293508, 32'sd-0.06524961386765869, 32'sd0.07030845912694009, 32'sd0.01923116671337368, 32'sd0.06828701581004218, 32'sd-0.0832126077836093, 32'sd0.04121946962278308, 32'sd-0.0608023325814033, 32'sd0.08474034364971031, 32'sd0.08771130968059468, 32'sd-0.008133744102124725, 32'sd-0.0018750403850289344, 32'sd-0.024975014766990197, 32'sd0.050092897961325614, 32'sd0.04499953238309415, 32'sd-0.010745622374929285, 32'sd-0.0113218590174679, 32'sd-0.02143073732745754, 32'sd-0.0625283511575957, 32'sd-0.0951549506028855, 32'sd-0.03982991548598258, 32'sd0.036962781190905056, 32'sd-0.07636590384184512, 32'sd0.012791206811224863, 32'sd0.047456453472323405, 32'sd0.049218191717808654, 32'sd0.05816216946548039, 32'sd0.025776757341627193, 32'sd0.010295673792485681, 32'sd-0.010946967878253142, 32'sd-0.034826484705480304, 32'sd0.09049469354216892, 32'sd-0.07268458511562884, 32'sd-0.016455711130527344, 32'sd0.06017046552398021, 32'sd0.03917768041967162, 32'sd-0.024410363982479606, 32'sd0.020601528030946562, 32'sd0.010338184872329001, 32'sd0.07838091487758937, 32'sd0.0177959347191572, 32'sd0.0594083633466805, 32'sd0.028669618495441435, 32'sd0.11085621225043933, 32'sd0.02157962983938423, 32'sd-0.01607417495595667, 32'sd-0.14652590358688414, 32'sd-0.01758949856255573, 32'sd-0.1377754809354816, 32'sd-0.018314539366356367, 32'sd0.08335056792019079, 32'sd-0.10122523871018964, 32'sd-0.04391494504628752, 32'sd0.10899715365274695, 32'sd0.003256766159620842, 32'sd-0.0734572200183515, 32'sd0.06944985141140625, 32'sd-0.020296607433645145, 32'sd-0.11377424057756731, 32'sd0.05757678359567234, 32'sd0.084955662563088, 32'sd-0.05481615833507423, 32'sd-0.011783417782088607, 32'sd-0.035649921644138265, 32'sd0.00016208121427534764, 32'sd0.01565146850029493, 32'sd0.022593403817178666, 32'sd-0.04672584359163451, 32'sd0.06718965127738884, 32'sd0.0193339684837756, 32'sd0.1248246377422293, 32'sd0.008397466083471396, 32'sd0.09952489738410102, 32'sd-0.04079506551473122, 32'sd-0.10220697771414505, 32'sd-0.0023482664600247187, 32'sd-0.048233181343038105, 32'sd-0.11454415535787525, 32'sd-0.09102063282243437, 32'sd-0.14726821396351839, 32'sd-0.05581629575481473, 32'sd0.0037178483571048172, 32'sd-0.1455571113447043, 32'sd-0.07762903402388419, 32'sd0.07393588818466099, 32'sd-0.019789796065541317, 32'sd-0.02911738643302867, 32'sd0.011984821090745786, 32'sd0.04765526590378938, 32'sd0.042738375542048776, 32'sd0.06197700718723604, 32'sd-0.01942310686878706, 32'sd-0.026152279141093644, 32'sd-0.030328244500297634, 32'sd-0.04044073773951961, 32'sd0.07997437390967838, 32'sd0.02021870571236561, 32'sd-0.03327269973770071, 32'sd0.14049939662786243, 32'sd0.20245747559965596, 32'sd0.1241019117988663, 32'sd-0.006906756337521763, 32'sd0.1166904913861268, 32'sd0.06832495517423348, 32'sd0.05157752697482296, 32'sd-0.06997687994169106, 32'sd-0.06730015862910424, 32'sd-0.07993400086528668, 32'sd-0.11161495629831794, 32'sd-0.04537336013488805, 32'sd-0.09227236850459387, 32'sd-0.07008191931851897, 32'sd-0.022246270846361917, 32'sd0.042969161256385814, 32'sd0.028768426099257418, 32'sd0.10511237724228634, 32'sd0.030490631229384953, 32'sd-0.021730050784936557, 32'sd-0.07881274338853046, 32'sd-0.08030416573317124, 32'sd0.0815599241250151, 32'sd-0.0347184668290212, 32'sd-0.05494982560447093, 32'sd0.05139609747181062, 32'sd0.0037034226660150674, 32'sd0.11185667836246671, 32'sd0.07090034699217819, 32'sd0.2299258156043813, 32'sd0.07326232511444225, 32'sd-0.004519003266989002, 32'sd0.13178416279360058, 32'sd0.08193329737559489, 32'sd0.11133250478676457, 32'sd-0.06141742488791228, 32'sd-0.0795888943285151, 32'sd-0.15388498893989938, 32'sd-0.0639769017450068, 32'sd0.034524607919996446, 32'sd0.02624665549480222, 32'sd-0.04122586837139954, 32'sd0.08567031237491325, 32'sd0.13999349864049362, 32'sd0.01397835966468646, 32'sd0.08405332340264797, 32'sd0.014387613139364142, 32'sd-0.008787105064610697, 32'sd-0.07155458173598488, 32'sd-0.09926471036338841, 32'sd-0.04626412818701123, 32'sd0.04690009481263867, 32'sd0.008936541074448485, 32'sd-0.0626088123605735, 32'sd-0.08712934667232876, 32'sd0.06044211145089039, 32'sd0.08339260123331368, 32'sd0.11558491872973223, 32'sd0.1998504226811549, 32'sd0.08609459460501488, 32'sd0.047007860332683706, 32'sd-0.011891992038668546, 32'sd0.03387262774781141, 32'sd0.047714497004444724, 32'sd-0.008935474063474148, 32'sd-0.08137600014037386, 32'sd-0.13589641816842726, 32'sd0.04639003942417795, 32'sd0.04757616012837932, 32'sd0.06916525550408592, 32'sd0.008132813077595462, 32'sd-0.03850769401086577, 32'sd0.046369683811370695, 32'sd0.012981132752851874, 32'sd-0.07256235741661946, 32'sd-0.0727041213106491, 32'sd-0.034871366813277946, 32'sd-0.114061210404576, 32'sd0.010924850639037467, 32'sd0.012264485201225627, 32'sd-0.005840134570972429, 32'sd0.0018908981207913802, 32'sd-0.057758558110661336, 32'sd-0.06051114602598991, 32'sd-0.16586209507416402, 32'sd-0.017664535056455752, 32'sd0.005188116609895098, 32'sd0.15524450064928078, 32'sd0.15933828250051138, 32'sd-0.03642204874091251, 32'sd-0.02816000176889803, 32'sd-0.17545861828658899, 32'sd-0.13387297718633207, 32'sd-0.03996221480731887, 32'sd-0.002265842890986254, 32'sd-0.02956578917075629, 32'sd-0.06881956770128972, 32'sd0.11202823923578079, 32'sd-0.03491983774257568, 32'sd-0.08592278296598135, 32'sd0.03359260076792348, 32'sd0.00615237661722637, 32'sd-0.029978276361260933, 32'sd-0.02996153902698383, 32'sd-0.07091140283930497, 32'sd-0.025604532057174847, 32'sd0.09932407031890704, 32'sd0.02802300378943037, 32'sd0.045982067766939555, 32'sd0.05638250182837741, 32'sd0.010716338369136272, 32'sd-0.07431729964093442, 32'sd-0.05160188248994933, 32'sd0.024690380505414913, 32'sd-0.054217860581642005, 32'sd-0.07323641231569702, 32'sd-0.15028116731615174, 32'sd-0.15882598445448431, 32'sd-0.1257847319430324, 32'sd-0.21652367039262546, 32'sd0.012210084426063441, 32'sd0.14098765282591105, 32'sd-0.08213911239731674, 32'sd0.016759202872036423, 32'sd-0.023145329017953967, 32'sd-0.12643116131275464, 32'sd-0.04216959893534948, 32'sd-0.01446129217738435, 32'sd-0.16189512298685702, 32'sd-0.13499150951598968, 32'sd0.04521439439308032, 32'sd-0.02813513899215082, 32'sd0.03427841561747757, 32'sd0.15500110117343857, 32'sd0.07070130050514503, 32'sd0.04313542718843079, 32'sd-0.07492995559957734, 32'sd0.004221005003320074, 32'sd0.06723373125130457, 32'sd0.04783062592490547, 32'sd-0.09022230735632605, 32'sd-0.04029884663663379, 32'sd-0.11436610802208522, 32'sd-0.22284198908885847, 32'sd-0.21654690263304194, 32'sd-0.2638600749726481, 32'sd-0.24106034127427234, 32'sd-0.10422039869829024, 32'sd0.06688028437624184, 32'sd0.17547317596699047, 32'sd-0.042680788549043884, 32'sd-0.029907463759010065, 32'sd-0.017766213380601505, 32'sd-0.004505915515950255, 32'sd-0.029101881658113494, 32'sd-0.12880111485561455, 32'sd-0.03978576538600398, 32'sd-0.0016822872598154712, 32'sd0.053118394662101165, 32'sd0.03970241419450415, 32'sd0.11909656033499834, 32'sd0.013561885239819806, 32'sd0.028330676911264042, 32'sd0.049261156103171756, 32'sd-0.06205819740411571, 32'sd-0.030081133685255737, 32'sd-0.022485406870089004, 32'sd0.10075793071673479, 32'sd-0.0023607299449700005, 32'sd-0.04965713670923848, 32'sd-0.05952661525141711, 32'sd-0.24930603206810178, 32'sd-0.30147961321662037, 32'sd-0.23736430092406374, 32'sd-0.09972990771917367, 32'sd0.004986551546605407, 32'sd0.1484622130118686, 32'sd0.14861738991591514, 32'sd0.03045419238725378, 32'sd0.11744888406884597, 32'sd-0.02095079819442637, 32'sd-0.03456172198380327, 32'sd-0.028831697077761113, 32'sd-0.08210211389803347, 32'sd-0.05926352986758735, 32'sd0.0001430272401348455, 32'sd0.1122789143060004, 32'sd0.017087484765893963, 32'sd-0.029625039659123123, 32'sd-0.10319087152516287, 32'sd-0.04336553692505312, 32'sd-1.0987905774501256e-122, 32'sd0.04563949427794038, 32'sd0.014562048562383866, 32'sd-0.04994891320557002, 32'sd-0.07259486254429177, 32'sd-0.11671346521677134, 32'sd-0.12544280727836163, 32'sd-0.2566308012135391, 32'sd-0.17515593559130962, 32'sd-0.21545894600136406, 32'sd-0.11065456821811957, 32'sd0.08370350632878293, 32'sd0.26721013054594595, 32'sd0.05813879606034499, 32'sd0.09847893428733955, 32'sd-0.045414614618864584, 32'sd0.06540217406964471, 32'sd0.11413567095241839, 32'sd0.07605669340189711, 32'sd-0.03321035187217564, 32'sd0.03530683480006967, 32'sd-0.1568922903895998, 32'sd-0.010393847901149562, 32'sd0.022362659224945094, 32'sd-0.014002045028232138, 32'sd-0.10182647083878807, 32'sd-0.10921679539673958, 32'sd0.030924825548692882, 32'sd-0.02301452068942507, 32'sd0.06898888717015203, 32'sd-0.10141538300083201, 32'sd-0.035770979406925876, 32'sd0.04328666489647579, 32'sd-0.08169739314094981, 32'sd-0.07654852780755497, 32'sd-0.30526691481016327, 32'sd-0.2565701846325001, 32'sd-0.1032124808439495, 32'sd0.1209284451986448, 32'sd0.11921424735274279, 32'sd0.26944316064094986, 32'sd0.20282642707795615, 32'sd-0.08635666321010634, 32'sd-0.09328504327297825, 32'sd-0.1388081454071575, 32'sd-0.0125463285168084, 32'sd0.009985038436275098, 32'sd0.06717497243506564, 32'sd-0.11161817361877295, 32'sd-0.14723441353789551, 32'sd-0.12400998206132584, 32'sd-0.06109142922578699, 32'sd0.04974134758501961, 32'sd-0.010681895819642953, 32'sd-0.050475018834400656, 32'sd-0.03046799742268942, 32'sd0.028401425795383878, 32'sd-0.08401566170913659, 32'sd-0.052548672479841615, 32'sd0.0807770194464514, 32'sd-0.043978186416135566, 32'sd-0.15457311514109515, 32'sd-0.1550711598505307, 32'sd-0.10297309029444703, 32'sd-0.07202541061011268, 32'sd0.048284514397156614, 32'sd0.05545541865449347, 32'sd0.14432145439542807, 32'sd0.1691656548118818, 32'sd0.0946199930151126, 32'sd-0.09213768296923253, 32'sd-0.1233242782253545, 32'sd-0.02813211320133642, 32'sd0.037148585149838625, 32'sd0.02950562810179788, 32'sd0.03403386757872961, 32'sd0.018576295846518463, 32'sd-0.013064022573294892, 32'sd-0.08714671543287203, 32'sd-0.07681967907984949, 32'sd-0.013219449667589851, 32'sd-0.11088247660030007, 32'sd-0.03871808756770202, 32'sd0.051296196118292614, 32'sd2.3769541022681145e-117, 32'sd-0.03151329691044663, 32'sd0.016866465186535427, 32'sd0.01234658906212967, 32'sd-0.061361395811275164, 32'sd-0.14211015129219312, 32'sd-0.15391937678933892, 32'sd-0.06229127790170974, 32'sd-0.028954555284398106, 32'sd-0.015877815036219378, 32'sd0.09355379625244585, 32'sd0.19981123189489938, 32'sd0.26272853864696505, 32'sd-0.014482584627755882, 32'sd0.02196306408567467, 32'sd0.02997897459055173, 32'sd0.04543528262790993, 32'sd0.04889243658417773, 32'sd0.1298072352752385, 32'sd0.01934173896722372, 32'sd-0.08722834102570849, 32'sd0.049445878076025615, 32'sd-0.09967765481165007, 32'sd-0.06465679236515938, 32'sd-0.07249408063645917, 32'sd-0.047243224296861355, 32'sd-0.050353157697540944, 32'sd0.04334754415103735, 32'sd0.09853979724473197, 32'sd0.0505145612502992, 32'sd0.03779390710530395, 32'sd-0.0182754842336188, 32'sd-0.09174462159611076, 32'sd0.0022710578606346455, 32'sd0.037383075704863794, 32'sd-0.039303490366830805, 32'sd-0.16904075083534922, 32'sd-0.009910202116168191, 32'sd0.02932710491301129, 32'sd0.07253050230087386, 32'sd0.15105903805030904, 32'sd0.015545897685424947, 32'sd0.027678257527273604, 32'sd0.06102614957992224, 32'sd0.05588208131632185, 32'sd0.08756641677462478, 32'sd0.07362167041827077, 32'sd0.10353077190977429, 32'sd-0.008705531106565198, 32'sd0.013940350805317176, 32'sd0.04651145644507429, 32'sd0.09549779550766085, 32'sd0.14187796770689667, 32'sd0.052713818318256826, 32'sd0.08000305008173042, 32'sd0.02516726432007522, 32'sd0.05470004322807032, 32'sd-0.030393587734287374, 32'sd-0.025446297404228557, 32'sd-0.05958664693762823, 32'sd0.026269291485481936, 32'sd-0.011063198047647002, 32'sd-0.015499637859201248, 32'sd-0.043924727404069656, 32'sd-0.16125467111576625, 32'sd0.011838697140109097, 32'sd-0.01277060336016615, 32'sd0.009916264745055133, 32'sd0.07484114701338744, 32'sd0.015962122434247456, 32'sd-0.05192343260225715, 32'sd-0.03876480850795294, 32'sd0.07209477328016374, 32'sd0.13153911074009902, 32'sd0.16026008036929507, 32'sd0.025433751052443613, 32'sd-0.07406909257685533, 32'sd-0.060495586850548046, 32'sd0.11584745777304949, 32'sd0.03992348697243953, 32'sd-0.001137265946444413, 32'sd0.05385483275146987, 32'sd0.07168758754214129, 32'sd0.037680732631483825, 32'sd1.4144352884607384e-118, 32'sd0.04972336761574943, 32'sd0.03819201995208316, 32'sd-0.06062200100882724, 32'sd-0.1094052842677378, 32'sd-0.029794694280926293, 32'sd0.0335113533942506, 32'sd0.02272513534826076, 32'sd-0.10527402659096854, 32'sd0.03403929612216842, 32'sd-0.06798104053503763, 32'sd0.0536022364452477, 32'sd0.03124313112429969, 32'sd0.13494918446017665, 32'sd0.045938357468822244, 32'sd0.16515473966516542, 32'sd0.07357675528396723, 32'sd0.08727853774125575, 32'sd0.003961131790941677, 32'sd0.09415823151827472, 32'sd0.027695317898530657, 32'sd-0.11868233054382989, 32'sd-0.0018897831638966544, 32'sd0.09995399424541496, 32'sd0.03209569823092608, 32'sd0.04202476112713764, 32'sd-0.02256230659861966, 32'sd-6.609120421303877e-128, 32'sd1.2950589690785086e-122, 32'sd6.046804456313183e-127, 32'sd-0.002092695788932614, 32'sd-0.07945218001921814, 32'sd-0.15653759767223258, 32'sd-0.050380258696947997, 32'sd-0.002895945288450113, 32'sd-0.09127315604705204, 32'sd-0.015520901315499491, 32'sd-0.08175698892210867, 32'sd-0.1081058407930244, 32'sd0.007951470778968845, 32'sd0.10839431311223036, 32'sd0.04599179450057663, 32'sd0.09504958655917427, 32'sd0.03144163545395423, 32'sd0.027542253872953715, 32'sd-0.037556720446042774, 32'sd0.07150875643358076, 32'sd0.08868024090772313, 32'sd0.08262633081540588, 32'sd-0.05479947375218958, 32'sd0.004626334079598281, 32'sd0.05104707359380123, 32'sd0.06346475970141731, 32'sd0.0743415238591581, 32'sd0.035106307502328876, 32'sd-2.957152810049522e-122, 32'sd3.4538780978267534e-124, 32'sd-1.0735667743659295e-121, 32'sd-0.023297814510036416, 32'sd0.032981688427156326, 32'sd0.05694493259737649, 32'sd0.020556076583331404, 32'sd0.12649040390774272, 32'sd-0.05209641781827804, 32'sd-0.044790025110743106, 32'sd-0.017380168803094696, 32'sd-0.06572461333132629, 32'sd0.009195474459976913, 32'sd0.07612707530866411, 32'sd-0.002484186507368407, 32'sd0.10600315149339315, 32'sd0.13197401634326536, 32'sd-0.051093590095889686, 32'sd0.003199764066484337, 32'sd-0.11774439934067876, 32'sd-0.03394009458922504, 32'sd-0.02621241585262256, 32'sd0.012323035848460477, 32'sd-0.09175774721618256, 32'sd-0.048618207600199595, 32'sd-0.00013916785796462756, 32'sd-0.0006059463564529071, 32'sd-0.002240899654951382, 32'sd-3.146124211752444e-120, 32'sd1.0715816638217655e-124, 32'sd-3.678475451195781e-125, 32'sd1.5727578729595705e-121, 32'sd0.033652102682019305, 32'sd-0.031444859071945504, 32'sd-0.006102133806258932, 32'sd0.045455080606562386, 32'sd-0.0465470551403973, 32'sd0.08890334929174339, 32'sd-0.008977142296598295, 32'sd0.000858540734612017, 32'sd0.07199446674129895, 32'sd-0.02354805366605972, 32'sd-0.041562197269530025, 32'sd-0.14033695016774764, 32'sd-0.06903446151574814, 32'sd-0.09346450289029795, 32'sd0.03817657764668774, 32'sd0.05255983421311176, 32'sd0.037022662397332165, 32'sd0.042393331527682834, 32'sd-0.0614898822499989, 32'sd0.1230924710879739, 32'sd0.03647148303601066, 32'sd-0.03590554609682272, 32'sd0.041786377774367986, 32'sd-4.659312152674603e-122, 32'sd1.2914817420655066e-124, 32'sd1.0974686055760086e-121, 32'sd3.385638638965049e-120, 32'sd-5.337919029845709e-118, 32'sd-3.209516138599097e-120, 32'sd0.10353199204284422, 32'sd0.06063508140692834, 32'sd-0.010411964067822724, 32'sd0.10129493518849939, 32'sd-0.05167592265016883, 32'sd-0.011345693494695436, 32'sd-0.050754254582259295, 32'sd0.005089862585719971, 32'sd0.05782810751911301, 32'sd0.11143805554638052, 32'sd0.1338094676754687, 32'sd0.06488019139684613, 32'sd0.1783305741319779, 32'sd0.11980308986323523, 32'sd0.05026120177632877, 32'sd0.07121283651270895, 32'sd0.00591541130834709, 32'sd0.02398213846107938, 32'sd0.012900760776877651, 32'sd0.003351748008616799, 32'sd2.330813102546962e-120, 32'sd-6.25617283880024e-118, 32'sd3.5631767228916125e-123, 32'sd4.905117906201472e-121},
        '{32'sd6.732116446403674e-124, 32'sd-9.281838966427261e-116, 32'sd-3.4624001693795927e-127, 32'sd-1.6829041375427163e-122, 32'sd3.1752140249221695e-120, 32'sd-1.6338020187035127e-121, 32'sd1.7696462110798766e-123, 32'sd1.7823793651550075e-123, 32'sd2.168584850493359e-125, 32'sd-7.128073565096033e-120, 32'sd3.6825322011012354e-122, 32'sd-9.61803207290355e-120, 32'sd-0.016908596970013633, 32'sd0.04499167840669021, 32'sd0.12168253861251552, 32'sd0.088856441607883, 32'sd-2.66357139586753e-117, 32'sd-1.1010503483914126e-128, 32'sd2.210997893159552e-116, 32'sd-1.3168496140150083e-125, 32'sd4.049171289532105e-115, 32'sd4.749326945104765e-118, 32'sd1.631600910327852e-115, 32'sd-1.0909487579023378e-119, 32'sd-1.1505752171994648e-116, 32'sd9.350132632698658e-120, 32'sd9.423607395453278e-120, 32'sd-3.206176135404008e-116, 32'sd-1.5406414850046975e-117, 32'sd-7.99454095750822e-121, 32'sd-2.535137007615012e-126, 32'sd1.3337738564048308e-118, 32'sd0.013227747992152922, 32'sd0.003460210355183451, 32'sd0.058158375809056806, 32'sd-0.051918767692888765, 32'sd0.04506468295676758, 32'sd0.046798504686800656, 32'sd0.0701195749840739, 32'sd0.06689971248634662, 32'sd-0.01903671622837241, 32'sd-0.053348869828272596, 32'sd0.041128035028332725, 32'sd-0.036771098110812174, 32'sd0.08541725131989888, 32'sd5.4777866540324977e-05, 32'sd0.026820820096302857, 32'sd0.0517450058182802, 32'sd-0.02455058594624474, 32'sd0.08344526751712074, 32'sd0.08952777428740269, 32'sd0.07437806502149115, 32'sd-3.027188089256357e-118, 32'sd-6.746828222756826e-126, 32'sd-3.9050625076093604e-119, 32'sd-2.835403634242706e-116, 32'sd-5.663655615824547e-127, 32'sd-2.8369537707393255e-123, 32'sd0.057686242043054115, 32'sd0.0519864992236797, 32'sd-0.11488142628119563, 32'sd0.07913466367133876, 32'sd0.07650537281241984, 32'sd0.07341609530846023, 32'sd0.01726743783475123, 32'sd0.012525600773306337, 32'sd0.020840094960799697, 32'sd-0.0365230957814003, 32'sd-0.019878480570740927, 32'sd-0.05702061355649037, 32'sd-0.033916049683308115, 32'sd-0.11372667898470966, 32'sd0.02294580984973814, 32'sd0.14270197994108633, 32'sd0.10642627625418666, 32'sd-0.15536034214665967, 32'sd-0.1222446312753069, 32'sd0.08316241757507005, 32'sd0.030628237891809126, 32'sd0.06742380938218699, 32'sd0.07145357349881269, 32'sd0.08492238583956539, 32'sd5.9175790015621486e-124, 32'sd3.292297998039331e-119, 32'sd-1.9751511242823612e-126, 32'sd2.2644116982066004e-126, 32'sd0.08093072352381231, 32'sd-0.02014396509999494, 32'sd-0.02224327813149212, 32'sd0.022826121041561412, 32'sd0.00781049873591478, 32'sd-0.056454814033471606, 32'sd0.0009345759523649151, 32'sd-0.0313369176936752, 32'sd0.05470315493880158, 32'sd0.012056131620749647, 32'sd0.06757135987360138, 32'sd0.0857766656094864, 32'sd0.06347292981536982, 32'sd-0.07957573863542, 32'sd0.027457032634686032, 32'sd0.016857683803306194, 32'sd0.08043293689189311, 32'sd0.04488153122614102, 32'sd-0.05668862541178325, 32'sd0.04698147583100479, 32'sd0.03989358072524248, 32'sd-0.058833714193319696, 32'sd-0.028883621916436477, 32'sd0.026349293094473897, 32'sd-0.10021781526148614, 32'sd-4.6293078375411567e-126, 32'sd4.258809271500359e-118, 32'sd-0.0014480154346317381, 32'sd0.04276879369816518, 32'sd0.012430903705406024, 32'sd0.08126448760309568, 32'sd-0.01666027370244736, 32'sd0.06112674113847732, 32'sd-0.02423826739701892, 32'sd0.020114603316105133, 32'sd-0.05038772093728931, 32'sd0.006738051620031507, 32'sd0.08863864189466795, 32'sd0.10640499912569555, 32'sd0.10764331365847957, 32'sd-0.017953386641797416, 32'sd-0.03068122942659164, 32'sd-0.0012829009972640357, 32'sd-0.12533297799526386, 32'sd-0.06653162288570214, 32'sd-0.1307824150901775, 32'sd-0.03341789787089594, 32'sd0.007345718366959393, 32'sd-0.0630015061609659, 32'sd0.00613576613418038, 32'sd0.06225664120371307, 32'sd-0.008669403073196297, 32'sd-0.057662416140162764, 32'sd0.07746898290018683, 32'sd2.8603530166777552e-118, 32'sd0.0514956203238144, 32'sd-0.03459373021384479, 32'sd-0.04590682075514602, 32'sd0.08602874590364601, 32'sd0.05784344595126574, 32'sd0.035042276598133304, 32'sd0.04557455123990819, 32'sd0.12593541774714365, 32'sd0.00950789962377158, 32'sd0.15632882312973218, 32'sd0.21576989447427283, 32'sd0.22545744189544026, 32'sd0.05736707258838734, 32'sd0.14351794890741756, 32'sd-0.036900621088564234, 32'sd0.060826829597786077, 32'sd-0.020867107851165433, 32'sd-0.20286607956619634, 32'sd-0.15982393114936327, 32'sd-0.061781371619724, 32'sd0.06061587531197238, 32'sd-0.01329349457028168, 32'sd0.0989774302491024, 32'sd0.05186505933334916, 32'sd0.020638827247243013, 32'sd-0.07508587904740324, 32'sd0.035929938270911545, 32'sd2.608649210350136e-124, 32'sd0.0412412745097449, 32'sd0.010632565569227334, 32'sd0.05827943374515469, 32'sd-0.0197459298494883, 32'sd0.0630423500489864, 32'sd0.0770029850191475, 32'sd0.07404735976906833, 32'sd0.16871618237505037, 32'sd0.11003391566426755, 32'sd0.22951124497528258, 32'sd0.10085042801127903, 32'sd0.19518785527439908, 32'sd0.07739187941881372, 32'sd-0.07554388641188092, 32'sd0.018066007815878807, 32'sd-0.06927133333805309, 32'sd0.04616983177568627, 32'sd-0.028326885259727888, 32'sd0.02564436998796911, 32'sd-0.04038183219027492, 32'sd-0.07138920114928662, 32'sd0.051759714218046336, 32'sd-0.0031604310647261272, 32'sd0.13253165218423985, 32'sd0.058057081857237444, 32'sd-0.052825945139669137, 32'sd-0.002570320468665741, 32'sd0.12065597978464607, 32'sd0.047382021271622776, 32'sd4.9330144519322884e-05, 32'sd0.05480508897402209, 32'sd0.11596821866386584, 32'sd0.12555506760037768, 32'sd0.02446168939060171, 32'sd0.029088137902943144, 32'sd0.04074369563257996, 32'sd0.2186670058061406, 32'sd0.21126444516620205, 32'sd0.1261413158693698, 32'sd0.04854735629461514, 32'sd0.02641350687338776, 32'sd-0.14385318346094014, 32'sd-0.14701449777758613, 32'sd-0.004007499423646708, 32'sd0.12057583523504856, 32'sd0.047730728826667526, 32'sd-0.04117339233920538, 32'sd-0.004486511432595136, 32'sd-0.05841924137577098, 32'sd-0.031166732281462026, 32'sd-0.040929771435198554, 32'sd0.216756858539231, 32'sd0.09456231120226202, 32'sd0.009220168082626207, 32'sd-0.009863596673890715, 32'sd0.07314106062124263, 32'sd0.09007809639225807, 32'sd-0.006302054960014969, 32'sd0.13290984867026895, 32'sd0.11040084820902009, 32'sd0.0722660979192567, 32'sd0.13578668164685045, 32'sd0.10197284223868408, 32'sd0.010405332227066817, 32'sd0.15031251288959974, 32'sd0.12291726813013741, 32'sd0.023314176299842757, 32'sd0.04925011999854331, 32'sd0.14008374026636575, 32'sd-0.08056140674462757, 32'sd-0.11829446874746109, 32'sd0.00866104933929197, 32'sd0.07503602509098953, 32'sd0.153073854241814, 32'sd-0.006897201761892293, 32'sd0.027273360996190318, 32'sd-0.13394093690393388, 32'sd-0.007702565799313091, 32'sd0.12683801873619768, 32'sd0.18593875126828063, 32'sd0.03268344742001818, 32'sd0.0010348458653871655, 32'sd0.008347664058356649, 32'sd0.04305039886167, 32'sd0.0013347493304828764, 32'sd0.15145775905251535, 32'sd0.1301654633709807, 32'sd-0.05563289602348509, 32'sd-0.0636484766717629, 32'sd-0.16279138867667772, 32'sd-0.14014017061454143, 32'sd-0.0780695608858614, 32'sd-0.01771445145002098, 32'sd0.0005199703671925499, 32'sd0.0004253620585746198, 32'sd0.05056681393279382, 32'sd-0.01956272093221968, 32'sd0.020607985405211304, 32'sd-0.04169710208056888, 32'sd-0.07867105548342238, 32'sd0.17920268834834938, 32'sd-0.03881385173699406, 32'sd-0.10548791302955896, 32'sd0.017330221557854394, 32'sd0.11017615568500458, 32'sd-0.023583627003218074, 32'sd0.1379161408823695, 32'sd0.05844565080564931, 32'sd0.032703957725061905, 32'sd-0.022811595835259425, 32'sd0.07128156570102075, 32'sd0.08032861364216384, 32'sd0.03787184900972134, 32'sd-0.017607467952387976, 32'sd0.09493048137417003, 32'sd-0.05699437481202473, 32'sd-0.10090933433804576, 32'sd-0.059138302905713924, 32'sd-0.18415357878451752, 32'sd-0.17388944295701395, 32'sd-0.07721643778427249, 32'sd0.05703951955895357, 32'sd-0.03159606183482359, 32'sd-0.11629381399127292, 32'sd-0.09124384031119855, 32'sd-0.19029976499614992, 32'sd0.055153961242629806, 32'sd0.023249319555187664, 32'sd0.1423713325647348, 32'sd0.012840336209883502, 32'sd-0.01652049286039868, 32'sd-0.04637382708055024, 32'sd-0.041586652922766774, 32'sd0.07400488600000786, 32'sd0.055717140202228, 32'sd0.01358089184403285, 32'sd-0.03340957184841783, 32'sd0.015273864680544888, 32'sd-0.0070368901281057114, 32'sd0.09254439390438088, 32'sd-0.013442977534691475, 32'sd0.040763925960947814, 32'sd-0.04532978257979864, 32'sd-0.09744752763401887, 32'sd-0.0647839091901819, 32'sd-0.16548573215253448, 32'sd-0.14388437867358972, 32'sd-0.08060144445115304, 32'sd0.014894339890804168, 32'sd-0.018373487588622634, 32'sd-0.09164765040250648, 32'sd0.00979228103689952, 32'sd-0.027429826160087812, 32'sd-0.11029851141562784, 32'sd-0.0601308929590329, 32'sd-0.010479849420042951, 32'sd0.0044505335540534685, 32'sd0.0451358541253532, 32'sd-0.08937284902192506, 32'sd-0.10968790501310186, 32'sd0.003437882114311356, 32'sd0.013872346636481073, 32'sd-0.018277687010934397, 32'sd0.0033285935121993124, 32'sd0.012626311655068067, 32'sd0.0007597974527210263, 32'sd0.023190842595327513, 32'sd0.05424165168345842, 32'sd0.07251113150123654, 32'sd0.06515503372994368, 32'sd-0.03986181633149828, 32'sd-0.03222886929034926, 32'sd-0.1980211473106865, 32'sd-0.21454740518058868, 32'sd-0.22194309666705525, 32'sd-0.12428930625361011, 32'sd-0.22277795257669486, 32'sd-0.14002542456214323, 32'sd-0.11232074264049896, 32'sd-0.02604401474681225, 32'sd0.028060955352205017, 32'sd-0.10368287923192641, 32'sd0.04794062764978668, 32'sd0.15488148379618535, 32'sd0.04940646726439099, 32'sd0.06346100107127403, 32'sd0.02183627249990914, 32'sd0.029364503967072655, 32'sd-0.007210500580575307, 32'sd-0.0075600363733832185, 32'sd0.05128224239080114, 32'sd0.10347313281102459, 32'sd0.004741203403679011, 32'sd-0.01891489847463465, 32'sd-0.004879012643198605, 32'sd0.06913856795299725, 32'sd0.0872127803363104, 32'sd0.07111268696089491, 32'sd0.029443132444210957, 32'sd-0.10810713418311992, 32'sd-0.15499803138841042, 32'sd-0.2558272975464294, 32'sd-0.1773106838472283, 32'sd-0.1483395045209753, 32'sd-0.16948716191308758, 32'sd0.05018312958354582, 32'sd0.02951039744539432, 32'sd0.08133812227572636, 32'sd0.10524863233259503, 32'sd-0.11582807523899948, 32'sd-0.0393503630853665, 32'sd0.05976254282337651, 32'sd-0.1299564694278023, 32'sd-0.023977062009649785, 32'sd0.024020416105905253, 32'sd0.04450018173725728, 32'sd0.07207434248970195, 32'sd0.037739878674104485, 32'sd-0.006692796492108261, 32'sd0.045449745083423185, 32'sd-0.13568561696314965, 32'sd-0.06643085007473873, 32'sd0.033868755147119387, 32'sd-0.02271813129635767, 32'sd-0.04944901625378842, 32'sd0.0316687457801118, 32'sd-0.056610919243487504, 32'sd0.08511237509911646, 32'sd-0.04895480390292839, 32'sd-0.03898460503565113, 32'sd-0.21915848244011119, 32'sd-0.22675651046206105, 32'sd-0.17527941081298232, 32'sd0.10292225955917313, 32'sd0.11874254171089779, 32'sd0.10854737870909992, 32'sd0.020645421581439328, 32'sd-0.03161141132888914, 32'sd-0.006218915703662149, 32'sd-0.1517758273006658, 32'sd-0.061450617750118945, 32'sd-0.0059843955163856564, 32'sd0.004504526505992762, 32'sd-0.06006837027353484, 32'sd0.07072055306143928, 32'sd-0.09057692132574385, 32'sd-0.09621223255093124, 32'sd-0.07128774930045031, 32'sd0.1373409623245855, 32'sd-0.048280172164544534, 32'sd-0.04303171207412559, 32'sd0.09185696131463622, 32'sd0.021669739378818928, 32'sd0.0745934535483753, 32'sd0.10790826039196563, 32'sd0.042263240419970316, 32'sd-0.06307355765797379, 32'sd0.0419886334720814, 32'sd0.013917379466618463, 32'sd-0.13472245681464837, 32'sd-0.0013513362501885737, 32'sd0.09470341519146762, 32'sd0.13602992695373256, 32'sd-0.030775181641532912, 32'sd0.00887532373915429, 32'sd-0.01947993023946328, 32'sd0.06856505870891832, 32'sd-0.039605156104189555, 32'sd0.004122759030274769, 32'sd0.08470100670810353, 32'sd0.004131505535499615, 32'sd0.010640021839904486, 32'sd0.07072634107448224, 32'sd-0.007563406745015133, 32'sd0.0864308999936443, 32'sd0.06977589540123512, 32'sd0.17594085822305977, 32'sd0.05549416981765539, 32'sd-0.025816369345555416, 32'sd0.07073220008961174, 32'sd-0.08312047449537405, 32'sd0.03598128530620854, 32'sd0.05280530197031611, 32'sd-0.08537642240434873, 32'sd0.09782071613230515, 32'sd-0.014633304847373326, 32'sd0.1319867881923445, 32'sd0.025964129339542057, 32'sd0.07448879407690116, 32'sd0.12030783595855339, 32'sd-0.039795957024838964, 32'sd-0.03182131761177254, 32'sd0.040337273829026, 32'sd0.020450417108029587, 32'sd-0.043603055224320904, 32'sd-0.03752928419253492, 32'sd0.14016781652088386, 32'sd0.07387769871415768, 32'sd0.10198250891479584, 32'sd-0.01152431022016063, 32'sd0.1246735353223659, 32'sd0.04201598570273828, 32'sd0.01820695946609011, 32'sd0.04035050536398644, 32'sd0.09071032329532375, 32'sd0.058597034362453226, 32'sd0.024632896917825522, 32'sd-4.3137477090548743e-125, 32'sd0.008092036758131149, 32'sd-0.02004145435422983, 32'sd-0.02173718707968618, 32'sd0.038778383348368674, 32'sd-0.026923431759272365, 32'sd-0.006347474823047792, 32'sd0.05913703236169181, 32'sd-0.023788891148898286, 32'sd0.15201370930976701, 32'sd0.02625560218137382, 32'sd0.021336369153959613, 32'sd0.014670950563552528, 32'sd-0.0005530865430238804, 32'sd-0.03358799469479333, 32'sd-0.07014715065233215, 32'sd-0.004904699782221141, 32'sd-0.120813139597439, 32'sd-0.030966524910383198, 32'sd0.04753938625830603, 32'sd0.06401414938118376, 32'sd0.059206666887650174, 32'sd-0.006198983175522359, 32'sd-0.021838189810951234, 32'sd-0.033984677711623966, 32'sd0.04843640503101052, 32'sd0.002008474191874838, 32'sd-0.016465272125948074, 32'sd-0.014470940487817621, 32'sd-0.011760022328677028, 32'sd-0.0258344651170674, 32'sd0.008932469261632398, 32'sd0.07800914792971211, 32'sd0.006981029388598817, 32'sd-0.06107759055255915, 32'sd0.017968525181594287, 32'sd-0.004175755717213733, 32'sd0.06316989288076377, 32'sd0.03190740709649352, 32'sd0.07225181081719767, 32'sd0.04432709996807674, 32'sd-0.0206234493707881, 32'sd-0.1364266371998578, 32'sd-0.003748916515741194, 32'sd-0.14185948106641458, 32'sd-0.057973652934539543, 32'sd0.010002584250735013, 32'sd-0.043012049828888475, 32'sd-0.0629757276560846, 32'sd-0.10451016772787453, 32'sd-0.015955210547231525, 32'sd0.03802591248157834, 32'sd0.053661224373955124, 32'sd0.02235475797086033, 32'sd0.04419812744285702, 32'sd0.026571478054982476, 32'sd0.05424782799691146, 32'sd0.0141008348965758, 32'sd0.07188639551798522, 32'sd0.09883369036413812, 32'sd0.020641471139052365, 32'sd0.01554197615625078, 32'sd-0.1313696522132445, 32'sd-0.07581706855714603, 32'sd-0.053976268832017636, 32'sd-0.0005979192775043207, 32'sd0.03445755571282676, 32'sd0.22188294354023444, 32'sd0.015352877863166577, 32'sd0.06933596198041017, 32'sd0.04594663882932524, 32'sd0.07006349974525518, 32'sd-0.09354920800920777, 32'sd-0.03689752950206818, 32'sd0.03448281174966995, 32'sd0.032209833959274896, 32'sd-0.0008374238142771002, 32'sd-0.0470397069966225, 32'sd0.07932353390262874, 32'sd0.05949770802976569, 32'sd0.036289651572065304, 32'sd-0.0007774065493128307, 32'sd0.010920439216107298, 32'sd-0.015005910596756785, 32'sd5.227425398890271e-127, 32'sd0.05760426318602416, 32'sd0.015273836198959676, 32'sd0.049353109680500905, 32'sd-0.1027615236900709, 32'sd-0.010503280955391957, 32'sd-0.1311179273333329, 32'sd-0.13237722579045735, 32'sd0.00740874908665986, 32'sd-0.08076005154671226, 32'sd0.07643929009809108, 32'sd0.1253398242398287, 32'sd0.018120432040630702, 32'sd0.04381417980255461, 32'sd-0.053519815699584986, 32'sd0.016643221887617066, 32'sd-0.11792579834342956, 32'sd-0.03879228769511194, 32'sd-0.11968010002696787, 32'sd-0.08073097351111894, 32'sd-0.09274233613378263, 32'sd-0.04050797539862884, 32'sd-0.07533652727362167, 32'sd0.03430290454211453, 32'sd0.001277079237866609, 32'sd0.0031809879656274002, 32'sd-0.05660398228917151, 32'sd0.043629255723854794, 32'sd0.04379817835993853, 32'sd-0.0334553761441087, 32'sd0.01671621367419, 32'sd0.05659327059479403, 32'sd-0.04340385846329173, 32'sd-0.06685303227193823, 32'sd-0.1555788558316307, 32'sd-0.13696768745226048, 32'sd-0.08368695721013043, 32'sd-0.07449470569874796, 32'sd0.035488760183355665, 32'sd0.09917806438618984, 32'sd0.01814611037801306, 32'sd0.11087497533417673, 32'sd0.1508515813603204, 32'sd0.05655474109693482, 32'sd-0.018291912531424308, 32'sd-0.08375828936147175, 32'sd-0.1171622712379619, 32'sd0.05023354764096265, 32'sd-0.15679237737309576, 32'sd0.020568236643021893, 32'sd0.11171857192601009, 32'sd0.07490662527560844, 32'sd-0.014562434305509301, 32'sd0.10795160679113805, 32'sd0.007658153233694876, 32'sd0.03993603243277676, 32'sd-0.023780779683346038, 32'sd-0.10936451124242796, 32'sd0.12079649912522245, 32'sd0.04342839080598917, 32'sd0.0823159396713821, 32'sd-0.04735748088780424, 32'sd-0.12128600934172999, 32'sd0.033506725916009165, 32'sd-0.0623038525502858, 32'sd-0.09187077069814854, 32'sd0.013183781614904518, 32'sd0.05664538477094408, 32'sd0.14071183205302465, 32'sd0.0959835253328929, 32'sd-0.07490632314551976, 32'sd-0.05456060709502551, 32'sd-0.0463371246677214, 32'sd-0.071581723412957, 32'sd-0.1535530938680007, 32'sd-0.12833599783685007, 32'sd0.04215024471144471, 32'sd0.09276560551471144, 32'sd0.0343090290378977, 32'sd0.030764213596110288, 32'sd-0.042434962774908276, 32'sd-0.029359247054358457, 32'sd-0.10355948886618356, 32'sd-0.03558890094073797, 32'sd-3.803177030627133e-129, 32'sd0.0820844403341878, 32'sd0.15339849061046154, 32'sd0.05103603458724059, 32'sd0.06397357925553161, 32'sd-0.1295379198179875, 32'sd-0.18039307775869937, 32'sd-0.030065691821097015, 32'sd-0.05540198243442426, 32'sd-0.07302047215325189, 32'sd0.043618041090735554, 32'sd0.0279960668462676, 32'sd-0.03636627841938352, 32'sd0.027133255768048575, 32'sd-0.02717219747472511, 32'sd-0.01773412385105868, 32'sd-0.013219485131119098, 32'sd-0.05059827700716602, 32'sd-0.07071722269675082, 32'sd0.04645345488064205, 32'sd-0.050320897305234924, 32'sd-0.05008146245832187, 32'sd-0.08447070633969969, 32'sd-0.09353077840432747, 32'sd-0.10012135435620606, 32'sd0.02918859067167182, 32'sd0.008749685750393985, 32'sd1.6935856241818216e-123, 32'sd-7.361961789994266e-115, 32'sd2.5437585729454966e-123, 32'sd0.0007443720476090817, 32'sd0.06357731183996672, 32'sd0.006090516283805771, 32'sd-0.09435317521781954, 32'sd-0.07977096565273184, 32'sd-0.008412057441426733, 32'sd0.14292686895688217, 32'sd0.0003112438269577305, 32'sd-0.06860857977657756, 32'sd0.01758223064479076, 32'sd0.020876227110673693, 32'sd0.10766390052043505, 32'sd0.14774070298136355, 32'sd-0.001892031806147659, 32'sd-0.07653254431497598, 32'sd0.028127275901825694, 32'sd-0.06014733775604359, 32'sd-0.03884169926837917, 32'sd-0.031585402230870765, 32'sd-0.16733807075387622, 32'sd0.05856092353101637, 32'sd-0.0216916596740463, 32'sd-0.004785048307508368, 32'sd0.002838885918730584, 32'sd0.062442269178666854, 32'sd1.6495074250630158e-125, 32'sd3.3126798740225455e-121, 32'sd-6.885911588259468e-120, 32'sd0.03892169097797964, 32'sd0.0085935316981027, 32'sd-0.0236130944573639, 32'sd0.03508293304396086, 32'sd-0.012003276075961617, 32'sd0.13283064582691945, 32'sd-0.024241660874805646, 32'sd-0.0498675874639817, 32'sd-0.052977913077943035, 32'sd0.041360114149850274, 32'sd0.009106888078307708, 32'sd0.02429551294294061, 32'sd-0.018352974406165692, 32'sd0.18522510333373443, 32'sd0.16822750922354238, 32'sd0.16060407560559428, 32'sd0.07742588951400056, 32'sd0.08491253082034257, 32'sd0.00569004048739743, 32'sd-0.03674446057125562, 32'sd-0.07103593412686697, 32'sd-0.10677530414287785, 32'sd0.042015705145977626, 32'sd0.003136683906899575, 32'sd0.01735087481076601, 32'sd-6.122452468606258e-124, 32'sd1.0765433919332954e-124, 32'sd8.086867829512829e-117, 32'sd5.392654843966017e-115, 32'sd0.12171711105718079, 32'sd-0.019703915875408564, 32'sd-0.012627737754063837, 32'sd-0.12805016501860433, 32'sd-0.02622101590061677, 32'sd0.01797827343995584, 32'sd0.032117815786308464, 32'sd0.04658709469768601, 32'sd-0.03098671225762618, 32'sd0.0626830840043656, 32'sd0.11979505209647733, 32'sd0.12553086490551094, 32'sd0.1255140057959465, 32'sd0.0489264074838065, 32'sd0.12876096015546318, 32'sd-0.006274705349839343, 32'sd0.028909830392989642, 32'sd-0.011252097839501716, 32'sd-0.025656569567230163, 32'sd-0.054365231988735684, 32'sd0.05227311682298388, 32'sd-0.0032043169051490824, 32'sd0.12793102190159977, 32'sd4.8393046044020344e-122, 32'sd2.2482863984794592e-123, 32'sd4.872931821086446e-123, 32'sd1.4243774809423457e-127, 32'sd-5.164776782568633e-121, 32'sd-5.260962971127992e-118, 32'sd0.10748628874936901, 32'sd0.05807764353148555, 32'sd0.01943393438381365, 32'sd0.09121439274948576, 32'sd0.09736153926946728, 32'sd0.01315632716153677, 32'sd0.07118269946959378, 32'sd0.0037939440872066165, 32'sd0.09238886089608372, 32'sd0.005159616113091684, 32'sd0.08809642283296942, 32'sd0.12299651908645251, 32'sd-0.022970366088820613, 32'sd0.0469330678618431, 32'sd0.026972843108682854, 32'sd-0.044682892469849786, 32'sd0.0188030526435065, 32'sd0.027097439082047325, 32'sd-0.08202109399266248, 32'sd0.1222449561133931, 32'sd8.087508283717463e-117, 32'sd-6.654132773538568e-120, 32'sd1.5924266630449017e-115, 32'sd4.249912421670738e-125},
        '{32'sd1.679103554612049e-122, 32'sd1.9387155862467185e-120, 32'sd-1.088988069391741e-118, 32'sd7.08065730113402e-127, 32'sd-1.4296188296539605e-118, 32'sd-2.084693237977046e-128, 32'sd2.64108029254826e-124, 32'sd-1.4346950436378355e-118, 32'sd7.404489195174161e-120, 32'sd1.0647021987027437e-117, 32'sd-7.875527568185616e-117, 32'sd-2.8263221709097425e-126, 32'sd0.0018084505282746203, 32'sd-0.055495945335266146, 32'sd0.03156712652411143, 32'sd-0.006315945977649271, 32'sd3.222460416355522e-114, 32'sd-2.676167234659634e-117, 32'sd3.271192040238911e-122, 32'sd-3.1309433025359355e-123, 32'sd-1.2055412537723735e-122, 32'sd9.682676419836057e-121, 32'sd6.043795605648317e-127, 32'sd3.604098740228447e-116, 32'sd-6.09915550654937e-115, 32'sd1.0774552754029007e-119, 32'sd1.235175661237987e-125, 32'sd3.0626710525622758e-121, 32'sd-7.73452882753895e-117, 32'sd-1.340622925593797e-122, 32'sd-2.0712203521444858e-117, 32'sd-3.12245663043909e-120, 32'sd0.07705952752374866, 32'sd-0.040232422153815894, 32'sd-0.04137430165149633, 32'sd-0.0531362939949174, 32'sd0.02122567595323452, 32'sd0.02986649774786475, 32'sd0.05895794972290398, 32'sd0.09560784916072194, 32'sd-0.0365550731046457, 32'sd-0.04574909430124306, 32'sd-0.03377990965627075, 32'sd0.07729089513840111, 32'sd0.019409062970714087, 32'sd0.037412057722826776, 32'sd0.041503261950609764, 32'sd0.0658189845991113, 32'sd0.07026290548204227, 32'sd0.06488515227935622, 32'sd0.08253394649451767, 32'sd0.028758313203867663, 32'sd-1.0452806338262553e-123, 32'sd8.81967324800848e-119, 32'sd4.938065257649432e-124, 32'sd-9.99019725685656e-121, 32'sd-1.2325796456596674e-118, 32'sd-4.579874814766572e-124, 32'sd0.054837089921708077, 32'sd0.0716485081253038, 32'sd0.029537004068416563, 32'sd0.0028991736902473962, 32'sd-0.0008694225638920551, 32'sd0.0442637510696831, 32'sd0.05324898914059641, 32'sd-0.09814150883860172, 32'sd0.0022243961739290613, 32'sd-0.0013602648131398126, 32'sd-0.11041870653904301, 32'sd-0.0784008528974824, 32'sd-0.1015561307293145, 32'sd-0.21205865340995722, 32'sd-0.049050631768825195, 32'sd-0.11779346857926494, 32'sd-0.14364209795654487, 32'sd-0.022887776002718557, 32'sd0.0018875436037497, 32'sd-0.008159411704577449, 32'sd0.053133966919229315, 32'sd-0.028062688060464233, 32'sd0.022999080217472143, 32'sd0.06108552586501287, 32'sd-6.949782558223704e-124, 32'sd-1.928070335277952e-119, 32'sd-4.7441433744923385e-127, 32'sd-1.3967006091452853e-125, 32'sd-0.005936234678445113, 32'sd0.05998249788009811, 32'sd-0.046530868213689285, 32'sd-0.07169581659797429, 32'sd0.07528304283829525, 32'sd-0.04127709265780542, 32'sd-0.020835096190092557, 32'sd0.097940493771507, 32'sd-0.08958378314968365, 32'sd-0.051609614171390955, 32'sd-0.17887075215614498, 32'sd-0.12065725149508859, 32'sd-0.1342775885813238, 32'sd-0.0019299124177835905, 32'sd0.02096252859596846, 32'sd0.07052609542722897, 32'sd-0.01272782463769369, 32'sd-0.18113611666583243, 32'sd-0.08235663495670303, 32'sd-0.14097661364709102, 32'sd-0.01994930397124892, 32'sd0.009958555530342991, 32'sd-0.08368388951697985, 32'sd-0.10402417286772417, 32'sd0.029037429584621497, 32'sd-6.919328874144256e-124, 32'sd-1.6610615717444756e-121, 32'sd0.01934790547138846, 32'sd-0.016868697311230807, 32'sd0.051187135689517604, 32'sd0.014292313234400425, 32'sd0.03056262848168917, 32'sd0.020282699007402736, 32'sd-0.15689947362704135, 32'sd-0.168042434633448, 32'sd-0.13641989131391474, 32'sd-0.2702657168436457, 32'sd-0.15667881206032813, 32'sd-0.22194008918973918, 32'sd-0.1156370227048014, 32'sd0.02300413944938964, 32'sd0.014161561517031278, 32'sd0.06275372593810814, 32'sd-0.031052614260268514, 32'sd-0.0173412617910138, 32'sd-0.02504614955216305, 32'sd-0.10968939835859301, 32'sd0.011241070644103547, 32'sd-0.02792960881481411, 32'sd-0.00569429374673587, 32'sd-0.06862065550784575, 32'sd-0.048519770326104224, 32'sd-0.09678668975634641, 32'sd0.03545986577771526, 32'sd6.91459503204119e-124, 32'sd0.05609736936462048, 32'sd0.08065319045847232, 32'sd-0.0541069915667801, 32'sd-0.0886977059248288, 32'sd-0.092830195177925, 32'sd0.03026465059185103, 32'sd-0.10476994194790182, 32'sd-0.07871975269592192, 32'sd0.07734367732776007, 32'sd-0.03829355388980076, 32'sd-0.09846638140829402, 32'sd-0.15294951166414875, 32'sd0.008849458438555386, 32'sd0.03730612883064899, 32'sd-0.0085473971861181, 32'sd-3.8481903000882415e-05, 32'sd-0.07121389934951378, 32'sd-0.1438286234262688, 32'sd-0.2593085444138052, 32'sd-0.15400566348018302, 32'sd-0.0012679300547403544, 32'sd0.03977684977869776, 32'sd-0.15819329366712528, 32'sd-0.006835391694379629, 32'sd-0.1043343183561705, 32'sd0.10685762726897186, 32'sd0.003038364119701372, 32'sd-2.321101390910213e-116, 32'sd0.05250103501274471, 32'sd-0.020129316179630423, 32'sd0.028493262725649237, 32'sd-0.034937852055648665, 32'sd0.041545201182691865, 32'sd0.009827658830002826, 32'sd-0.05262196518717186, 32'sd-0.13757515789484726, 32'sd-0.07025066482280365, 32'sd-0.012321622545317186, 32'sd-0.1364179229302745, 32'sd-0.030293034407124875, 32'sd-0.06348162107532238, 32'sd0.03241070259762285, 32'sd0.023447714019321577, 32'sd-0.06808930303132808, 32'sd-0.07382053761593527, 32'sd-0.11618405299644496, 32'sd-0.06654055847783842, 32'sd-0.06432883824023193, 32'sd0.014538412823415182, 32'sd0.02859280361099125, 32'sd-0.03179797719549465, 32'sd-0.056423103673030175, 32'sd0.0046158383501446534, 32'sd0.06977322966930084, 32'sd-0.004782709333502212, 32'sd0.029120542380256933, 32'sd0.003748517920635135, 32'sd-0.06562456407422021, 32'sd-0.07012149223146029, 32'sd-0.02702688475213973, 32'sd-0.0776079854332855, 32'sd0.05469084212650349, 32'sd-0.17120731287875893, 32'sd-0.05176414280270922, 32'sd0.14776371426348386, 32'sd-0.0739378986166986, 32'sd-0.08330359920878914, 32'sd-0.1813864627551723, 32'sd-0.1156045213696589, 32'sd-0.03598460174653022, 32'sd0.05698677348411377, 32'sd-0.07154122595245237, 32'sd-0.07080259602559297, 32'sd-0.02632939096966957, 32'sd-0.0639644645382115, 32'sd-0.044790694709201696, 32'sd0.013927982214616707, 32'sd0.04878668016556015, 32'sd0.026408999151615434, 32'sd-0.010981888532193923, 32'sd0.05080396644104253, 32'sd0.09451436543720709, 32'sd0.10052675512315709, 32'sd0.008563599776007017, 32'sd0.04999369177540891, 32'sd0.04971906581887941, 32'sd-0.04703650561791929, 32'sd0.012058875819926122, 32'sd0.030308596019198823, 32'sd0.09795656286760798, 32'sd-0.10361624333401026, 32'sd-0.06742780321902432, 32'sd0.03474031849982184, 32'sd-0.06956940615514622, 32'sd-0.09603146458559124, 32'sd-0.015895616351504216, 32'sd0.04171157233389845, 32'sd0.10217436268349026, 32'sd0.03414762681299967, 32'sd0.06442902486804997, 32'sd-0.07600580440688495, 32'sd0.06748969055141239, 32'sd0.012929392435003875, 32'sd0.023287571318275434, 32'sd0.014240668983613805, 32'sd0.08686688878077395, 32'sd0.02626021823551123, 32'sd0.09761462586938521, 32'sd0.04954089172087649, 32'sd0.09724373895352939, 32'sd-0.04220731043803409, 32'sd0.011377809065310593, 32'sd-0.015120392240222307, 32'sd-0.031110426822129396, 32'sd0.10565008551818768, 32'sd-0.04713786017536056, 32'sd-0.05178327594505175, 32'sd0.05162469686813865, 32'sd0.09153313032310885, 32'sd-0.0064900582659082155, 32'sd-0.07927119962819362, 32'sd0.0027768046198191677, 32'sd0.04973139343564736, 32'sd0.007935032549378376, 32'sd-0.04805028380456843, 32'sd0.09295603008866889, 32'sd0.07607752909088313, 32'sd0.09369328442999679, 32'sd-0.14185777753310955, 32'sd-0.05215624565321686, 32'sd0.11131281846293994, 32'sd0.08226452073667569, 32'sd0.018219706288040052, 32'sd-0.05218434606344292, 32'sd0.07601730292274483, 32'sd0.1616943451997714, 32'sd-0.011682189843673734, 32'sd0.11410949940712833, 32'sd-0.008784172036703147, 32'sd0.013761223242873377, 32'sd0.03811917024348422, 32'sd0.004530642063680245, 32'sd0.15599374304911837, 32'sd0.11022313959129737, 32'sd-0.009761896334918077, 32'sd0.06167484697022872, 32'sd0.10152230746037251, 32'sd0.07750442085523715, 32'sd0.10995986692338629, 32'sd0.09043897823478748, 32'sd-0.0384211913496526, 32'sd0.11811731086636922, 32'sd-0.0303048264831079, 32'sd0.0692632022720434, 32'sd0.038043692939976545, 32'sd0.004072319722335857, 32'sd0.08336097716044184, 32'sd-0.01761248604372774, 32'sd-0.002366741730214472, 32'sd0.09638222489686436, 32'sd0.06826600946567943, 32'sd-0.011615746965098962, 32'sd0.06072812654827135, 32'sd0.020837729158798706, 32'sd0.09875237440135597, 32'sd-0.03544127424212441, 32'sd0.05004278447898257, 32'sd0.002572160707801904, 32'sd0.13259905922911452, 32'sd0.06967081848049317, 32'sd-0.06250553503164581, 32'sd-0.05124317415179917, 32'sd0.10440706897314593, 32'sd-0.007727538611061083, 32'sd0.007460858692164852, 32'sd0.019621677271989397, 32'sd0.1394932855554319, 32'sd0.1831854227827366, 32'sd0.13542982388993305, 32'sd0.08950040825174363, 32'sd-0.0666453765870562, 32'sd-0.03934414557044167, 32'sd0.09369580265507033, 32'sd0.10895501187463397, 32'sd0.08561053786802363, 32'sd-0.10088337757896847, 32'sd-0.055298965175335016, 32'sd-0.008981095052533274, 32'sd-0.0033369203501407993, 32'sd-0.09509958780956955, 32'sd0.021125549365813543, 32'sd0.006930353678397203, 32'sd-0.022157924961080714, 32'sd-0.09210837779795467, 32'sd-0.06868389513732484, 32'sd0.04056596700191495, 32'sd0.026416268331653097, 32'sd-0.0029739096340133326, 32'sd0.019417810726597186, 32'sd-0.23174624952495032, 32'sd-0.15636185126989363, 32'sd0.0431688006921372, 32'sd-0.007079688867204441, 32'sd-0.07771007398711283, 32'sd0.13874137359888222, 32'sd0.03657162426435303, 32'sd0.03817918422567778, 32'sd0.08940433076066591, 32'sd0.09552113320887698, 32'sd-0.01923069153189808, 32'sd0.04220455481818102, 32'sd0.0698646470946141, 32'sd0.009128054550076788, 32'sd0.022772380452085905, 32'sd-0.06186640507928285, 32'sd0.02521125469718223, 32'sd-0.005928984779891153, 32'sd-0.07052537892146582, 32'sd0.03036369995699308, 32'sd0.06051116963732743, 32'sd-0.06479402694558588, 32'sd-0.012801631325579856, 32'sd-0.02126464677513789, 32'sd0.033381977168360964, 32'sd0.038830156493978064, 32'sd0.04332655078987708, 32'sd-0.006507593361204605, 32'sd-0.22552803081419429, 32'sd-0.011804632638961279, 32'sd-0.08828915585951362, 32'sd-0.07682887465293393, 32'sd0.06029089008211582, 32'sd0.11715764371791607, 32'sd0.008171624452304958, 32'sd0.14687998789249837, 32'sd0.10864860700306465, 32'sd-0.04198237036518814, 32'sd-0.06468406987444113, 32'sd0.053501058664278504, 32'sd0.008145001177536226, 32'sd-0.004093929900834436, 32'sd-0.08718048083010327, 32'sd-0.029991563541583825, 32'sd-0.024796587403339756, 32'sd-0.045695991366987966, 32'sd-0.033905812518197014, 32'sd0.025623858900339122, 32'sd-0.014639466544924245, 32'sd-0.03374663526100109, 32'sd-0.13011133706269742, 32'sd0.010846511726508875, 32'sd0.1101913994474591, 32'sd-0.04405611250789623, 32'sd-0.0050309792094932445, 32'sd-0.08111445934908802, 32'sd-0.09815560853835412, 32'sd0.03365299151447824, 32'sd0.054264458383314555, 32'sd0.11306072251889818, 32'sd0.03989185548067938, 32'sd0.0904522148307164, 32'sd0.1326472278005169, 32'sd0.16536501048229174, 32'sd0.07827539095739047, 32'sd0.03328014781088277, 32'sd-0.022978530447769818, 32'sd-0.09079515663243969, 32'sd-0.06247524556757196, 32'sd0.029407309241574867, 32'sd-0.0382631591251788, 32'sd0.05341696652585449, 32'sd-0.11463110986957972, 32'sd-0.07578295887528698, 32'sd0.051092540294069316, 32'sd0.03001376968915715, 32'sd0.10044250614380021, 32'sd-0.19142526740927032, 32'sd-0.08925481985164477, 32'sd-0.06485368311319874, 32'sd0.08259157134113897, 32'sd-0.06711447284357203, 32'sd-0.05341242722301936, 32'sd-0.00841969481134201, 32'sd-0.020442267476025486, 32'sd0.04947758435058268, 32'sd0.01694977758377779, 32'sd0.2175651228422755, 32'sd0.07209423179442488, 32'sd0.07715494714636667, 32'sd0.0923220727257659, 32'sd0.042055611622989236, 32'sd0.12750163491352476, 32'sd-0.16540792796350431, 32'sd-0.09385188252338424, 32'sd-0.034854681385595325, 32'sd0.015519420108974077, 32'sd-0.10335846888205394, 32'sd-0.02894757810561763, 32'sd-0.02047174618785666, 32'sd-0.08162877141444687, 32'sd-0.035529654311806255, 32'sd-0.022469122804814917, 32'sd0.12888306464753624, 32'sd0.22599320166486786, 32'sd-0.07632106312703615, 32'sd-0.10349141956331598, 32'sd0.008430027352270603, 32'sd0.016226055912727116, 32'sd0.004874811433760195, 32'sd-0.008461233398736105, 32'sd-0.05701958317372746, 32'sd-0.061903193234012215, 32'sd0.03159896952601904, 32'sd0.12870472354058912, 32'sd0.06415666235770456, 32'sd0.27663999489029767, 32'sd0.13828606704084145, 32'sd0.16962172533734196, 32'sd-0.010637864983418033, 32'sd-0.03696032234645483, 32'sd-0.1595245189665204, 32'sd-0.2146322125547067, 32'sd-0.04185774580122729, 32'sd-0.09592670928613523, 32'sd-0.03345694330434178, 32'sd-0.037666192806002495, 32'sd0.09038487229598818, 32'sd0.00826879355515606, 32'sd0.015460793835491381, 32'sd0.020497963476470437, 32'sd0.12715825271969358, 32'sd0.18014527034438516, 32'sd-0.06635096657728523, 32'sd-0.21501000604214693, 32'sd0.08185215035283114, 32'sd-1.8116594781817277e-123, 32'sd0.03210238016776825, 32'sd-0.011823651528201064, 32'sd-0.06297890989302649, 32'sd0.0235673260676156, 32'sd0.09133317884279706, 32'sd0.08456162715707123, 32'sd-0.052704103350471564, 32'sd0.16730102783882397, 32'sd0.18283405181871468, 32'sd0.13227671124786744, 32'sd0.06849779280977134, 32'sd-0.11880585318750857, 32'sd-0.11421321674094156, 32'sd-0.1275386741223048, 32'sd-0.0024360102621045388, 32'sd0.0857407134066217, 32'sd0.07272553677366153, 32'sd0.0103078369635441, 32'sd-0.007292605149448948, 32'sd0.1337542881726457, 32'sd0.08786227712043354, 32'sd0.05559164457888296, 32'sd0.07868628806880962, 32'sd0.004199962649761448, 32'sd-0.011351050007074922, 32'sd-0.056803194847574234, 32'sd-0.03159785000944424, 32'sd-0.04982329518748621, 32'sd0.0022085060609536708, 32'sd0.055528943000204445, 32'sd-0.02998618750072555, 32'sd0.131359012984804, 32'sd0.042853279020633545, 32'sd-0.07626092849045663, 32'sd0.005808528467260534, 32'sd0.19889061359461432, 32'sd0.1764070682195688, 32'sd0.04717842041099859, 32'sd-0.10581117728363873, 32'sd-0.06148259458244291, 32'sd-0.08199062272064842, 32'sd0.028590450734367303, 32'sd-0.05008607325648629, 32'sd0.05061780486709105, 32'sd-0.03628119965563122, 32'sd-0.07727213260501742, 32'sd-0.09290615476726584, 32'sd0.11391433960385362, 32'sd0.0005162469896261586, 32'sd-0.07692098463467377, 32'sd-0.052101266865766556, 32'sd0.0656354123600789, 32'sd0.05532554352105606, 32'sd-0.07045010228370317, 32'sd0.05365375846277347, 32'sd0.046036775042999564, 32'sd0.0184528218279484, 32'sd-0.055669748933028916, 32'sd0.06817888470952072, 32'sd0.015954742738785662, 32'sd0.015170955759588812, 32'sd-0.043633760987009725, 32'sd-0.10633919826457727, 32'sd0.16901902411999167, 32'sd0.15832296753950972, 32'sd0.054935782737237364, 32'sd-0.20785738842703477, 32'sd-0.153892397039393, 32'sd-0.045319077103152416, 32'sd-0.04061101379637715, 32'sd-0.11407559809242918, 32'sd0.03455972312265711, 32'sd-0.022146756578480968, 32'sd-0.07746461664019179, 32'sd-0.09371403397548123, 32'sd-0.032699760620814915, 32'sd-0.0785802103505115, 32'sd-0.204129201435035, 32'sd-0.08991287513536494, 32'sd0.11222252416027241, 32'sd-0.004078539584520687, 32'sd-0.08588691124931504, 32'sd0.08301212647207787, 32'sd-2.1175722355052784e-117, 32'sd0.01348090181141749, 32'sd-0.053755565117393364, 32'sd0.011803275165113526, 32'sd0.006574787588349301, 32'sd-0.025015015067864566, 32'sd0.014173429178981492, 32'sd-0.10973486175474645, 32'sd-0.008117187415215055, 32'sd-0.028108976306176765, 32'sd-0.07487190551235459, 32'sd0.02820873829674107, 32'sd-0.0699615445472816, 32'sd-0.07520894468611831, 32'sd-0.07417270829813183, 32'sd-0.07127613363995973, 32'sd-0.07795302014352683, 32'sd-0.010577102097004512, 32'sd-0.12321819884363737, 32'sd-0.06279385411103948, 32'sd-0.030052481588404033, 32'sd-0.18012376232917907, 32'sd-0.17390848102788872, 32'sd-0.0890094719611749, 32'sd-0.09961546780275038, 32'sd0.025317791447146985, 32'sd-0.06987328766833427, 32'sd0.032419892519218445, 32'sd0.046493855385624394, 32'sd0.09742609426958769, 32'sd-0.09761556785567321, 32'sd0.111321621699792, 32'sd-0.038522884753900054, 32'sd0.04459588633019092, 32'sd-0.057961321919855834, 32'sd-0.05244905845943038, 32'sd-0.011521557035566373, 32'sd-0.002719276751479659, 32'sd0.022536468239119353, 32'sd0.014441103350657883, 32'sd-0.1541303513926204, 32'sd-0.18798169976892365, 32'sd-0.22459360527204944, 32'sd-0.06408353258496488, 32'sd-0.016285957471720798, 32'sd-0.06519800246697416, 32'sd-0.10025605300755508, 32'sd-0.01704329431391046, 32'sd0.01446731760522356, 32'sd0.05334927058207228, 32'sd-0.032730539178684986, 32'sd-0.08246369203315372, 32'sd-0.11285441313323466, 32'sd-0.09728087683559988, 32'sd0.031594759072204055, 32'sd0.0047627599248302455, 32'sd0.048572250549302, 32'sd0.06645227329759908, 32'sd0.025694543194796325, 32'sd-0.047291828703362515, 32'sd-0.13287683590974064, 32'sd-0.011913102157145646, 32'sd0.015422247310738026, 32'sd0.06418442281176567, 32'sd0.03606147185208659, 32'sd0.05670968654809658, 32'sd0.023695234247713495, 32'sd-0.005130248404998731, 32'sd-0.009130671345117554, 32'sd-0.07032820530950909, 32'sd-0.024890113884070652, 32'sd-0.06186986198029583, 32'sd0.04381563706719255, 32'sd-0.08230422086860814, 32'sd-0.11838086906820935, 32'sd-0.06152437439751385, 32'sd0.015588504217896712, 32'sd0.02772786994878826, 32'sd-0.01744594195523837, 32'sd-0.03557140467972594, 32'sd-0.02414675020943972, 32'sd-0.12443011635629254, 32'sd0.018143092658964327, 32'sd0.036112738793550564, 32'sd-9.624063118149198e-121, 32'sd0.022488793743007975, 32'sd-0.007763482172783596, 32'sd-0.0777423749713994, 32'sd-0.05627142535761077, 32'sd0.05004850977033824, 32'sd0.03871456621108416, 32'sd-0.05799819839161557, 32'sd-0.013588620707885846, 32'sd-0.03813559452471733, 32'sd0.08976539960930943, 32'sd-0.05555848225335707, 32'sd-0.0032291929195654976, 32'sd-0.11806508658994655, 32'sd-0.07317708198323071, 32'sd0.042431414464046975, 32'sd-0.023549837739779683, 32'sd-0.08258903715529192, 32'sd-0.06782688832492838, 32'sd0.04410244154673811, 32'sd0.07012665521383797, 32'sd0.020397592670382117, 32'sd-0.007901232336156605, 32'sd-0.06392126633075762, 32'sd-0.0020953023226504214, 32'sd-0.05822887657501547, 32'sd0.02402706727600885, 32'sd3.0097777365750253e-122, 32'sd-3.820472006654242e-123, 32'sd-9.528902188708359e-124, 32'sd-0.02064193691622989, 32'sd0.013362145061107238, 32'sd0.07429575286798287, 32'sd0.03818370722727321, 32'sd-0.0819254950489536, 32'sd-0.048941468010996914, 32'sd0.05475513445466009, 32'sd0.08869922525141886, 32'sd0.06729462631359195, 32'sd0.008783526677320333, 32'sd-0.016372135450823586, 32'sd0.07599560734382334, 32'sd0.010494292892658491, 32'sd-0.08729323763622228, 32'sd-0.009162467197387511, 32'sd-0.08963281947937146, 32'sd0.0511262921375549, 32'sd0.04931240345788632, 32'sd-0.04253105427558694, 32'sd0.021506793001736288, 32'sd-0.06738446166643194, 32'sd-0.05950202213759923, 32'sd0.01123561983936034, 32'sd0.0828442879391402, 32'sd0.0044087972586080715, 32'sd-2.563901247380707e-126, 32'sd-2.006078764975972e-125, 32'sd2.716332955423176e-124, 32'sd0.042839446482172375, 32'sd-0.06031877367436212, 32'sd-0.07489496579952722, 32'sd-0.03113052277665014, 32'sd-0.10620474522975223, 32'sd-0.060268056793545334, 32'sd-0.03215983870648926, 32'sd0.10617674596806918, 32'sd-0.1631945410596838, 32'sd-0.023422614601501274, 32'sd0.02456469860055593, 32'sd-0.11431540460410697, 32'sd-0.05634707675090886, 32'sd-0.02669964642548583, 32'sd-0.13948916462574149, 32'sd-0.11655428158496695, 32'sd-0.020706349549525882, 32'sd-0.07778622050296516, 32'sd0.02739292322861656, 32'sd-0.010944101182349876, 32'sd-0.13531816070012523, 32'sd0.042973471494077334, 32'sd0.06669123548954285, 32'sd0.030057931892448226, 32'sd0.01631002054003941, 32'sd-1.2178068655245353e-117, 32'sd5.714270052993387e-119, 32'sd-6.127823134508667e-123, 32'sd-1.8624624267465176e-126, 32'sd0.06405712709416309, 32'sd0.005679933091460895, 32'sd-0.07154270216683978, 32'sd-0.1066795693171376, 32'sd-0.06888338630469423, 32'sd-0.15121099949357128, 32'sd-0.07011161499223886, 32'sd-0.025647576032430956, 32'sd-0.05446381298428578, 32'sd0.05392439774834029, 32'sd-0.06323291204529384, 32'sd-0.17181479067628755, 32'sd-0.14717235587271793, 32'sd0.013002009483370333, 32'sd0.007859876456452653, 32'sd-0.014056605699106684, 32'sd0.016261685838119655, 32'sd-0.0890639907723567, 32'sd-0.13396753475684953, 32'sd-0.02526583952323165, 32'sd-0.06227219336627438, 32'sd-0.010993403211205694, 32'sd0.020690048060320113, 32'sd2.438684056798753e-126, 32'sd3.713616061426933e-119, 32'sd1.9222389780809137e-121, 32'sd-1.3466657211721902e-115, 32'sd-1.1838449968600525e-118, 32'sd-4.410136745617717e-118, 32'sd0.07957016178487561, 32'sd0.0045811142117297395, 32'sd0.0034520570282975576, 32'sd0.08050056081969345, 32'sd-0.0006148794973075771, 32'sd-0.0027800222235620934, 32'sd-0.005399817580856012, 32'sd-0.07083681627046128, 32'sd0.06541516685660145, 32'sd0.029134881064499477, 32'sd-0.14483787594588002, 32'sd-0.14359934127786983, 32'sd-0.1356654783547619, 32'sd-0.02419712493273974, 32'sd0.0008553252475608618, 32'sd-0.01747479486012697, 32'sd-0.03740662275541935, 32'sd0.045973883486819925, 32'sd-0.00873385970605731, 32'sd0.00689409550968206, 32'sd-2.8435688727509226e-114, 32'sd-1.0225436510517852e-125, 32'sd-1.602611136676213e-117, 32'sd2.7753299352203527e-116},
        '{32'sd2.101206486560551e-117, 32'sd4.789117211304697e-118, 32'sd-6.758060023823991e-116, 32'sd4.312497340099715e-123, 32'sd3.8294527533566234e-125, 32'sd-3.365327600286977e-129, 32'sd5.256827415906486e-118, 32'sd1.2731140202196474e-117, 32'sd-4.688919478318981e-118, 32'sd-1.6896931887392358e-125, 32'sd-2.625438218318968e-121, 32'sd-9.591555032876726e-120, 32'sd0.14852843617181405, 32'sd0.15077259532433784, 32'sd-0.015259283631157007, 32'sd0.04139333239211169, 32'sd-3.503000073328145e-125, 32'sd9.117342111776273e-122, 32'sd-9.841794835958599e-125, 32'sd-3.274727452997635e-116, 32'sd-3.6274082442997486e-114, 32'sd-2.307750098066753e-126, 32'sd5.3336965037828214e-120, 32'sd3.0934060217546564e-115, 32'sd1.0484300225041393e-120, 32'sd-8.426825398441683e-127, 32'sd-4.858147911059069e-118, 32'sd4.187012792961671e-123, 32'sd5.240630126716073e-124, 32'sd1.1573311374988909e-118, 32'sd-6.152801829274975e-115, 32'sd5.95431088781888e-126, 32'sd0.12681536876742036, 32'sd0.02330087319774689, 32'sd0.01084233683689723, 32'sd0.052510162265906914, 32'sd-0.0032316887280630213, 32'sd0.09763622753618474, 32'sd0.07111305683247345, 32'sd-0.050250977216346915, 32'sd-0.005255181662302824, 32'sd0.17249918094041314, 32'sd0.001789981935932698, 32'sd0.1327566904158442, 32'sd0.04418215673661923, 32'sd0.06925552705148325, 32'sd-0.02692052692917511, 32'sd0.06482849274767137, 32'sd0.06318835741398617, 32'sd0.03316352435483473, 32'sd-0.03971614122704263, 32'sd0.04234792633076378, 32'sd1.9254033275337708e-121, 32'sd-3.1502208064086858e-115, 32'sd4.119733087172126e-124, 32'sd3.2644836824393225e-117, 32'sd1.3559417097826242e-123, 32'sd-1.664654271334775e-120, 32'sd0.05186193280906339, 32'sd0.09710934637856042, 32'sd0.05426624702131894, 32'sd-0.04550657903682166, 32'sd-0.08019444978171295, 32'sd0.04262274421908919, 32'sd0.14704143144165974, 32'sd0.14666382177287762, 32'sd0.016027367521005448, 32'sd0.14510245815696673, 32'sd0.08921238481344479, 32'sd-0.02915773747115666, 32'sd0.05341626709310876, 32'sd0.1329438599500621, 32'sd0.029532631962193894, 32'sd0.09935444193248853, 32'sd0.07541776578521014, 32'sd-0.06718263398502652, 32'sd0.003244127655775083, 32'sd0.049979130302699695, 32'sd-0.09561820925054727, 32'sd-0.08946977795930068, 32'sd0.0386322279954148, 32'sd0.13101580739751573, 32'sd-2.1083923461739608e-127, 32'sd-1.96177661157992e-126, 32'sd1.0412526891767114e-120, 32'sd-4.855706006893419e-126, 32'sd0.013392515496905833, 32'sd0.024634181736943095, 32'sd0.004821990227984172, 32'sd0.06138009949030692, 32'sd-0.012626092089881826, 32'sd0.10955170414884349, 32'sd0.14445337998365088, 32'sd0.1202531695865853, 32'sd-0.058147682034630395, 32'sd0.13280993301530866, 32'sd0.052764269440305954, 32'sd0.14116755249476276, 32'sd0.065421037156224, 32'sd0.09939904632409781, 32'sd0.04284941389299484, 32'sd-0.08736330154857101, 32'sd0.02856595907768642, 32'sd0.10176201185411542, 32'sd0.0327437424471632, 32'sd0.05606196359629213, 32'sd-0.005628774640740424, 32'sd0.02944420931084255, 32'sd0.03503775346832174, 32'sd-0.008600061362962548, 32'sd0.1116030060665412, 32'sd3.053004034255054e-118, 32'sd-2.1660805761323665e-121, 32'sd0.030893910886504374, 32'sd0.04395689288009255, 32'sd0.02799580027640078, 32'sd0.0677703792512714, 32'sd-0.022624199492396333, 32'sd-0.020934565742641752, 32'sd0.02783843545655794, 32'sd0.10587461557682432, 32'sd0.07282724687542047, 32'sd-0.017569662746508695, 32'sd0.002584754969231551, 32'sd0.17065100702129873, 32'sd0.1673100456991864, 32'sd0.05419421373999608, 32'sd0.1140766522740742, 32'sd-0.10790213612663392, 32'sd-0.043272357849925065, 32'sd-0.07928789316219521, 32'sd-0.09929121221154241, 32'sd-0.0352470337181902, 32'sd-0.004278551638485007, 32'sd-0.1093422265894004, 32'sd0.014302445074878083, 32'sd-0.0020055970932729927, 32'sd0.05195079175413463, 32'sd0.029206262653286144, 32'sd0.0880804458904091, 32'sd6.435026228999371e-120, 32'sd0.07688081052950764, 32'sd0.050487751966975185, 32'sd0.039524160264413986, 32'sd-0.005735874347055711, 32'sd-0.042330422964822735, 32'sd0.1385030883135108, 32'sd-0.01211329214892465, 32'sd-0.019236029905936914, 32'sd-0.14903667175112306, 32'sd-0.14240145288597544, 32'sd-0.03982145601120044, 32'sd0.05273979302548754, 32'sd0.02173273993077837, 32'sd0.016905825237247974, 32'sd0.0667544836563833, 32'sd-0.06683534483077236, 32'sd-0.018740506777350344, 32'sd-0.0973776559310337, 32'sd-0.032002628448330794, 32'sd-0.06220563474488412, 32'sd-0.03977005747861998, 32'sd-0.10451141371390389, 32'sd-0.09566277233780249, 32'sd-0.023888260231737565, 32'sd0.005462398146737902, 32'sd0.05895010984880936, 32'sd0.017965966605424377, 32'sd1.6953468339251386e-127, 32'sd0.041508359973510815, 32'sd0.029467071925128478, 32'sd-0.05049160314415474, 32'sd-0.11307918523973223, 32'sd-0.09605452902100846, 32'sd-0.020672400652903867, 32'sd0.016940348480895404, 32'sd-0.02321066243787102, 32'sd-0.041502190460268776, 32'sd0.0017484480391172761, 32'sd0.015636762302757862, 32'sd0.076734189484888, 32'sd0.12613054184413566, 32'sd0.1198625294306266, 32'sd0.06488161083023913, 32'sd-0.0840282957598454, 32'sd-0.05504397614515326, 32'sd-0.11129691327036177, 32'sd-0.12084844034418692, 32'sd-0.1724843552334367, 32'sd-0.039084023117741375, 32'sd-0.20157255140906327, 32'sd-0.07923362873674494, 32'sd0.007476842576686959, 32'sd-0.009709592742754692, 32'sd0.13204885966128316, 32'sd-0.049189794084740085, 32'sd0.03896858976211215, 32'sd-0.029637702870903636, 32'sd0.0036202995942755723, 32'sd-0.021196052425306172, 32'sd-0.06524019167765081, 32'sd-0.1289877224173805, 32'sd-0.1390866942049938, 32'sd0.049893807499486006, 32'sd0.05760353035323465, 32'sd-0.0898068243295931, 32'sd-0.022638810150822416, 32'sd0.12477645150519276, 32'sd0.1376557970474785, 32'sd0.20281459103397162, 32'sd0.10044229919475034, 32'sd0.06878881499035172, 32'sd-0.13629473079418403, 32'sd-0.23467628349293362, 32'sd-0.03018745809431426, 32'sd-0.15244886662090318, 32'sd-0.1437597261912378, 32'sd-0.19485769474112016, 32'sd0.010215657118502868, 32'sd-0.06709746166650447, 32'sd0.027607164246821695, 32'sd0.09949191970335543, 32'sd0.01913941462891986, 32'sd0.0559743937341681, 32'sd0.031331906278890306, 32'sd0.0722994629857483, 32'sd0.031841113320639686, 32'sd-0.1120348814323663, 32'sd-0.03899051832517517, 32'sd-0.05682569891995094, 32'sd-0.06624947036540228, 32'sd-0.03370965332881899, 32'sd-0.018944512051853792, 32'sd-0.005158092366118319, 32'sd0.106031811600053, 32'sd0.034250366837282595, 32'sd0.0018720700297413632, 32'sd0.17440159820703532, 32'sd0.002562108517598048, 32'sd-0.13968498314909777, 32'sd-0.18955479276430307, 32'sd-0.03913361983623778, 32'sd-0.01915479127012868, 32'sd-0.13278442517972652, 32'sd-0.12260292529952865, 32'sd-0.12498120762574501, 32'sd-0.05265893254434955, 32'sd-0.15024134993116706, 32'sd-0.07818070325802454, 32'sd0.07270599096676708, 32'sd0.12467896231786363, 32'sd0.016482330210496384, 32'sd0.0006825482411135164, 32'sd0.05127118896159893, 32'sd0.05971947285236655, 32'sd0.06300891472323403, 32'sd0.004760517894912725, 32'sd0.01041286627683818, 32'sd-0.023887399689576174, 32'sd0.10884382285101649, 32'sd0.0607245771148686, 32'sd0.13255220393953723, 32'sd-0.0008007619806899825, 32'sd0.0398472088195576, 32'sd-0.07933644158019076, 32'sd0.04805054301560351, 32'sd0.014857574384317252, 32'sd-0.11776283842710705, 32'sd-0.03587730321796778, 32'sd0.0230877404251285, 32'sd0.02917672619001618, 32'sd0.02713605464267636, 32'sd-0.029196950519872106, 32'sd-0.06582537430804403, 32'sd-0.001242590555320644, 32'sd-0.030837908968625042, 32'sd0.07831675304426254, 32'sd0.015183065191136403, 32'sd0.08787249745774135, 32'sd-0.022301713427292084, 32'sd-0.041030377356539936, 32'sd-0.01971587382353225, 32'sd0.008330848048442837, 32'sd-0.04565054566617397, 32'sd0.07549177227486335, 32'sd-0.023744936840962835, 32'sd0.02379636521667283, 32'sd0.03623773875164638, 32'sd-0.015244189870683109, 32'sd-0.10228528095138041, 32'sd-0.0052225422366425425, 32'sd-0.02808392943246919, 32'sd-0.019193606552401668, 32'sd0.07724955520162552, 32'sd-0.04600432421556688, 32'sd-0.1500904999105454, 32'sd0.02000084141208851, 32'sd0.047725442040629215, 32'sd-0.01951559820429506, 32'sd0.038226125625512516, 32'sd-0.037946583197579806, 32'sd-0.10000714532233682, 32'sd0.06258251962594812, 32'sd0.006924637028066405, 32'sd-0.10197860858036352, 32'sd0.03233734595683279, 32'sd0.12336123490630789, 32'sd0.02804397166141274, 32'sd0.07424880746362514, 32'sd-0.019971804756608216, 32'sd-0.00023951243521807175, 32'sd0.07448633779875874, 32'sd-0.022391711307809942, 32'sd0.023050444759376384, 32'sd0.02875842900214418, 32'sd0.025751582748989827, 32'sd-0.012383037480953972, 32'sd-0.017716225612583823, 32'sd-0.03659929645182083, 32'sd0.022247701385835005, 32'sd-0.04309179581331059, 32'sd0.08086576501860576, 32'sd0.04831555010186818, 32'sd-0.11435842296940231, 32'sd0.02673846604093009, 32'sd0.002084219430373578, 32'sd0.07755104415593911, 32'sd0.11675833979773594, 32'sd0.0911876612161964, 32'sd-0.0025932187159860808, 32'sd-0.05105079552521275, 32'sd-0.1065611880273726, 32'sd-0.05276432970146724, 32'sd0.04529574687159283, 32'sd0.047654831462729585, 32'sd0.05724663303599996, 32'sd0.0229373292466096, 32'sd0.020255872004553553, 32'sd-0.009262366668842722, 32'sd-0.09973079201199175, 32'sd0.11329942565284427, 32'sd0.027312657328813515, 32'sd-0.011310801936797857, 32'sd0.0026296197313016244, 32'sd-0.05025115339008721, 32'sd-0.020720453588464624, 32'sd-0.08798615024442971, 32'sd-0.058068407106679154, 32'sd-0.10639246834343469, 32'sd-0.08599198585792618, 32'sd0.05750118464492757, 32'sd-0.0590831100368904, 32'sd0.0668611687041334, 32'sd0.09365584175894388, 32'sd0.1242825538024494, 32'sd0.12035051832191104, 32'sd0.05822302418859686, 32'sd0.008328743779254863, 32'sd-0.07801720251648125, 32'sd0.021320906713648172, 32'sd0.16475091769656638, 32'sd0.09350906635416918, 32'sd-0.08805530968470528, 32'sd-0.005643759960433722, 32'sd0.00852615162297784, 32'sd-0.01899097816533814, 32'sd0.04110051911685609, 32'sd-0.06997445770407038, 32'sd-0.07880307147939801, 32'sd-0.0023477611111594812, 32'sd0.010927492455998606, 32'sd-0.03628004086327629, 32'sd-0.07978359317206851, 32'sd-0.004919015620182479, 32'sd-0.015244670670228864, 32'sd-0.08858808885378627, 32'sd-0.17933496557799405, 32'sd-0.17068769587250415, 32'sd0.02223732713375971, 32'sd0.06953314982816397, 32'sd0.11458176770195877, 32'sd0.09224750070905759, 32'sd-0.021433215091729185, 32'sd0.07040196098393958, 32'sd-0.01030792889851962, 32'sd0.057503732394352663, 32'sd-0.043796064938467945, 32'sd0.028704492876182566, 32'sd0.057818475691841856, 32'sd-0.006386623853477528, 32'sd-0.00934249498180574, 32'sd0.04762308140681894, 32'sd0.01706554531244327, 32'sd-0.043597221382598306, 32'sd0.044270543874508, 32'sd-0.089566071735235, 32'sd-0.18982004649474146, 32'sd-0.023462290492918342, 32'sd-0.05983561459029367, 32'sd0.0684315675543566, 32'sd0.032424201538941363, 32'sd0.009103303849344987, 32'sd-0.09810366185957613, 32'sd-0.12068388974880224, 32'sd-0.08695193627749971, 32'sd-0.0740027663815509, 32'sd-0.020844278519280595, 32'sd0.09137433242319218, 32'sd0.12705391297812732, 32'sd0.010179836297085559, 32'sd-0.009972364855523918, 32'sd-0.114896606034246, 32'sd-0.04831030104712184, 32'sd-0.06704536742239679, 32'sd0.0908297894952467, 32'sd0.036866932935586724, 32'sd-0.03783505734221329, 32'sd-0.035416736212601115, 32'sd-0.005589386606417776, 32'sd0.08295774163147852, 32'sd0.020990503565678244, 32'sd0.0036257700861895277, 32'sd-0.032012516631991346, 32'sd-0.06435340810335938, 32'sd-0.11749160963527705, 32'sd-0.01790074929894699, 32'sd0.03799615540646966, 32'sd0.049859070277023965, 32'sd0.01717762895776871, 32'sd-0.11992102519419591, 32'sd-0.1446910542881802, 32'sd-0.025704922438228788, 32'sd-0.05646559200604956, 32'sd-0.029432646743803928, 32'sd0.13196304970930245, 32'sd0.07316967912072621, 32'sd0.019549377145002163, 32'sd0.017583541287251526, 32'sd0.028274569682034442, 32'sd-0.006319420347222892, 32'sd0.024720340717036417, 32'sd0.014211557890322843, 32'sd0.02367016687052582, 32'sd0.05464987696808762, 32'sd0.03580756284692774, 32'sd-0.0704433017503107, 32'sd0.05631219157700337, 32'sd0.012635695810840139, 32'sd0.03324851618414212, 32'sd0.03285012070861591, 32'sd0.030202025795205124, 32'sd-0.009267170188416229, 32'sd-0.02178770521092377, 32'sd-0.0514430613273127, 32'sd-0.07536143579621991, 32'sd0.03781110578728273, 32'sd-0.015410840624013288, 32'sd-0.15161391893890522, 32'sd-0.18802723519901207, 32'sd-0.06855799653183237, 32'sd-0.0646553845425421, 32'sd0.09505611857139576, 32'sd0.11437687825556796, 32'sd0.07535000713789808, 32'sd0.004736673469049109, 32'sd0.06972103653830496, 32'sd-0.05578939028764101, 32'sd-0.14342939017129572, 32'sd-0.020239470027484704, 32'sd-0.05218430730730116, 32'sd-0.024536059843326824, 32'sd-0.014416610945459468, 32'sd0.08032186064723958, 32'sd0.06318642569675123, 32'sd0.021589964271133116, 32'sd0.05308059657215529, 32'sd-3.4695157873302815e-118, 32'sd0.029024462539136764, 32'sd-0.05819003497089179, 32'sd0.06779325741349947, 32'sd0.10737565475260222, 32'sd-0.0022043228168564205, 32'sd-0.012517260609044208, 32'sd-0.05550553134308734, 32'sd-0.14044162277527356, 32'sd-0.15743602361988518, 32'sd-0.08968523584972966, 32'sd-0.005346181024117361, 32'sd-0.004340340090213254, 32'sd0.14945286625604076, 32'sd0.022044341268412967, 32'sd0.08640478095313964, 32'sd-0.060772591771758463, 32'sd-0.0052261069150519365, 32'sd-0.06363340297145388, 32'sd-0.011038153956741344, 32'sd-0.03498640301175902, 32'sd-0.013443181188085837, 32'sd0.003332078518500044, 32'sd0.10551750677464085, 32'sd0.07056382715008462, 32'sd0.13237370491796382, 32'sd0.05704679057416076, 32'sd-0.06785867613906364, 32'sd0.09385896438424286, 32'sd0.06360961778497211, 32'sd-0.02168106620221679, 32'sd-0.03792499707202695, 32'sd-0.00022956469159282148, 32'sd-0.09682326235736625, 32'sd0.0031795578671186576, 32'sd-0.07140988191413929, 32'sd-0.13214886078633992, 32'sd-0.10221514957772161, 32'sd-0.10721780784391582, 32'sd-0.06420690263557899, 32'sd0.07374157910355854, 32'sd0.03378613542878476, 32'sd0.04985428758676198, 32'sd0.08851538285321288, 32'sd-0.042400630779371416, 32'sd-0.018692519579851186, 32'sd0.026930354534828897, 32'sd-0.01658567361365616, 32'sd-0.08097846815165646, 32'sd-0.04225591375185946, 32'sd0.014424381765585314, 32'sd-0.10570395411537595, 32'sd0.10027227173596731, 32'sd0.11855954066362079, 32'sd-0.08913227935425552, 32'sd0.013113347888293964, 32'sd0.04214935877011004, 32'sd0.06392096403300904, 32'sd-0.03108537290841278, 32'sd-0.16969288111219105, 32'sd0.09342081775082199, 32'sd-0.03843767472701477, 32'sd-0.039582943995317345, 32'sd0.00743576438970124, 32'sd-0.00027807795355346877, 32'sd-0.07580886888963535, 32'sd-0.007169048008430899, 32'sd-0.004949478116397902, 32'sd0.1293219927469107, 32'sd-0.10031259611946379, 32'sd-0.0020993967690785932, 32'sd0.0072070478908766505, 32'sd0.03426722911291882, 32'sd0.032354866508430453, 32'sd0.019636104800837783, 32'sd-0.0025211108390706134, 32'sd0.07732673062125599, 32'sd0.08587927537510263, 32'sd-0.07424500438826152, 32'sd-0.08932453382071236, 32'sd0.0026663331203669624, 32'sd-0.01126871036191857, 32'sd0.026165492155860413, 32'sd-0.04251984945486247, 32'sd-9.008942125988033e-128, 32'sd0.0445426293708572, 32'sd-0.08547501727030613, 32'sd0.020811541791636367, 32'sd-0.030489097428001256, 32'sd-0.13286640733902205, 32'sd-0.007688983348462168, 32'sd-0.09696059860448115, 32'sd-0.0608968136677028, 32'sd-0.026386285277847383, 32'sd0.15557279117312253, 32'sd0.06803133598691724, 32'sd0.1155331893459193, 32'sd0.014980044771101852, 32'sd0.21844337740202854, 32'sd0.15137407151199142, 32'sd0.12424400909599696, 32'sd0.04979734915891145, 32'sd0.14991093985932014, 32'sd-0.015004204088579418, 32'sd0.1159988923330234, 32'sd0.06687210038585041, 32'sd-0.053391362625269036, 32'sd-0.03666950427920978, 32'sd0.09843609448686537, 32'sd0.01011927507427657, 32'sd-0.028560315298897097, 32'sd0.04503790820747252, 32'sd0.0376899298412588, 32'sd-0.026865226506173644, 32'sd-0.0012115387481813772, 32'sd0.008464628595562884, 32'sd0.10065445020260541, 32'sd0.061677155158309085, 32'sd-0.07139969196945607, 32'sd-0.09662625127101263, 32'sd-0.03796057479828352, 32'sd-0.0374291737255196, 32'sd0.04337680453617682, 32'sd0.03437779206283137, 32'sd-0.03549595999324536, 32'sd0.07768408266040265, 32'sd0.09652382327733756, 32'sd0.20277647911193855, 32'sd0.10300258981378908, 32'sd0.14868161843537006, 32'sd0.1296177238663857, 32'sd0.05928783438554996, 32'sd0.025258750359113843, 32'sd-0.04064002791773316, 32'sd-0.1646169727897144, 32'sd0.07800759250067849, 32'sd0.15834871985009244, 32'sd-0.025444733796018557, 32'sd0.08082327492200107, 32'sd-0.003235938947677701, 32'sd0.0887987750228831, 32'sd0.023896618801728536, 32'sd-0.043786651658663876, 32'sd0.029270894116339635, 32'sd0.11011928435780824, 32'sd0.0733498062355674, 32'sd0.03536850293985605, 32'sd-0.03528913617813128, 32'sd-0.1150070233933351, 32'sd0.024105895980508836, 32'sd-0.11439035606701585, 32'sd-0.05031273857302551, 32'sd-0.004271994230382738, 32'sd-0.025398620697534804, 32'sd-0.04025919835172651, 32'sd0.0490166986998681, 32'sd-0.015217877619302912, 32'sd-0.01932667843793836, 32'sd0.05817944879997445, 32'sd-0.036595256466731535, 32'sd0.020648615999570446, 32'sd0.0007707184202542456, 32'sd-0.0643783899429577, 32'sd-0.07664563848876924, 32'sd-0.060316249250286946, 32'sd0.039190013860713246, 32'sd0.048062214648343336, 32'sd0.04563220064518398, 32'sd-4.421130357642363e-119, 32'sd-0.017075059774998493, 32'sd0.000792504487959213, 32'sd-0.05435537597718715, 32'sd0.06530919001049097, 32'sd0.04945996754463158, 32'sd0.0660526550497986, 32'sd0.023518371713555693, 32'sd-0.0034562677189827464, 32'sd-0.10073783563644727, 32'sd-0.04718064350789281, 32'sd-0.03027132910417016, 32'sd-0.08284301935800342, 32'sd-0.029054827305666414, 32'sd-0.07095128368650351, 32'sd0.07760595539236574, 32'sd0.09231550624862736, 32'sd0.09835889374575053, 32'sd0.03361080415642212, 32'sd-0.028751102448477124, 32'sd0.07547898165659625, 32'sd0.028199572303400602, 32'sd-0.02561352300112504, 32'sd0.04056093347677394, 32'sd0.031209404543701694, 32'sd-0.06091749085359352, 32'sd-0.017377553836593895, 32'sd2.3335926118003127e-124, 32'sd-3.0750471172687936e-126, 32'sd-1.4358735755677674e-115, 32'sd0.03392048845227889, 32'sd-0.006846639917185744, 32'sd-0.054169438846400374, 32'sd-0.038252151820495794, 32'sd0.02813815097567269, 32'sd0.005189894122917695, 32'sd-0.012036906093491262, 32'sd0.03184746947715957, 32'sd0.047010035954098146, 32'sd0.050415536002761885, 32'sd-0.027528279990810076, 32'sd-0.015831664716681116, 32'sd0.06396187202428387, 32'sd-0.0002465733476639722, 32'sd0.09698806184481802, 32'sd0.037749598192288916, 32'sd0.032337575830374346, 32'sd0.07789146989273257, 32'sd0.029748538720287706, 32'sd0.06567375627907884, 32'sd0.0518185637691201, 32'sd0.10605406942392887, 32'sd-0.002701545100930447, 32'sd0.00693224325858246, 32'sd0.014198702095215338, 32'sd-2.282657563811111e-115, 32'sd7.893896309060512e-120, 32'sd6.688593419347141e-124, 32'sd-0.08219590350574926, 32'sd0.09073568491078186, 32'sd-0.05263603768025761, 32'sd-0.0518118180653605, 32'sd-0.02003047863492572, 32'sd0.03781472604743543, 32'sd-0.011085220683393033, 32'sd-0.026007392836622848, 32'sd-0.05836701781319779, 32'sd-0.046180211321006935, 32'sd0.00980722333906979, 32'sd-0.03948906972294798, 32'sd-0.014668582686396021, 32'sd0.03250644426416223, 32'sd-0.08811410528172989, 32'sd-0.00449594457437647, 32'sd-0.04066665194430565, 32'sd0.009686493924631036, 32'sd-0.06396723185357105, 32'sd0.04757233381281565, 32'sd0.08784630479235118, 32'sd0.032034186941842555, 32'sd-0.047769934832093, 32'sd0.01982123039701763, 32'sd0.09964560331387552, 32'sd-4.3702449960118215e-127, 32'sd-3.415614548209917e-126, 32'sd-1.5545608997637746e-117, 32'sd3.797141522782114e-122, 32'sd0.012171581146005148, 32'sd0.013669276519685868, 32'sd0.04436156073783827, 32'sd-0.1263189787296683, 32'sd-0.023440833005011708, 32'sd0.014405662987885618, 32'sd-0.15027269371748717, 32'sd-0.028452016566399514, 32'sd-0.0007098995712346846, 32'sd-0.043922971675937894, 32'sd-0.18678726357081193, 32'sd0.014387112096832981, 32'sd-0.010845170615560194, 32'sd0.0807578018887095, 32'sd0.118137705433484, 32'sd0.14024640011413061, 32'sd-0.056706779478589577, 32'sd-0.042498502232355684, 32'sd-0.0019458326502448083, 32'sd0.07926784340760086, 32'sd0.08028256895965484, 32'sd0.002160883277841964, 32'sd0.01019022162790391, 32'sd-4.793311163395595e-127, 32'sd3.9781594892984724e-115, 32'sd-6.432416997532629e-124, 32'sd1.6634856225931078e-125, 32'sd-7.051224405474324e-127, 32'sd-4.217323300101419e-117, 32'sd0.04433809140777269, 32'sd0.010902748960618625, 32'sd0.009199236473518389, 32'sd0.012681391654489591, 32'sd-0.04464100590373464, 32'sd-0.015583207015179398, 32'sd-0.06154090737302055, 32'sd-0.023443756159089058, 32'sd-0.07759374754672124, 32'sd0.058750076582342256, 32'sd0.12047196031925149, 32'sd0.01603280888422399, 32'sd0.0761458619729494, 32'sd-0.07361522845829511, 32'sd-0.06038975343824136, 32'sd-0.012161860063623554, 32'sd-0.06899266038864207, 32'sd0.017576571199814633, 32'sd-0.0899085755102439, 32'sd0.06310438135373996, 32'sd3.8309543855881135e-123, 32'sd1.1113507002368712e-121, 32'sd-5.537706173055546e-115, 32'sd5.57255195462053e-121},
        '{32'sd4.713588873914971e-128, 32'sd2.7737021065375e-119, 32'sd-3.212278771210468e-120, 32'sd-5.3738340726386335e-117, 32'sd-4.976191742747889e-115, 32'sd-1.8133815998849944e-119, 32'sd-8.685134576192346e-127, 32'sd-3.0774939763825874e-118, 32'sd7.561018891740884e-124, 32'sd4.3520805066008166e-123, 32'sd4.3278738216670114e-125, 32'sd-3.11650804181975e-116, 32'sd0.010809152982063294, 32'sd-0.029467094777021575, 32'sd0.08390327239625128, 32'sd0.11194046116801927, 32'sd5.6691109624355393e-126, 32'sd1.5994032046906875e-126, 32'sd1.1747988610285207e-123, 32'sd-1.1167207334222785e-119, 32'sd4.171506685079291e-118, 32'sd-4.343746490070249e-121, 32'sd8.572931951077343e-117, 32'sd5.443200309432459e-125, 32'sd-3.686763546289077e-121, 32'sd1.2241249237160504e-126, 32'sd6.796556261760817e-123, 32'sd-4.2709901238576516e-117, 32'sd1.1670283829465428e-115, 32'sd-6.349647008590328e-119, 32'sd-8.831438827148182e-123, 32'sd1.3996718524966424e-125, 32'sd-0.02824088794276072, 32'sd0.01801216282153803, 32'sd-0.095891508203206, 32'sd0.03345382630691873, 32'sd-0.09532645299554506, 32'sd-0.005131413841738006, 32'sd-0.012206106809170256, 32'sd-0.014093930727555635, 32'sd-0.031351594443468744, 32'sd0.1027452480731113, 32'sd0.06938446459873308, 32'sd0.057685874400387284, 32'sd-0.03133187110901903, 32'sd0.011333937677248497, 32'sd-0.03405047585045742, 32'sd-0.05242099921466428, 32'sd0.024471452994221706, 32'sd-0.007551569598910738, 32'sd0.04234864979430962, 32'sd0.05556745537789756, 32'sd9.09845072467746e-123, 32'sd-1.5182833577256937e-123, 32'sd-1.198103908174496e-122, 32'sd3.671882104148228e-126, 32'sd5.326785473889361e-118, 32'sd3.9802658047695885e-124, 32'sd0.10411465118514028, 32'sd0.014033821763626218, 32'sd-0.022627236283283184, 32'sd-0.04468277218884481, 32'sd0.05350583623434859, 32'sd0.003682869244483294, 32'sd0.017659931530502885, 32'sd0.005761260289811714, 32'sd0.12691384605145184, 32'sd0.04016249012181663, 32'sd0.11670496683840315, 32'sd0.1767406025172925, 32'sd0.08595412467765201, 32'sd0.0791224205197354, 32'sd-0.05817373607797154, 32'sd0.036160349770283415, 32'sd-0.05762259930623436, 32'sd-0.024383069982250302, 32'sd-0.005756190285878851, 32'sd0.055974536136693474, 32'sd-0.022040378036211786, 32'sd0.14863201264379422, 32'sd0.058104853622065133, 32'sd0.09463672176990699, 32'sd-2.7463072814242493e-118, 32'sd2.8387873889965944e-123, 32'sd1.3408733235653254e-122, 32'sd-3.5339047097019403e-122, 32'sd0.06233194795708739, 32'sd-0.008973818001713813, 32'sd-0.00977511706978159, 32'sd0.08434368347389092, 32'sd0.0005959806737388046, 32'sd0.08565713649006171, 32'sd-0.025064184795087145, 32'sd0.08417840710183364, 32'sd0.14483841699704827, 32'sd0.17618749884642337, 32'sd0.2771726787921846, 32'sd0.20244282605900843, 32'sd0.17907298405601185, 32'sd0.06337645876324904, 32'sd0.1916220463213292, 32'sd0.11975791413120238, 32'sd0.1979246485865861, 32'sd0.08154989555962079, 32'sd-0.026502395288491944, 32'sd-0.11100688395449437, 32'sd0.021118321775994292, 32'sd-0.12192568501860998, 32'sd0.06609514871524329, 32'sd0.007948257136289699, 32'sd-0.08941822957411918, 32'sd2.336512970187456e-125, 32'sd1.9627860110618533e-126, 32'sd0.03905587408691613, 32'sd0.045345121511533984, 32'sd0.0181558663318089, 32'sd-0.025801889475043395, 32'sd0.03517160127150294, 32'sd-0.027408109092171697, 32'sd-0.02694044519014569, 32'sd-0.048517009434296224, 32'sd-0.061776552416981906, 32'sd0.23415485369250008, 32'sd0.1467636947391649, 32'sd0.07866045135354022, 32'sd0.12023698060413547, 32'sd0.20607377801214155, 32'sd0.13692705814582828, 32'sd0.18382931857188606, 32'sd0.09760049421142171, 32'sd0.07519358760504431, 32'sd0.07503843824199466, 32'sd-0.014282748390725923, 32'sd-0.06114364625347711, 32'sd-0.09745436323916984, 32'sd-0.1313432460857387, 32'sd0.01952649135731089, 32'sd0.03303074336753134, 32'sd-0.04850137326829097, 32'sd0.014533718477315754, 32'sd-8.572739883561462e-117, 32'sd0.12516652758499414, 32'sd-0.062311261749392756, 32'sd0.012168466690553235, 32'sd-0.060376255185043116, 32'sd0.018806702934440686, 32'sd-0.043112586530518714, 32'sd-0.009639900576495901, 32'sd-0.14388563882601826, 32'sd-0.12232912321485899, 32'sd0.052751086387633164, 32'sd-0.0768962116759079, 32'sd0.052943158115107886, 32'sd0.04562755016064636, 32'sd0.05775386055859916, 32'sd0.1550302167754511, 32'sd0.09094670567641919, 32'sd0.033691429906993794, 32'sd0.165464364852574, 32'sd0.10945208393644165, 32'sd0.04864144953387694, 32'sd-0.014261639773447821, 32'sd0.08453999010437904, 32'sd0.05099175891367443, 32'sd0.03856146496345181, 32'sd0.03440130713042421, 32'sd-0.09361513301743452, 32'sd-0.03270164130326606, 32'sd6.155346007669574e-125, 32'sd0.08251199367439556, 32'sd-0.03331712906512036, 32'sd0.07954402174648699, 32'sd-0.13513385063922817, 32'sd-0.0007585160662327532, 32'sd-0.038674990781098845, 32'sd0.008964772637103763, 32'sd-0.06403252582667772, 32'sd-0.019293479235271974, 32'sd-0.011994173984718724, 32'sd-0.08863656226248114, 32'sd-0.1024232407284868, 32'sd0.12975457946700222, 32'sd0.03082897985059793, 32'sd-0.007349772794017511, 32'sd0.09132151778935471, 32'sd0.03835945969429856, 32'sd0.0727707093841672, 32'sd0.04699414951516187, 32'sd-0.013681855593095859, 32'sd-0.03493090811976986, 32'sd0.00694642964515282, 32'sd-0.021514960720915376, 32'sd0.059386107016396156, 32'sd-0.10049887316761685, 32'sd0.017414394071985025, 32'sd0.049043757902366, 32'sd0.0886783391809257, 32'sd0.07678139719757666, 32'sd0.048156143097175357, 32'sd0.08460431880483328, 32'sd-0.023656229725946557, 32'sd-0.06585796164386643, 32'sd0.02435882500505177, 32'sd-0.12771629106975615, 32'sd-0.12184820237589737, 32'sd-0.05593833184703442, 32'sd-0.12792343913221768, 32'sd-0.033521436456366176, 32'sd-0.09524199065081412, 32'sd-0.06516295460355688, 32'sd0.03105951843257499, 32'sd0.09534624312315294, 32'sd0.046830413818462154, 32'sd0.11550416782870704, 32'sd0.1392315185140413, 32'sd0.041689418013607184, 32'sd0.03431971712093007, 32'sd0.04420458019302651, 32'sd0.08792929227010374, 32'sd0.06797286578189929, 32'sd0.0319146838346131, 32'sd-0.05391544727997319, 32'sd0.010497130410814398, 32'sd0.05106672639224898, 32'sd0.03416088915691843, 32'sd0.03603008132520514, 32'sd-0.00882458337779432, 32'sd-0.06369221419966628, 32'sd-0.02773636466528516, 32'sd-0.1295307566693657, 32'sd-0.08001116377017581, 32'sd-0.08209540267730422, 32'sd-0.029525628497618153, 32'sd0.10112664065278736, 32'sd-0.004800724846156721, 32'sd-0.16394495505298023, 32'sd-0.12068565430368006, 32'sd-0.16179977216765526, 32'sd-0.08197588513746774, 32'sd-0.09159500767937237, 32'sd0.04620841707251492, 32'sd0.12670034625703552, 32'sd0.04667150544149333, 32'sd0.09233771008371029, 32'sd0.04627382060752612, 32'sd0.0402301411283871, 32'sd-0.005590099217496658, 32'sd0.01682137306304068, 32'sd-0.15029406106443358, 32'sd0.026329637052240805, 32'sd0.007940794905310501, 32'sd0.06194880748217137, 32'sd0.014954213977766568, 32'sd-0.04170500915936419, 32'sd-0.043004794574164514, 32'sd0.08782818991562487, 32'sd-0.023925919948466073, 32'sd-0.10411503954316723, 32'sd-0.09649717240784475, 32'sd-0.08777898233736427, 32'sd-0.1630725622966383, 32'sd-0.04160276099145361, 32'sd-0.19494994315854258, 32'sd-0.3249072859615802, 32'sd-0.3215764188589842, 32'sd-0.286568961817987, 32'sd-0.0893198998382284, 32'sd-0.08293583598915318, 32'sd0.026451868190929387, 32'sd0.11965113860952176, 32'sd0.05260183296862559, 32'sd0.07714477301780683, 32'sd0.07606426851459555, 32'sd0.1157453246764381, 32'sd-0.05435016877904393, 32'sd0.006047601008568124, 32'sd-0.06453624680213672, 32'sd-0.029708047584965633, 32'sd-0.011774435864002718, 32'sd0.005578931050437378, 32'sd0.05417582102686271, 32'sd-0.06446233346131214, 32'sd0.0575272370965593, 32'sd0.06316102465688814, 32'sd0.03226664806082336, 32'sd-0.001470943418267691, 32'sd-0.10859003969203, 32'sd-0.22244933837495098, 32'sd-0.26140185665879767, 32'sd-0.1658810366129804, 32'sd-0.2319995031244143, 32'sd-0.3996586762196566, 32'sd-0.21893281990037236, 32'sd-0.17738591397741707, 32'sd0.056852425369550076, 32'sd-0.05025131758291568, 32'sd0.03764057602710154, 32'sd-0.0221497526709715, 32'sd-0.0036758550245675043, 32'sd-0.017352039528350502, 32'sd-0.0062071671576576105, 32'sd0.05250270263566315, 32'sd-0.0394697231124059, 32'sd-0.03649265457161631, 32'sd-0.06552588509239166, 32'sd0.024671147218781726, 32'sd-0.02316048516422793, 32'sd-0.04815063391199418, 32'sd-0.02134513072096698, 32'sd0.051038742570455084, 32'sd0.03765841464694719, 32'sd-0.04639720472735638, 32'sd-0.0711150624978682, 32'sd-0.20194325407815866, 32'sd-0.18932345699149133, 32'sd-0.23671125088667078, 32'sd-0.2590497776449477, 32'sd-0.15065549851055976, 32'sd-0.1624778298751745, 32'sd-0.2720139050065402, 32'sd-0.16626736700159353, 32'sd0.048521815798995754, 32'sd0.14346463611277768, 32'sd0.09364714333848884, 32'sd-0.1967619646167437, 32'sd-0.019261142949585905, 32'sd-0.08342247766970531, 32'sd0.02751939312032188, 32'sd-0.014636831167097733, 32'sd0.004522609729297693, 32'sd0.09056491779712202, 32'sd-0.0184189734258891, 32'sd-0.1717107818188698, 32'sd-0.020281374174867993, 32'sd-0.08687595372823569, 32'sd0.007338446483673774, 32'sd0.07376269043786465, 32'sd-0.07300426751754137, 32'sd-0.09748582545656934, 32'sd-0.0730988410251361, 32'sd-0.1758117306114292, 32'sd-0.08012229488359603, 32'sd-0.11330511748205165, 32'sd-0.1412190996456023, 32'sd-0.040251369231762875, 32'sd-0.028527314438205532, 32'sd-0.0316030071423673, 32'sd0.012052130394263085, 32'sd0.11007529201245661, 32'sd0.11207448082815118, 32'sd0.17888323308719636, 32'sd0.07143674729606274, 32'sd-0.10230824729679663, 32'sd-0.10912580894440106, 32'sd-0.007813140590585771, 32'sd-0.15834519409728684, 32'sd-0.17361745394618694, 32'sd0.02917422368733901, 32'sd-0.049840498259933995, 32'sd-0.018784956151521343, 32'sd-0.1551188431212078, 32'sd-0.10271502722880102, 32'sd-0.029895018330832624, 32'sd0.040398506680982105, 32'sd0.06421836116723942, 32'sd-0.04258553337271913, 32'sd0.01843623041927533, 32'sd-0.024524729470053193, 32'sd-0.026540025303879628, 32'sd-0.1104268079963789, 32'sd-0.09519350256307589, 32'sd0.035774296912181, 32'sd-0.002215433085727866, 32'sd0.13341310859095823, 32'sd0.11868772650299003, 32'sd0.18786461542678745, 32'sd0.135500405498253, 32'sd0.1535293490941635, 32'sd0.20510612457745853, 32'sd-0.01386904896832457, 32'sd-0.061941635766140715, 32'sd-0.1432703435505243, 32'sd-0.010296103082654419, 32'sd-0.15877097335071721, 32'sd-0.0031462112808894292, 32'sd0.021100048588004964, 32'sd0.036810975047669656, 32'sd0.11024756949218195, 32'sd-0.04050969432170025, 32'sd0.0035160759658722333, 32'sd0.015421134461339057, 32'sd0.07295917068808772, 32'sd0.057600348776788275, 32'sd-0.01844689828247562, 32'sd0.03445830632258352, 32'sd0.006976773403358526, 32'sd0.1599808145610909, 32'sd0.1256724195097125, 32'sd0.08258092793364584, 32'sd0.09400446276002697, 32'sd0.19438866012917033, 32'sd0.15565173283180067, 32'sd0.15364222470735645, 32'sd0.0400543116561809, 32'sd0.09773707757349309, 32'sd-0.0466777482887113, 32'sd0.02146964153528286, 32'sd-0.04014741424122224, 32'sd-0.026604126542767125, 32'sd0.03255114793678448, 32'sd0.11406968493994352, 32'sd-0.012726081780000889, 32'sd-0.07634284583097045, 32'sd-0.00490502529301015, 32'sd-0.010316950838083825, 32'sd0.05149742069724497, 32'sd0.03951417310921872, 32'sd0.01448716008922159, 32'sd-0.08359109904474767, 32'sd0.08420977169948335, 32'sd-0.06878205907240519, 32'sd-0.00014313956020368365, 32'sd-0.04372530432050575, 32'sd0.07492031857028804, 32'sd0.1348328224516303, 32'sd0.07112433667670293, 32'sd0.015503406391808234, 32'sd0.10206606641362177, 32'sd0.08751552756920558, 32'sd0.006018128037124817, 32'sd0.006466056414911061, 32'sd0.04886335334989602, 32'sd-0.11713226632046339, 32'sd-0.18109043735722302, 32'sd-0.10155216889021262, 32'sd-0.06978496455153088, 32'sd-0.01643837795052636, 32'sd0.07501128964208045, 32'sd0.028167101974377884, 32'sd-0.04130954216216003, 32'sd-0.13072391346128262, 32'sd0.052468017830921594, 32'sd0.022986348830263747, 32'sd-0.0782419865378755, 32'sd-0.06761686395981671, 32'sd-0.04941227930617381, 32'sd0.03979114666434608, 32'sd0.053496914956507, 32'sd0.07571799088909023, 32'sd0.07687593072567274, 32'sd0.016609587470101606, 32'sd-0.03305954606146289, 32'sd0.07282673007529027, 32'sd0.09669555908167125, 32'sd-0.02567062355390636, 32'sd0.08246841179865957, 32'sd-0.020482423254779978, 32'sd0.04359704903733148, 32'sd-0.019782112544081822, 32'sd0.015559770862889582, 32'sd-0.028784821879640505, 32'sd-0.136472688648362, 32'sd-0.16964853691080817, 32'sd0.050355191926336085, 32'sd0.03213663606569373, 32'sd0.22320149034833642, 32'sd0.07356649480808976, 32'sd0.06642586691960592, 32'sd-0.00248043333683055, 32'sd0.028897434800225427, 32'sd0.018165309881096593, 32'sd-0.012350639753800876, 32'sd-0.003918520466428085, 32'sd0.02306246951548991, 32'sd0.08955651537912597, 32'sd0.06920372625017787, 32'sd5.703340551999425e-124, 32'sd0.003173653275757202, 32'sd0.07445222492315924, 32'sd0.038466727579173576, 32'sd0.007512456067037591, 32'sd-0.016713671910094485, 32'sd0.04144123005352018, 32'sd0.0678029728938625, 32'sd-0.025682804821641106, 32'sd0.033414732366852704, 32'sd-0.04667487297169402, 32'sd0.027880810272391476, 32'sd-0.18533619234319704, 32'sd-0.21685763092890548, 32'sd-0.10236911749167717, 32'sd0.02750611984018655, 32'sd0.23739625401741457, 32'sd0.1455383526572352, 32'sd0.1561039059247564, 32'sd0.0918399845628874, 32'sd0.03433720353195714, 32'sd0.135140396447417, 32'sd0.019042589767372206, 32'sd0.022042274592597066, 32'sd0.06060231091531795, 32'sd0.04540459986898374, 32'sd0.010980966997334436, 32'sd0.03919782629290038, 32'sd0.02491570665529667, 32'sd0.0782856961755123, 32'sd0.1003592235004638, 32'sd0.12486032812381216, 32'sd0.03583091337523244, 32'sd0.07784637766983953, 32'sd0.028114704672576964, 32'sd0.029966463381270972, 32'sd0.009843832887387828, 32'sd0.022204103095963885, 32'sd-0.06092219926886588, 32'sd0.030301539094667318, 32'sd-0.19235037287084802, 32'sd-0.12109280571959585, 32'sd0.015452401082693091, 32'sd0.08001412745879244, 32'sd0.10611336708103403, 32'sd0.12387194699649288, 32'sd0.08184815535980156, 32'sd-0.04949471076344423, 32'sd0.016928637279111307, 32'sd0.040289372914571235, 32'sd-0.006442975098159557, 32'sd0.023046201922557092, 32'sd-0.05557069906405803, 32'sd0.06443641012989657, 32'sd-0.07471108244420593, 32'sd0.011225268001162001, 32'sd0.07142918079831445, 32'sd-0.024277912726677113, 32'sd-0.025030734858346074, 32'sd-0.033507411154935045, 32'sd-0.014177465289130432, 32'sd0.02797478610529085, 32'sd0.04077244130305591, 32'sd0.052784851918795526, 32'sd0.02662964615249291, 32'sd-0.033640934855364166, 32'sd-0.016529572486863025, 32'sd-0.11370713235573907, 32'sd-0.018709967185943005, 32'sd0.04595746145173994, 32'sd0.022395247788894374, 32'sd0.22755044085269094, 32'sd0.09682217921709112, 32'sd-0.02196499793731679, 32'sd-0.01778795452452906, 32'sd-0.09198587746776224, 32'sd-0.08877678335223221, 32'sd-0.026201101783271136, 32'sd-0.019559410085120393, 32'sd-0.08244465012429011, 32'sd-0.04971834866200679, 32'sd-0.11255335296574825, 32'sd0.07823999201297759, 32'sd0.0014811662494434515, 32'sd-4.581017366634545e-118, 32'sd0.053426303062643295, 32'sd0.08437507638965643, 32'sd0.0712685673945568, 32'sd-0.057695118935740974, 32'sd0.01686251989720322, 32'sd0.12611533879330025, 32'sd0.07194153671130128, 32'sd0.038859128730468324, 32'sd0.047474820700407955, 32'sd0.08250330722686683, 32'sd0.07020905252993602, 32'sd0.14013631676695487, 32'sd0.059976725090261356, 32'sd-0.017742350640301607, 32'sd-0.1156557415443799, 32'sd0.09336845224262323, 32'sd0.04537746559737883, 32'sd-0.07950300996582067, 32'sd-0.1448834067043724, 32'sd-0.0914995854460871, 32'sd-0.12104314531381413, 32'sd-0.033891193256270304, 32'sd-0.08082405342005454, 32'sd-0.0014273505043425232, 32'sd-0.07629146584060652, 32'sd-0.03632163179102486, 32'sd0.0445479757213522, 32'sd-0.0157744008747399, 32'sd-0.03473616161137983, 32'sd0.010066142641633236, 32'sd0.10627274648037426, 32'sd0.042605331857473776, 32'sd-0.07723654945671789, 32'sd0.07825796580908072, 32'sd0.016968074474386297, 32'sd0.13433240509293487, 32'sd-0.05743107859482347, 32'sd0.012755529917130843, 32'sd0.05370136779487479, 32'sd0.07772527633952421, 32'sd-0.06348148981275994, 32'sd-0.10836472834165478, 32'sd-0.13598090692396728, 32'sd-0.09029272814081223, 32'sd-0.06110068002439528, 32'sd-0.0977387967925267, 32'sd-0.052061952649075635, 32'sd-0.018918407092771074, 32'sd-0.019357024283409175, 32'sd0.0220006852602129, 32'sd0.1022796937471154, 32'sd-0.13209651225004318, 32'sd0.0058637552765527165, 32'sd0.02939789068893449, 32'sd0.010191312261310917, 32'sd-0.011727463465578876, 32'sd0.06311543733889516, 32'sd0.07409694336732957, 32'sd-0.048405168574453435, 32'sd-0.027138083095378348, 32'sd-0.08551665772236854, 32'sd0.11515183370283803, 32'sd0.11647054696467418, 32'sd0.001588644698843463, 32'sd-0.07416926764678533, 32'sd-0.02143505455171051, 32'sd3.9648946443945185e-05, 32'sd0.038597710598817746, 32'sd0.06279036236242502, 32'sd-0.04590559556006543, 32'sd-0.028117638511947707, 32'sd-0.07363205830971037, 32'sd-0.054016510378840164, 32'sd-0.03098591427105729, 32'sd-0.01171851476163358, 32'sd-0.03780872191542429, 32'sd0.07409044267474171, 32'sd0.08083325335394684, 32'sd-0.06524717699149968, 32'sd0.028405714810892865, 32'sd-0.01726949985958659, 32'sd-0.04341590499852661, 32'sd0.07131814462013428, 32'sd2.0022729703333189e-116, 32'sd0.06574736719784818, 32'sd-0.05871405492491691, 32'sd-0.023110693579752917, 32'sd0.05263070682981631, 32'sd-0.03634597947311368, 32'sd-0.0405764515806636, 32'sd-0.0243274841293653, 32'sd-0.07984339234874674, 32'sd0.06115304072113684, 32'sd0.06870324877764061, 32'sd0.11704952797496661, 32'sd0.15809744889907498, 32'sd0.025655961693844865, 32'sd0.0529775408801077, 32'sd-0.07909743426767324, 32'sd-0.07620586151804717, 32'sd-0.15083250497744333, 32'sd-0.1868480726829186, 32'sd-0.0152016154921079, 32'sd0.03435416399749469, 32'sd-0.010816893423208853, 32'sd0.017476929057145475, 32'sd-0.12111446432717378, 32'sd0.05553445525744147, 32'sd0.06345258993375322, 32'sd0.062197145543198065, 32'sd-4.327018197411949e-125, 32'sd-8.069592844311294e-118, 32'sd-8.691037050379299e-128, 32'sd-0.00744663755388275, 32'sd0.039630761920962744, 32'sd0.08663696359372441, 32'sd-0.02695069844454985, 32'sd0.014716758534151534, 32'sd-0.006376632646164977, 32'sd0.12999399566813233, 32'sd0.06235842676376187, 32'sd-0.10803376822161172, 32'sd-0.0007589381581551068, 32'sd-0.03396690817681119, 32'sd-0.02891461732916995, 32'sd0.04645551434798777, 32'sd0.06971564742401179, 32'sd-0.14089371985370297, 32'sd-0.16326088389573673, 32'sd-0.08810685968551478, 32'sd-0.06024911542839833, 32'sd0.07997526934157667, 32'sd-0.05714568242339129, 32'sd0.030723842111797135, 32'sd0.03773918677131916, 32'sd0.04634098831944694, 32'sd-0.00673614926098317, 32'sd0.07740656388509337, 32'sd-8.903826890898e-127, 32'sd2.4740800169290727e-117, 32'sd-1.3142944261528025e-122, 32'sd0.09055003394198233, 32'sd-0.06288595675905495, 32'sd0.020529426792477396, 32'sd0.008782779869028319, 32'sd-0.02414938812781218, 32'sd-0.14418292254884957, 32'sd-0.038517782929442024, 32'sd-0.08112173756232854, 32'sd-0.1367094054919934, 32'sd-0.03333898786239195, 32'sd-0.10424482443355126, 32'sd-0.012343969706917994, 32'sd0.02179128825210423, 32'sd-0.06428877610409334, 32'sd-0.011715639054076672, 32'sd0.018627932545312798, 32'sd0.01295469461898409, 32'sd0.08344414423017349, 32'sd0.05421054771877751, 32'sd-0.03803356689829162, 32'sd-0.04738922736497144, 32'sd-0.11199891652581183, 32'sd0.009576808350984, 32'sd0.03656920838891924, 32'sd-0.05384509608940687, 32'sd6.965284117138896e-121, 32'sd1.5748181508097428e-125, 32'sd1.6123759449809133e-125, 32'sd1.0775699471490713e-124, 32'sd0.0974135261147584, 32'sd0.027633076930406026, 32'sd0.06887222913996004, 32'sd0.027988458629822126, 32'sd0.0010779189199772387, 32'sd-0.059396533114616394, 32'sd0.011193663579433003, 32'sd0.09208168571699125, 32'sd-0.003347293369323064, 32'sd0.0345686253461147, 32'sd0.08277746096974048, 32'sd0.12795028012886014, 32'sd0.09169386041224586, 32'sd0.031375355119376516, 32'sd-0.026650807539361623, 32'sd0.061335318354635744, 32'sd-0.004387443170558067, 32'sd0.012196148133810213, 32'sd-0.05050096459854837, 32'sd-0.027554747110147042, 32'sd-0.012201481137568951, 32'sd0.02073428333213612, 32'sd0.03141434473872971, 32'sd-1.6153978920848175e-115, 32'sd-4.7125339489901474e-123, 32'sd7.659439980705893e-121, 32'sd2.4275599732113302e-126, 32'sd-5.061523235634357e-118, 32'sd4.7481704738339556e-123, 32'sd0.07217429133693033, 32'sd-0.02154347700215209, 32'sd0.07269457837770113, 32'sd-0.051723545016263035, 32'sd0.04743860634487606, 32'sd-0.003705406757635343, 32'sd0.05636892242750938, 32'sd0.0717829967454534, 32'sd0.05460578678795196, 32'sd0.07299412521131225, 32'sd0.08771230604114101, 32'sd0.07508451728492001, 32'sd0.08592304432424144, 32'sd0.14223058429305874, 32'sd0.05048431354386904, 32'sd0.07202503847122105, 32'sd0.028599136808309986, 32'sd-0.013029425603040221, 32'sd0.09544627051090535, 32'sd0.0538454582236887, 32'sd2.471741288636203e-124, 32'sd-8.555494534816719e-126, 32'sd8.128031635038046e-117, 32'sd3.509766378707519e-115},
        '{32'sd-3.7041488165993343e-116, 32'sd-3.7766866681522155e-128, 32'sd1.2868924977672362e-118, 32'sd-2.6375907575887196e-124, 32'sd-9.852827182992159e-118, 32'sd-2.6272076079803646e-116, 32'sd5.899697450134656e-116, 32'sd3.210388971348045e-121, 32'sd5.39385741439986e-118, 32'sd3.55765466602173e-114, 32'sd-3.0071454952325037e-119, 32'sd4.840689624625377e-128, 32'sd-0.004135142355679971, 32'sd-0.0003237971801643967, 32'sd0.0014468247772041884, 32'sd-0.03405848223243477, 32'sd2.3734292838395237e-122, 32'sd-1.5926357842976516e-121, 32'sd-8.955436658075706e-120, 32'sd-1.542312297081881e-123, 32'sd1.4547752010627164e-127, 32'sd-7.87731230820166e-121, 32'sd-1.4898723815956762e-117, 32'sd6.349778064414776e-119, 32'sd-2.0562117522842626e-115, 32'sd-4.296219062791963e-125, 32'sd1.3898181725514346e-116, 32'sd1.0108003910246849e-123, 32'sd-1.7153136430042573e-125, 32'sd-3.8901568423715603e-119, 32'sd-4.62582983739863e-123, 32'sd-2.7196677746897835e-116, 32'sd0.0011532516381201074, 32'sd-0.04853617868635363, 32'sd-0.009671379878999537, 32'sd0.004410801456439582, 32'sd0.009617102405734497, 32'sd-0.011433309109724139, 32'sd-0.03430368720460937, 32'sd0.04464995183833517, 32'sd-0.04814786577926199, 32'sd0.03222153752899917, 32'sd-0.0056349733815257794, 32'sd0.025130176738660207, 32'sd0.043120652062397825, 32'sd0.041495946263346156, 32'sd-0.009872951979955882, 32'sd0.04518099371366996, 32'sd-0.07462468172336921, 32'sd0.029981948597701945, 32'sd-0.008074266530497184, 32'sd-0.026260805538644173, 32'sd-5.984981167182643e-123, 32'sd3.738891720119678e-129, 32'sd9.641536152479591e-121, 32'sd3.9515028863185735e-125, 32'sd7.335826195683415e-117, 32'sd-6.102267165054473e-126, 32'sd0.025851406924119212, 32'sd-0.04757750222390769, 32'sd-0.03868400986542637, 32'sd-0.011278049721857782, 32'sd-0.07666712597077524, 32'sd0.04470196064145077, 32'sd0.07461130622385263, 32'sd-0.08075279753814378, 32'sd0.0047663689391405, 32'sd-0.0041296667924335135, 32'sd-0.00889505133822837, 32'sd0.06882925323408756, 32'sd-0.0011080507189616712, 32'sd-0.10070148063375543, 32'sd-0.103560277778068, 32'sd-0.06254423235086062, 32'sd0.017295743815666814, 32'sd-0.017490643937041903, 32'sd0.02327724722080926, 32'sd-0.09016532733824623, 32'sd0.04971841110615386, 32'sd-0.07486902942200936, 32'sd0.02301947400985256, 32'sd0.02126012895518425, 32'sd3.908990256149326e-124, 32'sd-7.100230339018982e-126, 32'sd1.4108669965814018e-118, 32'sd1.0409999284662986e-124, 32'sd0.04264991261110113, 32'sd-0.04904276526154323, 32'sd0.0320254828926374, 32'sd-0.08197326499305664, 32'sd-0.0752551490566105, 32'sd-0.057949248074697673, 32'sd0.040877844936897424, 32'sd-0.06081019177504311, 32'sd-0.0782584249325095, 32'sd-0.07776179160134003, 32'sd-0.05350079816059981, 32'sd-0.03703158023799334, 32'sd-0.11439487433018805, 32'sd-0.05348053249769458, 32'sd-0.07003870390707695, 32'sd0.01991543622361494, 32'sd0.044562242918504996, 32'sd0.02326423064760415, 32'sd0.027457255994038313, 32'sd0.08529533574472302, 32'sd-0.01811114970937452, 32'sd-0.025479070910626112, 32'sd0.08610119837635606, 32'sd-0.01603005073799357, 32'sd0.05377112436111255, 32'sd2.2524967022604284e-121, 32'sd-3.4219387772510596e-125, 32'sd0.017554422828098975, 32'sd0.0068435092867974775, 32'sd0.0038781130447196597, 32'sd-0.08971560437181565, 32'sd-0.08027726346853012, 32'sd-0.07966142645602944, 32'sd-0.10528094011914853, 32'sd-0.11951061156898071, 32'sd-0.15275238141400746, 32'sd-0.17838809560770694, 32'sd-0.05833511263764722, 32'sd-0.08136812288519954, 32'sd-0.08741390077362972, 32'sd-0.1607787670486298, 32'sd-0.1026601607694703, 32'sd-0.0331031448307124, 32'sd0.0701958418723283, 32'sd0.19510816354252788, 32'sd0.1691419920652651, 32'sd0.032678973532161426, 32'sd-0.012169806098944967, 32'sd0.05583330360909754, 32'sd-0.08735148868619304, 32'sd0.011027399480210273, 32'sd-0.09729223909994748, 32'sd0.09965730136446178, 32'sd0.05306490811700808, 32'sd-1.9317335993168277e-125, 32'sd-0.03271700215423605, 32'sd0.07952910033880813, 32'sd-0.002339295618263894, 32'sd-0.05646316873111512, 32'sd-0.037442710171143506, 32'sd-0.04980443874082898, 32'sd-0.1253052852764122, 32'sd-0.09238128974835728, 32'sd-0.08455793394040559, 32'sd-0.11171020618711582, 32'sd-0.06623901821116028, 32'sd-0.07048928156075376, 32'sd-0.05892794101567439, 32'sd-0.021050132481667965, 32'sd-0.06745810083298798, 32'sd-0.07226273635540668, 32'sd-0.09514882886320852, 32'sd0.11265825383253891, 32'sd0.14724625795953403, 32'sd0.10525479420981079, 32'sd-0.009732231616079312, 32'sd0.07931969257661535, 32'sd-0.028192236662022845, 32'sd-0.011333367774519054, 32'sd0.10919211440206203, 32'sd0.06552600064288605, 32'sd0.02736897222961538, 32'sd-2.5844138408670846e-124, 32'sd-0.004889121862547487, 32'sd-0.022454575575421958, 32'sd-0.02251260021836387, 32'sd0.06381748110280264, 32'sd-0.056267595094544945, 32'sd0.05046044500070395, 32'sd-0.053231713035902635, 32'sd-0.14310085574744866, 32'sd-0.007565580990840802, 32'sd-0.09284321687873234, 32'sd-0.023606947458193965, 32'sd-0.11655000479517043, 32'sd-0.014946167902448806, 32'sd0.09992143261493636, 32'sd0.010883487960792143, 32'sd0.018379359449264842, 32'sd0.022204014937183464, 32'sd0.019696767742420494, 32'sd-0.09082158987576709, 32'sd-0.14045251176296067, 32'sd-0.07115734282977951, 32'sd-0.09070544024165236, 32'sd-0.005218611102106566, 32'sd0.003796530661367764, 32'sd0.027986507973603445, 32'sd0.040818087336914395, 32'sd0.04290985894356727, 32'sd0.019821674445273024, 32'sd-0.06426779625251378, 32'sd0.008353620950658927, 32'sd-0.046168568220393225, 32'sd-0.005186586220200341, 32'sd-0.006109779719856775, 32'sd-0.043171122955556473, 32'sd-0.12516066821118618, 32'sd-0.08217623660409536, 32'sd-0.19857653686189705, 32'sd-0.11464754942111353, 32'sd-0.050952375827397076, 32'sd0.025736397441793353, 32'sd0.05602103703372009, 32'sd0.006353045564314876, 32'sd0.10320656876002879, 32'sd0.0030496723469265363, 32'sd0.04044367475857124, 32'sd0.04007438652218075, 32'sd0.004655865589015455, 32'sd0.07346930038600011, 32'sd-0.07082196763443344, 32'sd0.06965318347035951, 32'sd0.04488420226873522, 32'sd-0.0492515906375551, 32'sd0.01234597019238344, 32'sd0.05045372074958812, 32'sd0.008107645570436686, 32'sd-0.03973814734119293, 32'sd0.061871803217289495, 32'sd-0.025206590191247973, 32'sd-0.07989330571218273, 32'sd-0.006175364414846166, 32'sd-0.07129760052610232, 32'sd-0.11440602532017369, 32'sd-0.1228687602618594, 32'sd-0.0875616921183507, 32'sd-0.07064511348398776, 32'sd-0.0671451165470574, 32'sd-0.023951912756901953, 32'sd0.1054729531716065, 32'sd0.0160558429890137, 32'sd0.01250235421280373, 32'sd0.0007492365338074074, 32'sd-0.01661322913949487, 32'sd0.04314631176289953, 32'sd-0.012040419874699226, 32'sd0.15795081551575268, 32'sd0.07153581744750837, 32'sd-0.015420379515860644, 32'sd0.05908023819344037, 32'sd-0.12458838756366562, 32'sd0.01510610189185755, 32'sd-0.009613242615669797, 32'sd0.04987977318073886, 32'sd0.057908748635256434, 32'sd-0.04252898953737517, 32'sd-0.013782042537350232, 32'sd-0.054416279982741365, 32'sd-0.08467209637268247, 32'sd0.08494947765546056, 32'sd-0.08395241176280897, 32'sd-0.031899080697515514, 32'sd-0.12084439029266716, 32'sd-0.06179758085365535, 32'sd0.1152490343982287, 32'sd0.19977981264840333, 32'sd0.017367130472429895, 32'sd-0.017744324301303283, 32'sd0.04479339043617672, 32'sd-0.20463716206480084, 32'sd-0.13449432361287184, 32'sd-0.0179570959454226, 32'sd0.18285699667077618, 32'sd0.1796442015422375, 32'sd0.11995371003389924, 32'sd0.07201404464828089, 32'sd0.139539684003555, 32'sd-0.07046321525837125, 32'sd-0.09813667203189567, 32'sd-0.08622282874198244, 32'sd0.03165122355671253, 32'sd0.01849529248765711, 32'sd-1.3985476610875682e-05, 32'sd-0.061681924733141553, 32'sd-0.008934110136323559, 32'sd-0.16271049477125296, 32'sd-0.06604592549146847, 32'sd-0.0004551912248256195, 32'sd-0.07577898818393394, 32'sd-0.10336471953077861, 32'sd0.03549153628811155, 32'sd0.13527188491084172, 32'sd0.18404491683357754, 32'sd0.051249029529010066, 32'sd0.03582093892307587, 32'sd-0.017920176061946184, 32'sd-0.1623450016458891, 32'sd-0.050682537183030694, 32'sd-0.04275568981377509, 32'sd0.07630414073076956, 32'sd0.09249387401688323, 32'sd0.18673450814814843, 32'sd0.12755421178427184, 32'sd0.055970806857158974, 32'sd-0.05024571462424685, 32'sd-0.01650204951918083, 32'sd-0.006953722215409393, 32'sd-0.15229651688279247, 32'sd0.03780645786309562, 32'sd0.06085149389126068, 32'sd0.08701407272242241, 32'sd-0.006764045555988129, 32'sd-0.06238029614018581, 32'sd-0.11725096830856764, 32'sd-0.0801842994108062, 32'sd-0.012273402406045896, 32'sd-0.009616013622986096, 32'sd0.07117619543004201, 32'sd0.04803277952676108, 32'sd0.09831703498624006, 32'sd0.05780131427983883, 32'sd-0.07560775206949676, 32'sd-0.18641252463408542, 32'sd-0.19503097928963664, 32'sd-0.15120673609192142, 32'sd-0.05094999807838365, 32'sd0.03531336023305418, 32'sd0.15286090506389255, 32'sd0.14992839901515567, 32'sd0.11200715609302056, 32'sd0.14311456411644616, 32'sd0.1835976428561385, 32'sd0.06268505754837762, 32'sd-0.02695644928099521, 32'sd-0.10793336337245141, 32'sd-0.09414677769579674, 32'sd0.06336559705572213, 32'sd-0.011997813110552015, 32'sd-0.0006298290120910143, 32'sd-0.035375377161296406, 32'sd-0.0004504591127048399, 32'sd-0.05233012111318458, 32'sd-0.04992999672911005, 32'sd0.07554167068959276, 32'sd0.08151961876608851, 32'sd0.07422461844133804, 32'sd0.06578495184866985, 32'sd-0.009596745754192969, 32'sd-0.05216628829905482, 32'sd-0.18899772339024962, 32'sd-0.12460667481047182, 32'sd-0.07473872290353822, 32'sd0.014509232513034188, 32'sd0.1153814783162874, 32'sd0.22522903534705513, 32'sd0.19576656473589107, 32'sd0.21866347248960075, 32'sd0.19483187203254818, 32'sd0.18112846002455713, 32'sd0.16133861490058682, 32'sd0.02212931811828339, 32'sd0.025999142340108524, 32'sd0.012255491598719592, 32'sd-0.12497714964145758, 32'sd0.034966308853480434, 32'sd0.03752465595433956, 32'sd-0.04170845567921764, 32'sd0.051666005549866945, 32'sd-0.044437775563634686, 32'sd0.052611309721600275, 32'sd-0.12616058114368023, 32'sd0.011832366536872281, 32'sd0.0241388683483552, 32'sd0.11225043162598437, 32'sd-0.07624811993848861, 32'sd-0.031404186169629575, 32'sd-0.18949668858853091, 32'sd-0.13886262297690424, 32'sd-0.08181486243302445, 32'sd-0.06909686142171104, 32'sd0.11725506655945582, 32'sd0.29237446763614877, 32'sd0.20438831723043116, 32'sd0.13988496719107915, 32'sd0.13831026188992793, 32'sd0.1692072575709376, 32'sd0.060499180492274526, 32'sd-0.06710484061861165, 32'sd-0.0032784354264981524, 32'sd-0.03986704286314013, 32'sd-0.15638345038041673, 32'sd-0.15078181426144224, 32'sd-0.06476854831763641, 32'sd0.03832470777428478, 32'sd-0.06261811936995235, 32'sd-0.04022975832402921, 32'sd-0.02683861456483175, 32'sd-0.10614886311392907, 32'sd-0.10985590167874987, 32'sd0.03594939437716428, 32'sd-0.062458246116803666, 32'sd-0.027825603966046393, 32'sd-0.10715105333087561, 32'sd-0.04450766421930053, 32'sd-0.09044137074343833, 32'sd-0.02392331323286807, 32'sd0.07896052218447547, 32'sd0.14653766619791855, 32'sd0.11438188811571923, 32'sd0.23346141217506727, 32'sd0.16183767523367135, 32'sd0.0909244171329411, 32'sd0.0016761099625918665, 32'sd0.08225244583372825, 32'sd-0.04797111483970869, 32'sd-0.11938415417417762, 32'sd-0.1582062614141102, 32'sd0.01838220701708845, 32'sd0.06833150813295324, 32'sd-0.009778625119939498, 32'sd0.07885045617143842, 32'sd0.005438789307156673, 32'sd-0.025504147304691988, 32'sd0.05327101630531655, 32'sd-0.040845663458354144, 32'sd-0.07945019398771236, 32'sd-0.08740628290795897, 32'sd0.0456581050504383, 32'sd0.007607792518581848, 32'sd-0.02415271480784986, 32'sd-0.009841970981124777, 32'sd-0.020477580500496348, 32'sd-0.1089171662171056, 32'sd-0.1284444618778144, 32'sd-0.036836071393669526, 32'sd0.11241455908489188, 32'sd0.14025375533740125, 32'sd0.07429325126635551, 32'sd0.023017391481973324, 32'sd0.11946289216572857, 32'sd-0.031540744187548306, 32'sd-0.17199004521736633, 32'sd-0.08029344410234592, 32'sd-0.06526299428383592, 32'sd-0.09978482974232458, 32'sd-0.030533669276503275, 32'sd0.01121818543993894, 32'sd-0.008677684599036875, 32'sd-0.08773061013286203, 32'sd-0.02703480748512799, 32'sd0.022624630873092817, 32'sd0.06809393385915007, 32'sd-0.06173513075676541, 32'sd0.04824283334427561, 32'sd0.0038939442786839846, 32'sd-0.05244916892175724, 32'sd-0.14091955689006996, 32'sd-0.03125619337565902, 32'sd0.09647088868863915, 32'sd0.08455932349210052, 32'sd0.08977447223129682, 32'sd0.0702959825609655, 32'sd0.1908436404050924, 32'sd0.08297221823997912, 32'sd0.2160156463228044, 32'sd0.10897750614514999, 32'sd-0.05409885202463194, 32'sd-0.04542182411309016, 32'sd-0.07282618539601918, 32'sd-0.1688523144531022, 32'sd-0.07856304491114557, 32'sd-0.11331262942081907, 32'sd-0.04871275447109242, 32'sd-0.11205653294475552, 32'sd0.018504034800514033, 32'sd0.1207651654152299, 32'sd-0.016460138065703893, 32'sd-0.08785167560839047, 32'sd-0.043052214816791924, 32'sd-3.6266843151754895e-116, 32'sd-0.059666990805482316, 32'sd0.05073895007993627, 32'sd-0.0997174863997278, 32'sd-0.17200408213429735, 32'sd-0.16013379369268207, 32'sd-0.10057288887959648, 32'sd0.054990850952046, 32'sd0.13197744233318884, 32'sd-0.0004271174017063713, 32'sd0.08040616548444912, 32'sd0.21096813589103486, 32'sd0.15269323893376635, 32'sd0.26641931666053575, 32'sd0.016488202189896394, 32'sd-0.19810403786521125, 32'sd-0.0750040478360336, 32'sd-0.11514144373715036, 32'sd-0.10256398707816354, 32'sd-0.04872806212783579, 32'sd-0.027855067817911753, 32'sd-0.14780632988513617, 32'sd-0.08581930998984144, 32'sd-0.0005490438579531957, 32'sd0.03465028907008961, 32'sd-0.05564367413944743, 32'sd-0.05097273739755898, 32'sd-0.04691189665600499, 32'sd0.0059992326984744685, 32'sd0.03188422414795132, 32'sd-0.024799211941348025, 32'sd0.06864559146527115, 32'sd-0.0014043820045312027, 32'sd-0.07894251206844566, 32'sd-0.08988604856173237, 32'sd0.07576035519655752, 32'sd0.03465522079409935, 32'sd0.004736658244826024, 32'sd0.0632571267552191, 32'sd0.05767135402918541, 32'sd-0.03627915200138697, 32'sd-0.0012745988552608576, 32'sd0.0333939980512305, 32'sd-0.041746273333728955, 32'sd-0.135359757990643, 32'sd-0.02131018105557392, 32'sd-0.07857343312412599, 32'sd-0.12405026608701616, 32'sd-0.033716884744037376, 32'sd-0.08081393229111922, 32'sd-0.04418851036509935, 32'sd0.0040620278486942964, 32'sd-0.02032471558111651, 32'sd0.024518280712995052, 32'sd-0.033429366419086726, 32'sd-0.023068352712948995, 32'sd0.03950357222106527, 32'sd-0.05121933805097875, 32'sd-0.046367754676311, 32'sd0.12237243599029662, 32'sd0.006715421239830637, 32'sd-0.004893706570625611, 32'sd-0.00588080637129939, 32'sd0.10939083905424685, 32'sd0.018766067858705618, 32'sd-0.10335343051109847, 32'sd-0.19797854359030362, 32'sd-0.14457081740783273, 32'sd-0.164185052362483, 32'sd-0.07260945389453025, 32'sd-0.01693013773284803, 32'sd-0.03314885760131955, 32'sd0.12268266485534399, 32'sd0.00045660287960503585, 32'sd0.041133492241552154, 32'sd-0.10221627243622752, 32'sd-0.0711899223098127, 32'sd-0.0535338762924976, 32'sd0.032658994719311406, 32'sd-0.037813580685839426, 32'sd-0.13091799480632818, 32'sd0.008615625353178297, 32'sd-0.103149480187831, 32'sd0.11018570225365674, 32'sd6.59227504498e-125, 32'sd-0.044056443133276064, 32'sd0.06598820526662848, 32'sd0.03666190411715311, 32'sd0.08297907488789272, 32'sd-0.04399680389712281, 32'sd-0.030978104695848302, 32'sd0.05986125346250648, 32'sd0.014044238942532749, 32'sd-0.06827132669264825, 32'sd-0.16092449689993654, 32'sd-0.1014321645493638, 32'sd-0.045651958146519296, 32'sd-0.12101278200097347, 32'sd-0.05994273658052649, 32'sd0.10663350053784791, 32'sd0.03342182098639789, 32'sd0.024196441989750673, 32'sd0.052624965059052994, 32'sd-0.10969852433918312, 32'sd-0.0456446746051493, 32'sd-0.0429611276826009, 32'sd0.0123621134071161, 32'sd-0.08165637905575428, 32'sd0.07013331717060696, 32'sd-0.05882560703068478, 32'sd-0.09786359427355482, 32'sd0.004919469015702021, 32'sd-0.004280031356243403, 32'sd-0.0613206454301819, 32'sd0.09828046522972905, 32'sd0.05363557283744287, 32'sd0.036945065742208544, 32'sd0.08429195261556587, 32'sd0.039816854084872504, 32'sd0.066461222653852, 32'sd0.07765146075755573, 32'sd0.010699515699062856, 32'sd0.06514964518663503, 32'sd-0.12651614023876595, 32'sd-0.12908871180158793, 32'sd-0.10004988090984797, 32'sd-0.0009557291527740634, 32'sd-0.02749199709652616, 32'sd0.10190780010298062, 32'sd-0.04591225742705941, 32'sd0.017490240210148677, 32'sd0.0038907874348203244, 32'sd-0.004433686626109401, 32'sd-0.10002196836562954, 32'sd0.007415832369932844, 32'sd0.04410157737249279, 32'sd-0.015517169088528867, 32'sd-0.015960471982995956, 32'sd-0.05711405760314898, 32'sd-0.03216494981903551, 32'sd-0.014650961334749786, 32'sd-0.04972769277347332, 32'sd-0.05514400389933293, 32'sd-0.059341047789234914, 32'sd0.002116920062382316, 32'sd0.13512592092239537, 32'sd0.06476896586228457, 32'sd0.006440536703002819, 32'sd0.020683052254699935, 32'sd0.03365513828123828, 32'sd-0.017289680664232192, 32'sd-0.05873551628256149, 32'sd-0.13212774923733095, 32'sd-0.06315025793892365, 32'sd-0.15858026073961995, 32'sd-0.06244835314247451, 32'sd-0.048585516099178626, 32'sd-0.04871928805008048, 32'sd-0.06455238156301782, 32'sd-0.12381743742530597, 32'sd-0.05205963181714184, 32'sd-0.09193973211391286, 32'sd-0.06891168712250724, 32'sd0.030689444944642773, 32'sd-0.1100390308239193, 32'sd-0.058039501734881115, 32'sd-0.014224718345951596, 32'sd-0.016209633582214326, 32'sd7.597345755442968e-127, 32'sd-0.01543689509237421, 32'sd-0.04597731950023601, 32'sd-0.09367323124366597, 32'sd-0.017261669423979567, 32'sd0.07184921904329497, 32'sd-0.07241719541412422, 32'sd0.044696864234667975, 32'sd0.08555621106486089, 32'sd0.06351279865577068, 32'sd0.009320402637039406, 32'sd0.09623891315309263, 32'sd-0.02467566212461154, 32'sd-0.009991251150281596, 32'sd-0.10182690463499162, 32'sd-0.059997201939112565, 32'sd-0.03971993360069697, 32'sd-0.09158556221301223, 32'sd0.08605794235632055, 32'sd-4.010130175552351e-05, 32'sd-0.06778231864576847, 32'sd-0.09140649558497356, 32'sd-0.011284433648954605, 32'sd-0.012766911005109833, 32'sd0.06740208359097168, 32'sd-0.033395444223819445, 32'sd0.09178406466323931, 32'sd3.009653020287363e-126, 32'sd-1.2913742068940284e-118, 32'sd-1.2205007330312928e-125, 32'sd0.04843069976692473, 32'sd-0.13753173237766544, 32'sd0.10422854845926656, 32'sd-0.030174459903126123, 32'sd-0.0189907606447374, 32'sd0.05713723077716665, 32'sd-0.05591811063097451, 32'sd-0.012362304123252791, 32'sd-0.010097638357189652, 32'sd-0.04001440328463451, 32'sd-0.0009203109073838921, 32'sd-0.051213523831090985, 32'sd0.021252484741614744, 32'sd-0.07263263460689048, 32'sd0.02470909692332891, 32'sd-0.029627033943153674, 32'sd-0.004178136509147448, 32'sd-0.08042669608038264, 32'sd-0.08673039510001702, 32'sd0.011980471394680782, 32'sd-0.014121288979285374, 32'sd-0.024202701415441105, 32'sd0.10467789768245252, 32'sd-0.060781011495857254, 32'sd-0.041077688307623345, 32'sd-1.5473796733272684e-125, 32'sd1.872444543799359e-125, 32'sd-6.312567177314636e-123, 32'sd-0.03891614880706139, 32'sd-0.015283234515602448, 32'sd0.028455170654188202, 32'sd0.11638953237660604, 32'sd0.029353923767310035, 32'sd0.0968338655776905, 32'sd0.15172437614082662, 32'sd0.0372004307920867, 32'sd0.0633066991053967, 32'sd0.041164336373222754, 32'sd0.005641183515248912, 32'sd0.09118534072126326, 32'sd-0.02632635153170738, 32'sd0.108968315705108, 32'sd0.040130668227875574, 32'sd-0.07259800148201434, 32'sd-0.005382956599909454, 32'sd-0.11396382205475629, 32'sd-0.08454929346030206, 32'sd-0.07023616848276286, 32'sd0.038982702356545565, 32'sd0.010356182800411673, 32'sd-0.1208740478789367, 32'sd-0.008959156070505885, 32'sd-0.02241076491468805, 32'sd-3.1938606341989367e-124, 32'sd-8.40996900753099e-118, 32'sd8.368902284177166e-122, 32'sd-5.806370573976169e-124, 32'sd-0.03477437249926584, 32'sd-0.0020271355930024273, 32'sd0.039703343915062285, 32'sd0.08119240719607897, 32'sd0.1014152026858305, 32'sd0.19724983896911394, 32'sd0.1098848809331976, 32'sd0.08077944011287856, 32'sd0.08891941429534504, 32'sd0.007729597481654063, 32'sd0.06900449341594483, 32'sd0.08942486347156178, 32'sd0.016509567232536368, 32'sd-0.07601143778587309, 32'sd0.016982531179294116, 32'sd-0.007453044999955228, 32'sd0.09392345486824571, 32'sd0.08788229367072212, 32'sd0.07725569527602352, 32'sd-0.030510749472433398, 32'sd-0.07315845944352632, 32'sd0.0632689519262039, 32'sd-0.03309423551601062, 32'sd-4.208373336412398e-126, 32'sd4.299657054711411e-118, 32'sd-8.153663689384324e-119, 32'sd-3.9624918270589774e-116, 32'sd1.618101978941903e-127, 32'sd-1.3439859707353694e-124, 32'sd0.04019144734085993, 32'sd0.06555591102575434, 32'sd0.05152132517256436, 32'sd-0.04041953791332546, 32'sd0.0429606079990597, 32'sd0.008831913117042123, 32'sd-0.11786931376339681, 32'sd-0.013454383185793893, 32'sd0.03880032664546478, 32'sd0.008042285622943991, 32'sd-0.018043100908281116, 32'sd0.08664695795361567, 32'sd0.026224214848284213, 32'sd0.041293343068543854, 32'sd-0.02015631229419508, 32'sd0.06722907200810647, 32'sd-0.02300873180288167, 32'sd-0.04566740226857254, 32'sd-0.02187632305714253, 32'sd-0.020207909852384593, 32'sd-5.270257327900731e-120, 32'sd1.7856623762676613e-125, 32'sd-2.1307206853511303e-122, 32'sd-2.6218361496411605e-116},
        '{32'sd7.951480568497643e-124, 32'sd-7.496696800132359e-115, 32'sd-1.3338598293138386e-117, 32'sd-6.561159008847667e-126, 32'sd1.213415732761292e-123, 32'sd-2.8131778127605322e-126, 32'sd-4.443634993490649e-116, 32'sd9.169506484537946e-125, 32'sd-3.2097953080649026e-122, 32'sd-3.9593707454107465e-121, 32'sd2.1074218852313485e-117, 32'sd-7.175151826078977e-116, 32'sd-0.04699721011176289, 32'sd-0.05949241253479799, 32'sd0.032959309205010626, 32'sd-0.042613698926388784, 32'sd6.786455931522562e-117, 32'sd1.2116331712979907e-124, 32'sd-3.978104434005707e-128, 32'sd-6.833537642450716e-122, 32'sd-8.450104276929571e-121, 32'sd-9.338927485346433e-122, 32'sd8.624270086256126e-127, 32'sd-2.3684751128697893e-119, 32'sd-1.456895083272299e-127, 32'sd-1.7396281979448917e-125, 32'sd1.0925666537345635e-119, 32'sd-3.2695607736802663e-122, 32'sd1.659826671885347e-123, 32'sd-1.5749777039624626e-123, 32'sd2.8224554077554845e-116, 32'sd1.967904458809042e-114, 32'sd0.050912958185010036, 32'sd0.03399667645867993, 32'sd-0.04800139058235043, 32'sd-0.0476828144853508, 32'sd0.05289168223482673, 32'sd-0.134642021009149, 32'sd-0.07432247122757066, 32'sd0.049600902196977395, 32'sd0.07365315078978166, 32'sd0.00887966355020274, 32'sd0.0011355729120245527, 32'sd0.01883892991632663, 32'sd0.05579073212639839, 32'sd-0.011724793963392328, 32'sd0.06697934075812646, 32'sd0.10241099160492728, 32'sd-0.009243942557469213, 32'sd0.07557671571971873, 32'sd0.07880270279081, 32'sd0.005448465232816968, 32'sd1.7191155698149736e-124, 32'sd-9.185738875193651e-121, 32'sd-6.626938774220797e-120, 32'sd-7.371174182660322e-123, 32'sd1.161536835999029e-122, 32'sd-9.941059968592682e-116, 32'sd0.004816471164146988, 32'sd0.08518374648643615, 32'sd0.03166715927176895, 32'sd0.0038304174137357688, 32'sd-0.05902037883088177, 32'sd-0.03555119146999887, 32'sd0.023992621728806344, 32'sd-0.021553224377549373, 32'sd-0.12025743628302993, 32'sd0.029081358958419536, 32'sd0.061012901663004514, 32'sd-0.023959524912510657, 32'sd0.08518653291980018, 32'sd0.12103424588412182, 32'sd0.0063817787334337775, 32'sd0.007121452366020012, 32'sd-0.03963273616967945, 32'sd0.022669396126359927, 32'sd0.06474811312138838, 32'sd-0.022508395630913204, 32'sd0.0978130534122488, 32'sd0.05740724612618707, 32'sd0.049954949793407394, 32'sd0.10387507924842111, 32'sd3.11972984942362e-120, 32'sd-2.5295971674157107e-126, 32'sd-3.8672797423218256e-126, 32'sd8.730586838525166e-123, 32'sd0.02613147634921421, 32'sd-0.014815095911524292, 32'sd0.031710771329576434, 32'sd-0.04993022916587384, 32'sd-0.07274324952174156, 32'sd-0.08950440891627018, 32'sd-0.040414468885036026, 32'sd-0.030675213868629734, 32'sd0.12405331617562783, 32'sd0.07531362407382247, 32'sd0.06136123428704608, 32'sd0.029002920752078765, 32'sd0.15647067620536903, 32'sd0.028931877082304675, 32'sd0.08196377732211173, 32'sd-0.044810443821418335, 32'sd0.03637361813127548, 32'sd-0.018012996191384745, 32'sd0.070913354042114, 32'sd0.049745695531829406, 32'sd-0.0053929519914276, 32'sd0.0075246832177274445, 32'sd-0.026443453992338325, 32'sd0.048153997850643566, 32'sd-0.0042318151236328885, 32'sd-2.5378481740499718e-116, 32'sd4.899736896276494e-126, 32'sd0.0475496146280416, 32'sd0.05714491331824329, 32'sd-0.09056899949198488, 32'sd0.014460163043419003, 32'sd0.0017516642051255446, 32'sd-0.08636173334237256, 32'sd-0.04279476363952975, 32'sd-0.03447200535182039, 32'sd0.09774963930900238, 32'sd0.045283461360830814, 32'sd0.05953309660838091, 32'sd0.021130742171918328, 32'sd-0.014428945546681306, 32'sd0.13971516469360662, 32'sd0.14876993562531918, 32'sd0.05397823078441906, 32'sd0.030296358383424028, 32'sd-0.03707536670552524, 32'sd0.023587150168472834, 32'sd0.07297250139604441, 32'sd0.03306141047321631, 32'sd-0.0016977638513227089, 32'sd-0.08348192527635886, 32'sd-0.041726937601605736, 32'sd-0.053668101297381796, 32'sd-0.010518488757815476, 32'sd0.08961243189396444, 32'sd3.525174352137794e-116, 32'sd0.032208708623652806, 32'sd-0.009410418024289295, 32'sd-0.07086656327177522, 32'sd-0.03998390024056205, 32'sd-0.09585258564322814, 32'sd-0.0630444108614633, 32'sd0.002756762227370647, 32'sd-0.03201151697098146, 32'sd0.016925330728265683, 32'sd0.07111089206268438, 32'sd0.07290864279995878, 32'sd0.09639835858180444, 32'sd0.014047726759231452, 32'sd0.1644524277278519, 32'sd0.049903978787740264, 32'sd-0.03660900534326015, 32'sd0.07495213751679916, 32'sd0.04181429756471406, 32'sd-0.050023691001383284, 32'sd-0.0778416051594684, 32'sd0.003068446229969968, 32'sd0.04139618677515682, 32'sd-0.038305233833278884, 32'sd0.06192924137662796, 32'sd0.06639918156099023, 32'sd0.031098221395060945, 32'sd0.031838433511733114, 32'sd-1.3593300101212308e-117, 32'sd0.031397312464294974, 32'sd0.03610447299164259, 32'sd-0.033972081733865296, 32'sd-0.02183355173382909, 32'sd-0.15646055937539644, 32'sd-0.049200952370889166, 32'sd0.032374537463862214, 32'sd0.006273259858406886, 32'sd-0.0518479441072125, 32'sd0.054114401875082735, 32'sd0.060645559967382565, 32'sd0.07719171898015055, 32'sd0.1260752441522284, 32'sd0.05050485668301635, 32'sd-0.059414110454828965, 32'sd-0.14551248466265604, 32'sd0.05852615708313148, 32'sd-0.029363081577734134, 32'sd0.009613374716671643, 32'sd0.011182963408050512, 32'sd-0.05019441911275445, 32'sd0.1290271453975909, 32'sd-0.026966315329935653, 32'sd0.009203387038324821, 32'sd0.042139576301008216, 32'sd-0.006995040069170878, 32'sd0.03537163898254246, 32'sd0.007949911985790568, 32'sd0.04234298173736934, 32'sd-0.035108974195360895, 32'sd-0.016333283563035716, 32'sd-0.1297557354667411, 32'sd-0.19949271670431076, 32'sd-0.06097490640143803, 32'sd-0.03796552468480152, 32'sd-0.07072115510141251, 32'sd0.06939237468929513, 32'sd0.06771219733008438, 32'sd0.12160620247095504, 32'sd0.025832955178159506, 32'sd0.05183477833582597, 32'sd-0.04909363256648829, 32'sd-0.03213869466803027, 32'sd-0.13103072915554395, 32'sd-0.07426714982361383, 32'sd-0.04097634707032648, 32'sd-0.09572911491933073, 32'sd0.03438807854583756, 32'sd0.11230536588574341, 32'sd0.23284468739117342, 32'sd0.008162253156424548, 32'sd0.005977229390630696, 32'sd0.04191218353091297, 32'sd-0.0678971209438914, 32'sd0.0372893018811647, 32'sd0.018204726498052968, 32'sd0.0784603816432983, 32'sd-0.09857204512077648, 32'sd-0.01770461184208329, 32'sd-0.17300890807099575, 32'sd-0.13574233281764242, 32'sd-0.024598152281523265, 32'sd-0.05227422145418569, 32'sd0.05227189844862631, 32'sd0.06101934870568359, 32'sd0.1062473116992926, 32'sd0.08872323154059644, 32'sd0.03687137046173629, 32'sd0.03627128306020824, 32'sd-0.07331963570568942, 32'sd-0.06561440073563, 32'sd-0.0773224616433935, 32'sd-0.13762669879975034, 32'sd-0.07266657280239837, 32'sd-0.11723817244807803, 32'sd0.004977266143741724, 32'sd-0.0145830132731648, 32'sd0.008789631494973506, 32'sd-0.021996782965619088, 32'sd-0.07309803982014201, 32'sd-0.09576333567194793, 32'sd-0.008555260772971428, 32'sd0.014438297491798901, 32'sd-0.029207537969592263, 32'sd0.002057916943888798, 32'sd0.01596334420104768, 32'sd0.10359294215081896, 32'sd-0.04120098626315115, 32'sd-0.15521806777930866, 32'sd0.07491952931293937, 32'sd0.010956142902560678, 32'sd0.08005458074942264, 32'sd0.09998140809173711, 32'sd0.013899825988347703, 32'sd-0.0325375476791805, 32'sd-0.018779747082919507, 32'sd-0.16812072298227895, 32'sd-0.2239159441542647, 32'sd-0.08889326970785401, 32'sd-0.044406173332894455, 32'sd-0.1352162726547111, 32'sd-0.0979190930498269, 32'sd-0.1588907892295873, 32'sd-0.03347955971776948, 32'sd-0.03519068864118472, 32'sd0.012947827844408852, 32'sd-0.06638974722315302, 32'sd-0.02188542375888095, 32'sd-0.009521325102522274, 32'sd-0.04811496423125869, 32'sd-0.01089708034190337, 32'sd0.005295393639792004, 32'sd0.05825141049667568, 32'sd-0.02282337093055762, 32'sd-0.07086038367495495, 32'sd-0.17518094428970868, 32'sd-0.07843690510464214, 32'sd0.03675512588805589, 32'sd0.10932361536113178, 32'sd0.12558516704864683, 32'sd0.16004504436059466, 32'sd0.03360780574405796, 32'sd-0.15801060786914536, 32'sd-0.024677431708575705, 32'sd-0.1458697003068174, 32'sd-0.19831370153255481, 32'sd-0.12848957036447992, 32'sd0.010858959791430192, 32'sd0.06486459112652479, 32'sd-0.08686732195908717, 32'sd-0.16083024343346047, 32'sd-0.0182483787207983, 32'sd-0.03763941439333572, 32'sd-0.06888633236372019, 32'sd-0.012410684685234001, 32'sd0.14615855844972933, 32'sd0.06376958487158443, 32'sd-0.03931525953223845, 32'sd0.009943841699161968, 32'sd0.01243467467710557, 32'sd-0.011700255203828837, 32'sd0.032763331921769834, 32'sd-0.03026003208856217, 32'sd-0.09778310759443551, 32'sd-0.06175417750883132, 32'sd-0.032923648694110665, 32'sd0.1294247558308647, 32'sd0.1929219163973235, 32'sd0.07420596461779361, 32'sd-0.08655794414324684, 32'sd0.002321890586873696, 32'sd0.13895329349890564, 32'sd0.05115497719418726, 32'sd-0.0987503704633157, 32'sd-0.12191314431645707, 32'sd-0.013615838167921763, 32'sd0.21280198044547716, 32'sd0.04082809681105894, 32'sd-0.0958527259720901, 32'sd-0.15040272110466818, 32'sd-0.12657639810877974, 32'sd-0.07429822995884974, 32'sd0.12264613170070139, 32'sd0.09600405415196968, 32'sd-0.011702164087209742, 32'sd-0.04103129411499532, 32'sd-0.03172734416100207, 32'sd0.018788778763267507, 32'sd-0.03342706943423693, 32'sd0.008274977608055812, 32'sd-0.04833410556041501, 32'sd-0.12483143189786713, 32'sd-0.09404834051039627, 32'sd0.018881478761831168, 32'sd0.006757705858211787, 32'sd0.10546145540414091, 32'sd0.11781934323210608, 32'sd0.004076225414709794, 32'sd0.043528060749653395, 32'sd0.04900750766829282, 32'sd0.13044222989057996, 32'sd-0.03210218341088578, 32'sd-0.08982191906347144, 32'sd-0.038268011092840434, 32'sd0.1273227646676408, 32'sd0.14348707648976222, 32'sd0.034040835581824275, 32'sd-0.09295646372623825, 32'sd-0.09430142995616571, 32'sd-0.1721425264953877, 32'sd-0.060326025506917985, 32'sd0.11705559947281297, 32'sd-0.13182406342769695, 32'sd-0.006582836563390464, 32'sd0.07010168721469813, 32'sd0.006083636742061007, 32'sd-0.0280463925772904, 32'sd-0.023313234549751462, 32'sd-0.07348707985040139, 32'sd-0.2708273396938104, 32'sd-0.19080866163575944, 32'sd0.015154672723153918, 32'sd0.13578121191195539, 32'sd0.08737552654359858, 32'sd0.05238737534023391, 32'sd0.03182058148119841, 32'sd0.06230943559352467, 32'sd0.1284650973626212, 32'sd0.06787459598286333, 32'sd0.13959223468120652, 32'sd0.09299669182084688, 32'sd0.04986990202695491, 32'sd-0.11526722071510409, 32'sd0.05842051625908025, 32'sd0.06530378293100468, 32'sd0.07423707531431724, 32'sd-0.06326353685029244, 32'sd-0.052523753218736535, 32'sd0.04610077876867965, 32'sd-0.0026938991599534867, 32'sd-0.1138721332305799, 32'sd-0.0014691677987096058, 32'sd0.039555913940295694, 32'sd0.09379500442623659, 32'sd-0.016837441779102246, 32'sd0.011519456876198096, 32'sd-0.00340262162136147, 32'sd-0.15990190041830976, 32'sd-0.09004819694827786, 32'sd-0.1057996995967266, 32'sd-0.05108150726028991, 32'sd0.11895219801809753, 32'sd-0.04440088816517602, 32'sd0.010358181505334506, 32'sd0.008454896519603051, 32'sd-0.016205797862423876, 32'sd-0.011445786786897586, 32'sd0.095531334435383, 32'sd0.04875770264557614, 32'sd0.02636185661021532, 32'sd0.07444717639094986, 32'sd0.019420900807773887, 32'sd-0.032347972670960956, 32'sd0.053511652419116075, 32'sd-0.039091433140087194, 32'sd0.07992718281724438, 32'sd0.031423301050865854, 32'sd0.0759304549675668, 32'sd-0.012111175329953866, 32'sd0.03608218438069565, 32'sd-0.024135073203428312, 32'sd0.004963795166362664, 32'sd0.05299402656256147, 32'sd0.10642190828432999, 32'sd0.009386490144851399, 32'sd-0.020725053220369688, 32'sd-0.09359377359682293, 32'sd0.001534654637995585, 32'sd-0.005667954912978105, 32'sd0.07093761527789458, 32'sd0.008216706721628424, 32'sd-0.017456346592910593, 32'sd0.005317926885174995, 32'sd-0.00716490101885092, 32'sd0.02266380912871643, 32'sd0.07525481273669168, 32'sd0.03668991859091673, 32'sd0.037994228928003006, 32'sd0.026737567752387444, 32'sd0.07044094045075923, 32'sd-0.09278851902382661, 32'sd-0.003135177307064778, 32'sd-0.03469843295343324, 32'sd-0.05463342140930234, 32'sd-0.00922726337153667, 32'sd-0.029589597291743115, 32'sd-0.10637505434159628, 32'sd0.05508232507050836, 32'sd0.06014343939907547, 32'sd0.03748701272255449, 32'sd-0.04315722307289305, 32'sd-0.0011083724709577535, 32'sd-0.025284585492391095, 32'sd0.0626184941957767, 32'sd0.009582758226686819, 32'sd-0.06000519448436459, 32'sd0.028486116528948217, 32'sd0.1210079931912485, 32'sd0.07168530450013076, 32'sd-0.061473737573230526, 32'sd0.06926175853956305, 32'sd0.037978521252219795, 32'sd0.1384113668375694, 32'sd0.05747090422076038, 32'sd-0.0038417887310348156, 32'sd0.13821059143142048, 32'sd0.0716920448680895, 32'sd0.09393689804595587, 32'sd-0.05279368800051085, 32'sd-0.13359811419183915, 32'sd-0.08507768914356384, 32'sd-0.09711413282052277, 32'sd0.07493735803593977, 32'sd-0.08838826998516505, 32'sd0.05447382179309683, 32'sd-0.02208375197676996, 32'sd0.0750069265111606, 32'sd-6.377549118106049e-121, 32'sd0.037445401526256826, 32'sd0.08446833854156531, 32'sd-0.10817623520051632, 32'sd-0.00031143605773760187, 32'sd-0.09004662260147217, 32'sd-0.01838802104236537, 32'sd0.004307324934872053, 32'sd-0.09343572846304213, 32'sd-0.05274056163564469, 32'sd0.06421952511215435, 32'sd0.10207195880849551, 32'sd0.17317297321601194, 32'sd0.13268268351869808, 32'sd-0.12114024077739124, 32'sd0.01965970329298619, 32'sd0.1732271831863251, 32'sd0.015665107787260314, 32'sd0.04176507856397524, 32'sd-0.03470196129030101, 32'sd0.04096183165188463, 32'sd0.011248179506857435, 32'sd0.14647222260537843, 32'sd0.04642922453640216, 32'sd-0.020674458636654205, 32'sd0.00844000656648649, 32'sd-0.07000131648755309, 32'sd0.03949503912163502, 32'sd0.008265408377296172, 32'sd-0.02395286759601756, 32'sd-0.015163033215506381, 32'sd-0.0010316723944308799, 32'sd-0.13154561534330036, 32'sd-0.12839207965290791, 32'sd-0.07363459091000338, 32'sd-0.09159757694809995, 32'sd-0.0008216984453080444, 32'sd-0.05759102584403925, 32'sd-0.08285181432156906, 32'sd-0.06738692249034622, 32'sd0.012970971152774145, 32'sd0.08325101064825159, 32'sd-0.13231865042267232, 32'sd-0.07488677769187099, 32'sd-0.05631200829936464, 32'sd0.0013571593426956788, 32'sd0.08668201388250703, 32'sd-0.05531872612803461, 32'sd0.023491334236191007, 32'sd0.007112636666780636, 32'sd0.050334878384691195, 32'sd-0.01830102314869509, 32'sd-0.005662514620088473, 32'sd0.09757411663467425, 32'sd-0.02526591168509778, 32'sd0.0004115822010972066, 32'sd0.015335627867941543, 32'sd-0.008696715285214403, 32'sd-0.018817934762692952, 32'sd-0.018684837308597282, 32'sd-0.1265525812965474, 32'sd-0.14377569077845648, 32'sd-0.049597718557060216, 32'sd-0.11772183197164139, 32'sd0.08686836763106776, 32'sd0.09354164975246108, 32'sd-0.09716125713229577, 32'sd-0.1312729833869844, 32'sd0.2013897287672457, 32'sd0.02853112817397979, 32'sd-0.017478519475552755, 32'sd-0.06390904087241187, 32'sd-0.17296701082510918, 32'sd-0.04011981085765871, 32'sd0.10244971257162297, 32'sd0.03532908753958994, 32'sd-0.029017140932669695, 32'sd0.12703550972190508, 32'sd-0.011548033978362246, 32'sd-0.04361053234163919, 32'sd-0.0597102192295019, 32'sd0.05055192230026045, 32'sd-0.14114251528694385, 32'sd-0.12667471341048045, 32'sd9.313112291832259e-115, 32'sd-0.004052616014550037, 32'sd-0.11883719567516757, 32'sd0.004468258274375596, 32'sd-0.10509931027840604, 32'sd-0.0620393609256116, 32'sd-0.00367539449780048, 32'sd-0.031110516999811134, 32'sd-0.08134035109210806, 32'sd0.0888016477305199, 32'sd-0.08394418205366048, 32'sd-0.0015907826579696753, 32'sd-0.014597338076695568, 32'sd0.09577292783419357, 32'sd-0.008120131878615412, 32'sd-0.023163926033227235, 32'sd-0.11102337812910404, 32'sd-0.07096646296073944, 32'sd0.048891695520403095, 32'sd0.0401869267588305, 32'sd0.07410760687367475, 32'sd0.10241248204706678, 32'sd0.09413617602683755, 32'sd-0.0923857054567332, 32'sd-0.13066548165072733, 32'sd0.007507457559109396, 32'sd-0.014250059864498364, 32'sd0.053648411310123274, 32'sd0.03274441460261553, 32'sd-0.04190857394591446, 32'sd-0.01871600530047864, 32'sd-0.006400040241372868, 32'sd0.05768909529230481, 32'sd0.06320725100553119, 32'sd0.02919151298522017, 32'sd-0.031981479221276254, 32'sd0.0911188609842065, 32'sd0.028902984479427875, 32'sd0.02468293179498251, 32'sd-0.022355808514266926, 32'sd0.05724979458986449, 32'sd-0.018563912406389632, 32'sd0.05744059055003146, 32'sd-0.016511263599040187, 32'sd-0.032871167156505225, 32'sd0.11442479182030746, 32'sd0.11274111858618908, 32'sd0.12751977255273236, 32'sd0.04909017316201662, 32'sd0.08144312386605171, 32'sd0.018895337389803857, 32'sd0.010842533906128028, 32'sd-0.0070988703912748365, 32'sd-0.06910580634239165, 32'sd-0.05668867107318295, 32'sd0.032554113641520596, 32'sd0.06754811418274238, 32'sd0.0964899227535734, 32'sd0.027320072557608283, 32'sd-0.12060940628235478, 32'sd-0.04310206598336428, 32'sd0.0005995258333163932, 32'sd-0.03355582648289609, 32'sd-0.06968011039777806, 32'sd-0.033796736635131164, 32'sd0.01930206996764073, 32'sd0.015711354025782578, 32'sd0.02620943862371007, 32'sd-0.11894633955402142, 32'sd-0.07879222388942088, 32'sd-0.0348850055927524, 32'sd0.05529315071622706, 32'sd0.026304365313763657, 32'sd0.10492023214513828, 32'sd0.08752669426144999, 32'sd0.08153102870439904, 32'sd-0.0485755701801372, 32'sd-0.11648590365954434, 32'sd-0.05730965085885273, 32'sd-0.011684449997492739, 32'sd-0.05640376679205307, 32'sd0.03076099589434014, 32'sd-0.1073601348100815, 32'sd0.04348895179811615, 32'sd-2.851026857541417e-121, 32'sd0.04721294730417495, 32'sd-0.08019044483176416, 32'sd0.03902893275625289, 32'sd0.0735521896019602, 32'sd0.07867345978889598, 32'sd-0.035174434733633526, 32'sd-0.08573443159923819, 32'sd0.1112012318651817, 32'sd-0.050813776388468394, 32'sd0.013077600336623104, 32'sd0.0050283548509912675, 32'sd0.014954144791118456, 32'sd-0.07225762225501266, 32'sd0.072630388231452, 32'sd0.0733048828632842, 32'sd0.06213480830883372, 32'sd0.1655161873967757, 32'sd-0.028675582671103383, 32'sd0.018202190066657017, 32'sd-0.0057326048027626355, 32'sd-0.16897580823086863, 32'sd0.0019300579855226964, 32'sd-0.01474631863523343, 32'sd0.04745864512705386, 32'sd-0.06718179568825552, 32'sd-0.0012039433649351672, 32'sd1.3126664712432105e-122, 32'sd8.719029468866408e-117, 32'sd-1.712432263390698e-127, 32'sd0.042817919987254024, 32'sd-0.08519407662156436, 32'sd-0.039292537047350924, 32'sd0.01953405136937066, 32'sd-0.06551783252193412, 32'sd0.017773170119530595, 32'sd0.0043374228350812, 32'sd0.052553175597701576, 32'sd-0.0939571474567731, 32'sd-0.06862361548963018, 32'sd0.06943123551712214, 32'sd0.11651894335795233, 32'sd-0.0022404439167103157, 32'sd0.09241266133229704, 32'sd0.18046541797858773, 32'sd-0.05523802086116331, 32'sd-0.09199460999468641, 32'sd-0.001636259630189841, 32'sd0.04871674686806118, 32'sd-0.07322479789620588, 32'sd-0.04292122035774182, 32'sd0.027847201362976755, 32'sd0.05289067888599446, 32'sd0.04028949179383756, 32'sd0.07762349798936838, 32'sd1.5799102434226868e-125, 32'sd8.412882805568751e-123, 32'sd-2.6143511596252806e-126, 32'sd-0.001685139812149529, 32'sd-0.006897179958728646, 32'sd0.053941519732036536, 32'sd-0.006426174618081209, 32'sd0.00035688361666186486, 32'sd-0.013655730081668255, 32'sd0.009552980323341703, 32'sd-0.03028240431190945, 32'sd0.07212021471526106, 32'sd0.0970148732412929, 32'sd0.15978228851096438, 32'sd0.04591324828329149, 32'sd0.04597613733558488, 32'sd0.10124658815163387, 32'sd0.04417985959255512, 32'sd0.08884182767115689, 32'sd0.16424158910838166, 32'sd0.04945640874076981, 32'sd0.0876693677461893, 32'sd0.09613568970565102, 32'sd0.010159474324570683, 32'sd0.08334543262745647, 32'sd0.08989199943995714, 32'sd0.05799447990564636, 32'sd-0.06770656308701944, 32'sd-1.1427882799847157e-122, 32'sd2.2581807053148297e-118, 32'sd3.9935939615558666e-121, 32'sd2.323518528112311e-117, 32'sd0.0722799088587055, 32'sd0.0317582060969739, 32'sd-0.08268636333824647, 32'sd-0.07354034026239227, 32'sd0.03050091252120547, 32'sd0.02175387197975402, 32'sd-0.028171698061666514, 32'sd-0.02006819521334369, 32'sd0.02379135261440472, 32'sd0.04519046793971783, 32'sd0.013512907936711506, 32'sd0.010893526229549847, 32'sd0.036759891738908354, 32'sd-0.03057736588750667, 32'sd0.0952069561780798, 32'sd0.017319659365850244, 32'sd0.03406971310164506, 32'sd0.030920349095978687, 32'sd0.004806534195424166, 32'sd0.06062169208845125, 32'sd0.12201049199389086, 32'sd0.02364460168966619, 32'sd0.03408506764546855, 32'sd-1.5119280871478733e-122, 32'sd-9.141888545602273e-127, 32'sd1.709014739628183e-123, 32'sd-1.9647911589408943e-119, 32'sd8.721476189812874e-127, 32'sd4.552449761547482e-126, 32'sd0.013547916157042216, 32'sd0.015048085910463771, 32'sd0.06773835186979872, 32'sd0.01192327512850726, 32'sd-0.011007934590312072, 32'sd-0.01775882771581719, 32'sd-0.010977101140209942, 32'sd-0.011063202677253489, 32'sd0.01002284812197597, 32'sd0.044222657842817543, 32'sd0.06304420869708006, 32'sd0.07336843938917417, 32'sd0.012032383623086272, 32'sd-0.08010785084268603, 32'sd0.06638916598292424, 32'sd0.03282228901506244, 32'sd0.029735107287167828, 32'sd-0.11379526476107282, 32'sd-0.008993629820362245, 32'sd-0.0009512141149772196, 32'sd-6.369154272768971e-116, 32'sd3.8316124056348255e-115, 32'sd-6.375726641059043e-125, 32'sd-4.221528825889207e-121},
        '{32'sd-6.493087792485083e-125, 32'sd-3.961101767673277e-116, 32'sd-6.790328242952538e-124, 32'sd-1.9975787720541944e-127, 32'sd-3.370208635412704e-120, 32'sd1.8480835054965913e-116, 32'sd-2.5505749080655532e-124, 32'sd6.383580199239049e-127, 32'sd-4.3483137773107063e-126, 32'sd-1.3309015751157765e-118, 32'sd4.514913582502383e-115, 32'sd-2.42459123538884e-124, 32'sd0.007335138532554862, 32'sd-0.029367445746014843, 32'sd0.010866999360834113, 32'sd0.024699740637656346, 32'sd-4.2973111974275903e-125, 32'sd-9.490518549804363e-124, 32'sd2.7207050098534142e-121, 32'sd-1.0715739021364708e-124, 32'sd5.298735483851802e-118, 32'sd4.173319919918554e-123, 32'sd7.786153085496978e-125, 32'sd7.499990308445732e-126, 32'sd4.412623114162358e-124, 32'sd-2.4721423274452384e-122, 32'sd-1.3093669275762834e-122, 32'sd3.7605962448670677e-119, 32'sd6.847911925267463e-127, 32'sd8.891922553309799e-118, 32'sd3.999394553172594e-116, 32'sd3.61800995763763e-123, 32'sd0.062043373144264946, 32'sd0.08979747948449668, 32'sd-0.059851245182860925, 32'sd-0.04740084448694345, 32'sd-0.033249863852085615, 32'sd-0.08337687950555057, 32'sd0.03219698430840754, 32'sd-0.052122993627396016, 32'sd0.01545279827055107, 32'sd0.0024755552011334753, 32'sd0.05028627050078777, 32'sd-0.0435639970555317, 32'sd0.03956585503581318, 32'sd0.11555300847356087, 32'sd0.027300799285322818, 32'sd0.09282123086553687, 32'sd0.0029745312245145436, 32'sd0.08389797441223397, 32'sd0.09331473602093622, 32'sd0.061558548199060564, 32'sd8.200790754555507e-126, 32'sd1.1847984767069102e-125, 32'sd-4.1968217546857207e-125, 32'sd-5.133376136732138e-118, 32'sd2.5616477340302855e-126, 32'sd-1.0100962860929115e-121, 32'sd0.041323517302932496, 32'sd0.0718683424213455, 32'sd0.05330761041017453, 32'sd-0.01929812398601317, 32'sd-0.03298538027830834, 32'sd-0.006961708705144075, 32'sd-0.024778295326527852, 32'sd-0.07017677502920013, 32'sd0.021926652402154537, 32'sd-0.06120672026132114, 32'sd-0.012776088710351973, 32'sd0.1367675999678685, 32'sd0.0461852161109213, 32'sd0.015913619462113678, 32'sd0.03560789557250952, 32'sd0.09259139924765002, 32'sd0.09874341694303465, 32'sd0.1382918832114097, 32'sd0.04450936303501338, 32'sd0.013973892193836756, 32'sd0.09039847087325865, 32'sd0.01180222023144098, 32'sd0.024662338835963842, 32'sd0.10578263021755664, 32'sd4.1075318547307477e-125, 32'sd-9.399592449130122e-122, 32'sd1.0267872238644813e-122, 32'sd6.771189756608094e-122, 32'sd0.1154900249375703, 32'sd0.050066364769620154, 32'sd0.006386445519105098, 32'sd-0.07559887670368073, 32'sd0.007190260687568994, 32'sd-0.05076178146332665, 32'sd-0.13325089475615073, 32'sd0.034105410195425276, 32'sd0.0973853918267733, 32'sd-0.20109284034285457, 32'sd-0.05515353299972287, 32'sd0.016505943233415518, 32'sd0.019684780323563106, 32'sd-0.03720660868170014, 32'sd0.10442801974092109, 32'sd0.13922317138289036, 32'sd0.21478368964405517, 32'sd0.059866199313874616, 32'sd0.12854317754982408, 32'sd0.07461836313460478, 32'sd-0.02000449452382098, 32'sd-0.001251604015312811, 32'sd-0.0006625834049079331, 32'sd-0.019932954669756142, 32'sd-0.03261866228745993, 32'sd6.312562643032702e-126, 32'sd1.5111188951565246e-121, 32'sd0.040684885359340346, 32'sd0.03588466071700186, 32'sd-0.05473727414709999, 32'sd-0.038712919755839785, 32'sd-0.03161760687188435, 32'sd-0.07515626672553963, 32'sd0.024190606603304424, 32'sd-0.09563117799551463, 32'sd0.07827764131047726, 32'sd-0.06431300161640074, 32'sd-0.16705357584069963, 32'sd0.022403780905424345, 32'sd0.020390582432973665, 32'sd0.01239653832394506, 32'sd0.0898625111328079, 32'sd0.004875099798780456, 32'sd0.04524619018274828, 32'sd0.04822910616930803, 32'sd-0.026315841884597856, 32'sd0.024206883844594757, 32'sd0.16766821750605118, 32'sd0.029756576492368483, 32'sd0.052984576832213894, 32'sd-0.035827450003904186, 32'sd-0.021444769714544662, 32'sd0.053406339165541765, 32'sd0.05579446419126936, 32'sd1.5269374995122015e-126, 32'sd0.059906297971557054, 32'sd-0.07769801700083016, 32'sd0.011758939465312873, 32'sd0.009197187157036593, 32'sd-0.006497986397218972, 32'sd-0.00406780906976896, 32'sd0.04898759490708287, 32'sd0.10123265884464272, 32'sd-0.05900481410920008, 32'sd-0.07871485390705324, 32'sd-0.02079306583225515, 32'sd-0.1335399984805254, 32'sd-0.08700922424919384, 32'sd-0.045439355409008224, 32'sd0.05989372189680716, 32'sd0.03754175616550884, 32'sd0.08485094045075581, 32'sd0.1612993607860951, 32'sd0.004419854510189609, 32'sd0.09437441477605192, 32'sd-0.007708165047448934, 32'sd0.06850385393051392, 32'sd0.08634471146442149, 32'sd-0.06595949750653866, 32'sd0.042802782109903334, 32'sd-0.03096050229299073, 32'sd0.003414246501174338, 32'sd-3.442719269941849e-123, 32'sd0.012392375671188992, 32'sd0.04753023380827657, 32'sd-0.01513241963393372, 32'sd-0.07429953625060584, 32'sd-0.010381756496382993, 32'sd0.05886794035791326, 32'sd0.09010545902660302, 32'sd0.05046594459030591, 32'sd-0.0008829768392897669, 32'sd0.01576400850713696, 32'sd0.08974692999207419, 32'sd0.13297531900090806, 32'sd0.09889253196283244, 32'sd0.11723184692559882, 32'sd0.07831116809371284, 32'sd0.16834625823953822, 32'sd0.19353392228164268, 32'sd0.12875393085648, 32'sd0.20280575962854583, 32'sd0.06903073670371535, 32'sd0.07289048530872322, 32'sd-0.04065083690467208, 32'sd0.061677448340188415, 32'sd0.07803655624541372, 32'sd0.12980255851582087, 32'sd0.03429172157034083, 32'sd0.030564616027656876, 32'sd0.10726970726211454, 32'sd0.040748912619586186, 32'sd0.03694087909474937, 32'sd0.009147982350805888, 32'sd0.026702979000890862, 32'sd0.025287921919900456, 32'sd0.011299933194364753, 32'sd0.108426883702189, 32'sd0.026809201912159207, 32'sd0.03844335237213088, 32'sd0.06324541684884533, 32'sd0.004057679502125221, 32'sd0.015129427774043453, 32'sd0.08192689441238786, 32'sd0.05340064384799065, 32'sd0.04774437983395455, 32'sd0.13869235059195528, 32'sd0.16684545547411916, 32'sd0.21633191688073594, 32'sd0.08616367446463062, 32'sd0.16954982013807066, 32'sd0.010850906106764266, 32'sd0.05522003510272272, 32'sd0.1302166339242919, 32'sd0.06070396219404528, 32'sd0.09284408731867677, 32'sd0.048985518780106006, 32'sd0.02422572916894061, 32'sd0.0444285090703932, 32'sd0.1038869939913046, 32'sd0.08005712999021652, 32'sd-0.07997856251690588, 32'sd-0.07724697985056171, 32'sd-0.02773927119846711, 32'sd0.015556002606137808, 32'sd0.156901387275394, 32'sd-0.06753802103163563, 32'sd0.12083242829620806, 32'sd0.09338315111983693, 32'sd0.027743880468684992, 32'sd-0.038745020232500205, 32'sd-0.0003275759322160126, 32'sd0.002901862724045861, 32'sd0.07007002091282818, 32'sd0.0518790751400547, 32'sd0.0390462037461112, 32'sd0.014807080960648453, 32'sd-0.14840132349497875, 32'sd0.003725548642903451, 32'sd-0.08415159318577999, 32'sd-0.09920287406658876, 32'sd0.06750387227965436, 32'sd0.004255784716711679, 32'sd-0.10985826227493198, 32'sd0.010341604132038185, 32'sd-0.009846141802335083, 32'sd0.028075995581061025, 32'sd0.06331603420445862, 32'sd-0.09911786209997608, 32'sd-0.021483120572965544, 32'sd0.05156711961047145, 32'sd-0.0668804331371098, 32'sd0.13237267478188627, 32'sd0.02954963646997873, 32'sd-0.04221404133259947, 32'sd0.009265896420711288, 32'sd0.14258197721528013, 32'sd0.09169648423193548, 32'sd0.050109598198255334, 32'sd0.06612237488317177, 32'sd0.04084972867111832, 32'sd-0.02324109365402641, 32'sd-0.2918382802578361, 32'sd-0.18805192008685942, 32'sd-0.21101856771822283, 32'sd-0.21589647858533456, 32'sd-0.19174988705897109, 32'sd-0.14549501426222095, 32'sd-0.12851193433776245, 32'sd-0.10048869672821219, 32'sd0.0764432799896076, 32'sd-0.04575292092681493, 32'sd0.03866493984351102, 32'sd-0.00716461945513464, 32'sd0.1081109537885842, 32'sd0.05810090587375204, 32'sd0.022165830772946628, 32'sd-0.07318910000377596, 32'sd0.04806642919964506, 32'sd0.04604192007326173, 32'sd0.11949420048441341, 32'sd-0.03884777245222242, 32'sd0.08458737589438287, 32'sd-0.016654384626364163, 32'sd0.18051451549169475, 32'sd0.07250572389439025, 32'sd0.07246026749619613, 32'sd0.04394180750633967, 32'sd-0.11922108856509439, 32'sd-0.12969889963808884, 32'sd-0.1171408234495282, 32'sd-0.21573486451921828, 32'sd-0.11501970319417336, 32'sd-0.2180619200048384, 32'sd-0.29431850815715954, 32'sd-0.2325054292478877, 32'sd-0.12859800964149032, 32'sd-0.09130398956845148, 32'sd-0.12270868440104588, 32'sd-0.10237742183528242, 32'sd0.012905736468431458, 32'sd0.01230850761313208, 32'sd0.07864410226360974, 32'sd-0.006809628108373036, 32'sd-0.03316232671001673, 32'sd0.045338923883044474, 32'sd0.01261767479594146, 32'sd0.09167527558880754, 32'sd0.08764207906575704, 32'sd0.002920991315310017, 32'sd-0.07311195977322303, 32'sd-0.05478472662861158, 32'sd-0.038382582213776405, 32'sd-0.014731626757142445, 32'sd-0.12298274335159662, 32'sd-0.196580056672779, 32'sd-0.13952303785820688, 32'sd0.05544186864786843, 32'sd0.04659068254522525, 32'sd0.007653932561010238, 32'sd-0.04064651033423475, 32'sd-0.18149323739841783, 32'sd-0.2137142887095671, 32'sd-0.19846009071864318, 32'sd-0.03810994955730654, 32'sd-0.0725315571668538, 32'sd-0.12307164577811432, 32'sd-0.0372375055204179, 32'sd0.04112006138525235, 32'sd-0.071300184316642, 32'sd0.019683803732450544, 32'sd-0.06429656961507399, 32'sd-0.006892913917956416, 32'sd0.0935368442749679, 32'sd0.09381946413063665, 32'sd0.04115088017271314, 32'sd0.021196397068539027, 32'sd0.01606388087494868, 32'sd0.06619969106283301, 32'sd0.05599943710258065, 32'sd0.031319300461874526, 32'sd-0.03501518612182174, 32'sd-0.0951303593980122, 32'sd-0.065697077098009, 32'sd-0.008852255295961174, 32'sd0.0737183087594638, 32'sd0.07162713769756489, 32'sd0.07712868122019767, 32'sd0.08527718331132081, 32'sd-0.04521229646389257, 32'sd-0.08388278843518557, 32'sd-0.16915602316128073, 32'sd-0.006494843441845131, 32'sd-0.14897771428011017, 32'sd-0.010631558929900727, 32'sd-0.08254555154849724, 32'sd0.057227038315254115, 32'sd-0.03968515628380144, 32'sd0.043233039114294484, 32'sd0.07946967560300656, 32'sd-0.014525708743472846, 32'sd0.05468636236634658, 32'sd0.10352652662262071, 32'sd0.06406490249357558, 32'sd-0.022265765617981454, 32'sd-0.025244386163816798, 32'sd0.025573158019413365, 32'sd-0.15524014200427844, 32'sd-0.14572797727283987, 32'sd-0.04944928331538467, 32'sd-0.13103534420835486, 32'sd-0.12241304938211674, 32'sd-0.054296837639642104, 32'sd-0.012979680188771546, 32'sd0.05816454015105673, 32'sd0.0829385327461548, 32'sd0.002083043631845101, 32'sd0.07091737229030161, 32'sd-0.09427305102758836, 32'sd-0.04370667056088281, 32'sd0.023421697731515013, 32'sd-0.04925382977874861, 32'sd-0.08870997256043817, 32'sd-0.059112765472862046, 32'sd0.06215606280976574, 32'sd0.028712498276486798, 32'sd0.05183698729089646, 32'sd-0.043568705237439, 32'sd0.011796999435318744, 32'sd0.025940005446892296, 32'sd-0.007600180954574685, 32'sd0.0408395957499871, 32'sd-0.04820589138253486, 32'sd-0.0988230654661825, 32'sd-0.05880301435821096, 32'sd-0.14321525664910037, 32'sd-0.07084115768438647, 32'sd-0.10292660877441487, 32'sd-0.12287439357138105, 32'sd-0.06572500739410288, 32'sd-0.079740046447117, 32'sd0.14762360469823368, 32'sd0.23693566247251163, 32'sd-0.009163884765164946, 32'sd-0.04586630492669293, 32'sd0.06063080137310737, 32'sd0.06215920002491232, 32'sd0.035747655245318824, 32'sd0.008545668223623541, 32'sd0.007999781299016994, 32'sd-0.006414775312658779, 32'sd-0.04737880041585646, 32'sd-0.017684919261227096, 32'sd0.0021854503904781097, 32'sd0.1094428714552145, 32'sd0.030693899828740753, 32'sd-0.02252254560708388, 32'sd-0.013587073223739709, 32'sd-0.03397065325053534, 32'sd0.07055898907090301, 32'sd-0.03688831511620139, 32'sd-0.15278840962288748, 32'sd-0.03962397082245575, 32'sd-0.032311621838129606, 32'sd0.032519592402703766, 32'sd-0.15067142779188725, 32'sd-0.12400266766386668, 32'sd-0.11943568490237069, 32'sd0.04571996778912806, 32'sd0.18628551491912643, 32'sd0.17742181768818122, 32'sd0.08183806565517339, 32'sd0.03874942600448342, 32'sd0.06908476343580351, 32'sd-0.011836512319077444, 32'sd0.011617480248907073, 32'sd-0.010752959819916844, 32'sd-0.08266856130929622, 32'sd-0.05498310509123007, 32'sd-0.0891307529738242, 32'sd0.009683271684248125, 32'sd0.062380297026878084, 32'sd0.07005455242158998, 32'sd0.04005403368278065, 32'sd0.0224827012978647, 32'sd0.04545093223261373, 32'sd-0.0702727144258449, 32'sd-0.06455378047286378, 32'sd0.01762398806180572, 32'sd-0.026146031993854377, 32'sd-0.06386471209022354, 32'sd-0.015391104678781232, 32'sd0.030422306189510754, 32'sd0.019695504589645394, 32'sd-0.0376080351224182, 32'sd-0.025113831613979166, 32'sd0.1529841619099326, 32'sd0.32048684086317497, 32'sd0.16459267385277668, 32'sd0.08686653690664807, 32'sd-0.009368034234685184, 32'sd0.12729988739519282, 32'sd0.04856070501330379, 32'sd0.13210208727788966, 32'sd-0.03454096755202443, 32'sd0.02057050417470819, 32'sd0.09392161936060985, 32'sd0.04194142291178281, 32'sd-0.011292232303306296, 32'sd0.06626453664062422, 32'sd1.3664145951081222e-122, 32'sd-0.0050658017475345846, 32'sd0.08276415311815775, 32'sd0.08465263882049887, 32'sd-0.02787475908536459, 32'sd-0.08495498291921655, 32'sd0.07332497269819628, 32'sd-0.003947474652273648, 32'sd0.1571829307276412, 32'sd0.08038747443559836, 32'sd-0.028107751723925944, 32'sd-0.06488611739115704, 32'sd-0.05835758868005208, 32'sd-0.0645009247566886, 32'sd0.15533583733067746, 32'sd0.24015435726684872, 32'sd0.157456401280759, 32'sd0.10062038852579712, 32'sd0.045599957345631006, 32'sd0.015197859893187603, 32'sd0.1523118060265033, 32'sd0.036051924728775546, 32'sd-0.04264593781252217, 32'sd0.038723928588547576, 32'sd0.10007532004698026, 32'sd0.014343474848628503, 32'sd0.10189261163152112, 32'sd0.03504101013908704, 32'sd-0.006616818111950431, 32'sd0.032095235064407555, 32'sd0.08540249026985694, 32'sd0.024385442911135827, 32'sd0.01320071986824426, 32'sd-0.06683222132822424, 32'sd0.0640538027013167, 32'sd0.008168847758711314, 32'sd0.06410431614753292, 32'sd-0.0078766627293477, 32'sd-0.09972132802416747, 32'sd-0.12240654175691261, 32'sd-0.28918839816083197, 32'sd-0.12807005849478623, 32'sd0.11647362869334993, 32'sd0.20581128493775286, 32'sd0.18798074391321185, 32'sd-0.019637004115942148, 32'sd-0.08510682302172108, 32'sd0.06528263353344194, 32'sd0.003840301660434388, 32'sd0.009962286423175945, 32'sd0.06772621126404851, 32'sd0.05072392812364879, 32'sd0.03161892248083745, 32'sd0.031634755971436224, 32'sd-0.05048097900392913, 32'sd-0.029397198033596042, 32'sd0.08724664155181726, 32'sd-0.006831177130381051, 32'sd0.043548548018416615, 32'sd0.0319084801446302, 32'sd0.07445384087367558, 32'sd-0.0002579174816148594, 32'sd-0.12039170333895455, 32'sd-0.04836934440173076, 32'sd-0.04526111116637134, 32'sd0.0076078194558283916, 32'sd-0.15894968112254215, 32'sd-0.10342335896100135, 32'sd-0.14877588940214728, 32'sd-0.09973793107152755, 32'sd0.15078041902179512, 32'sd0.1392648724641336, 32'sd0.13744152884746863, 32'sd-0.0323011904111778, 32'sd0.06358998225339291, 32'sd-0.028003569678679775, 32'sd0.07298427895172395, 32'sd0.06528506458415854, 32'sd0.06330728163273053, 32'sd-0.022669489714722962, 32'sd0.11512489368696609, 32'sd0.03271850887332052, 32'sd0.0012237345757751385, 32'sd-0.1231092038776458, 32'sd-9.253275791493011e-123, 32'sd0.0505772474774483, 32'sd0.08696835502312321, 32'sd-0.006130047855145, 32'sd0.08092008992143188, 32'sd0.05918783865649363, 32'sd0.02043867340398795, 32'sd-0.06576199063443433, 32'sd-0.07560069257197446, 32'sd-0.05586957088384621, 32'sd-0.09689072971487137, 32'sd-0.11141067702854317, 32'sd-0.09732593969741905, 32'sd0.046940463162536035, 32'sd0.08516519034022113, 32'sd0.09755026970976961, 32'sd0.19766545453101173, 32'sd0.13166783718025596, 32'sd0.22802519652437864, 32'sd0.021541749074221933, 32'sd0.03846322287971793, 32'sd0.0740872503719077, 32'sd0.08090761894192729, 32'sd0.03361209793702717, 32'sd0.07740828462024253, 32'sd-0.09522659297445851, 32'sd-0.09246244935921732, 32'sd0.0774415546949319, 32'sd0.07272951866039166, 32'sd-0.03594240087372379, 32'sd0.026836319452518544, 32'sd0.07881876504005202, 32'sd0.11958501514437976, 32'sd0.07994789090495574, 32'sd0.02721907339266351, 32'sd-0.014056696999519573, 32'sd0.026324494837694636, 32'sd0.06600404011879865, 32'sd-0.033293586941611504, 32'sd0.009242069803008927, 32'sd0.07649624542051381, 32'sd0.06079386854802619, 32'sd0.12060820211889735, 32'sd0.09076643036439895, 32'sd0.1452627181780103, 32'sd0.10936868681824957, 32'sd0.12851221238267432, 32'sd0.017425055965182623, 32'sd-0.0270839124443754, 32'sd0.06521546674406639, 32'sd0.07606928082592442, 32'sd-0.03233914288726614, 32'sd0.06185649745017792, 32'sd0.031002871476947958, 32'sd0.03987268230974956, 32'sd-0.003553830148623945, 32'sd0.045183193467456244, 32'sd-0.000408816884423336, 32'sd-0.03791929820273572, 32'sd-0.041951358853551585, 32'sd0.13220391483735422, 32'sd-0.031493164244541266, 32'sd-0.11654581741081642, 32'sd0.05417487101585433, 32'sd-0.014300355124415645, 32'sd0.055959420656724566, 32'sd0.03990961574381319, 32'sd0.029842495733002412, 32'sd0.0022737562256513882, 32'sd0.02163048358678657, 32'sd0.1968580679318962, 32'sd0.19292744127750944, 32'sd0.03546424495366296, 32'sd-0.015043687667642575, 32'sd0.028213696320755658, 32'sd0.01095595346562697, 32'sd0.0033636045605902197, 32'sd-0.09195434877884019, 32'sd-0.18760034646020432, 32'sd0.0239850780644702, 32'sd-0.005049293618747524, 32'sd0.03851807692882066, 32'sd-0.10736645881054903, 32'sd0.023904234826189596, 32'sd-7.474361580445115e-127, 32'sd0.06353960041159926, 32'sd-0.0564775720119613, 32'sd0.02662683355049002, 32'sd-0.03381289446335978, 32'sd-0.06352566113742081, 32'sd-0.07247266004799051, 32'sd0.049810323380966144, 32'sd-0.06301179411164555, 32'sd0.027110707376060583, 32'sd0.07050634355941639, 32'sd-0.11812818941526654, 32'sd0.02636400629250126, 32'sd0.08397303898158925, 32'sd0.1241720192210926, 32'sd0.11743734181181581, 32'sd-0.06128525487049164, 32'sd-0.012844213688202518, 32'sd-0.16807881762496726, 32'sd0.035599878055722844, 32'sd-0.08604370802921739, 32'sd-0.21626797254114807, 32'sd-0.19955566866170033, 32'sd-0.08457545916288313, 32'sd-0.18948205548746314, 32'sd-0.10307728538731424, 32'sd-0.020128648197377863, 32'sd-6.413114591791615e-115, 32'sd1.3783228481208913e-117, 32'sd6.249598787189899e-117, 32'sd-0.02423192006562919, 32'sd0.0019093978831668205, 32'sd-0.0031239979657852472, 32'sd0.009627705915306114, 32'sd0.035802805147927184, 32'sd0.007661528051036281, 32'sd0.020335317656601144, 32'sd0.03698562276187474, 32'sd-0.06744667452146251, 32'sd0.008513515486524409, 32'sd0.05551270941774317, 32'sd-0.05226642680855727, 32'sd0.07708988023392935, 32'sd0.004680813908520283, 32'sd-0.09024103610798102, 32'sd0.02721025548313098, 32'sd-0.08010165226250046, 32'sd-0.02309397331996343, 32'sd-0.05913704614617507, 32'sd-0.04907784878896156, 32'sd-0.0006173804275059815, 32'sd0.0025983961587112553, 32'sd0.08304277230630912, 32'sd0.10318658100171979, 32'sd0.04444481589214551, 32'sd-1.1051663989456805e-115, 32'sd7.941865063895199e-125, 32'sd-1.8646061432751288e-127, 32'sd-0.00251374105494629, 32'sd0.021716291539738444, 32'sd-0.04394798233964257, 32'sd0.03200142830056731, 32'sd0.021108379114987467, 32'sd-0.08446668687268404, 32'sd-0.09738709081309173, 32'sd0.053732402205482116, 32'sd-0.04885248886265974, 32'sd-0.010925274973472187, 32'sd0.08294903117051682, 32'sd0.15681816997894263, 32'sd0.14523859743182116, 32'sd0.07770820482539169, 32'sd-0.06671410130804907, 32'sd-0.09206035351844974, 32'sd0.0047967640750663796, 32'sd0.022275925797453265, 32'sd0.004412367269323645, 32'sd0.08333717422232154, 32'sd-0.05697290727589632, 32'sd-0.04319403271775142, 32'sd0.058521433552765414, 32'sd0.06817908846140966, 32'sd0.033767750930470505, 32'sd4.6967650011277107e-122, 32'sd1.947021705459326e-114, 32'sd-1.0388814344418434e-123, 32'sd-5.785337557378575e-117, 32'sd0.03949960861841092, 32'sd0.05775725495717523, 32'sd-0.04208536267413089, 32'sd0.1715822501514802, 32'sd-0.03195702212812031, 32'sd-0.03816591567548035, 32'sd-0.03972770332825019, 32'sd-0.010637426327671062, 32'sd0.01558839916720182, 32'sd-0.11855871949106163, 32'sd0.012020526748212001, 32'sd-0.01138558370903831, 32'sd-0.025456321603756722, 32'sd0.09513278168393123, 32'sd-0.04502661925851864, 32'sd0.053177349146349535, 32'sd0.04403808896397979, 32'sd0.06670035115664733, 32'sd-0.0897473537970527, 32'sd-0.023104040229843484, 32'sd-0.0557678065883464, 32'sd0.0852068173358663, 32'sd0.08444608952116346, 32'sd-7.643295666228347e-127, 32'sd-1.3215942444882272e-122, 32'sd1.8173299205098818e-123, 32'sd1.0888019698016567e-125, 32'sd-2.1139994741860844e-127, 32'sd-3.082114677645217e-125, 32'sd0.11909334054994235, 32'sd0.041893783851153846, 32'sd0.06157967792496763, 32'sd0.08816589173202505, 32'sd0.03682818610660784, 32'sd0.06690676829760116, 32'sd-0.00717620628704431, 32'sd0.06449379621799399, 32'sd0.12578415280220437, 32'sd0.06315569500160034, 32'sd0.08372804404212089, 32'sd0.06953091166061087, 32'sd0.0010380184181025486, 32'sd0.08667171480145681, 32'sd0.08997632556986712, 32'sd-0.024847590241812618, 32'sd-0.058057187269995515, 32'sd0.029500684784079023, 32'sd-0.03314405101708578, 32'sd0.041468079836591745, 32'sd-1.0985983129458586e-114, 32'sd3.309783174816478e-119, 32'sd-1.132274086233112e-117, 32'sd-1.802845757859349e-123},
        '{32'sd-2.0524650604698404e-118, 32'sd-5.8349820875548866e-120, 32'sd1.1782695272662472e-122, 32'sd3.553490412159783e-116, 32'sd7.708741497967194e-117, 32'sd-1.3402111986372093e-127, 32'sd-4.7164507915098985e-119, 32'sd5.9209866175586025e-127, 32'sd4.628074250812244e-118, 32'sd3.092762325941508e-120, 32'sd-3.443450560799795e-114, 32'sd2.0465953890012907e-127, 32'sd-0.05874711249486108, 32'sd-0.045985881608872715, 32'sd-0.02030154488322199, 32'sd0.028493938374370434, 32'sd2.881911096695432e-122, 32'sd1.4872486936838964e-127, 32'sd-3.4577272111288314e-118, 32'sd-4.831873284956975e-118, 32'sd5.61695247252935e-124, 32'sd7.285737046898218e-125, 32'sd-1.0295140579651814e-123, 32'sd-2.600417826777905e-124, 32'sd-2.564263709633182e-126, 32'sd7.339218050260731e-121, 32'sd1.5486197645006335e-117, 32'sd-4.039309531954532e-118, 32'sd1.0530764893175685e-121, 32'sd3.2457138097212925e-121, 32'sd-2.811519858652752e-121, 32'sd2.730763855904955e-122, 32'sd0.049169814294196354, 32'sd0.10303537515343363, 32'sd-0.1035749132698456, 32'sd-0.02633322787595957, 32'sd0.015359045516865726, 32'sd-0.11433119531517172, 32'sd0.007874537119589234, 32'sd0.03761877985865268, 32'sd-0.020047306102103698, 32'sd0.06707904182487297, 32'sd0.059498092922336196, 32'sd-0.0374547590140032, 32'sd0.05157760146423232, 32'sd0.12797505243485718, 32'sd0.05456509586839255, 32'sd0.055034578071210885, 32'sd0.05065484229661779, 32'sd0.08850104327234264, 32'sd0.026025700653050165, 32'sd0.05090518675076474, 32'sd6.311891286998575e-124, 32'sd-2.8921028236153315e-115, 32'sd3.112347712812365e-114, 32'sd3.993405493911018e-124, 32'sd-2.8442313942020364e-114, 32'sd-2.427952454384627e-122, 32'sd0.04846494225497736, 32'sd0.10042646861220804, 32'sd0.024529881480037513, 32'sd0.07046510723613507, 32'sd0.04142028267621527, 32'sd0.0023652813933124155, 32'sd-0.06986144139921752, 32'sd-0.03620307748170771, 32'sd-0.026529841340547543, 32'sd-0.029311106449449616, 32'sd0.07901025160348168, 32'sd-0.02689634580546368, 32'sd0.01281677101897535, 32'sd-0.10878521050809835, 32'sd0.03219078631704646, 32'sd-0.0010361526529118906, 32'sd0.03239116934812954, 32'sd0.06628002713511302, 32'sd-0.006669016049228584, 32'sd-0.017628749645549443, 32'sd0.05964249438359792, 32'sd0.04794929990468464, 32'sd-0.017295552570348822, 32'sd0.04879104950966564, 32'sd-2.627282498685635e-117, 32'sd7.151235202540191e-115, 32'sd4.562135027636618e-123, 32'sd-1.6257673525236854e-115, 32'sd-0.025177983000295702, 32'sd0.007691757395431897, 32'sd-0.02450631485024264, 32'sd-0.008894595942337491, 32'sd0.0983491402291214, 32'sd0.09601743296818428, 32'sd0.14033103806347336, 32'sd-0.04776814656439742, 32'sd0.03947008413034343, 32'sd-0.01977054208082917, 32'sd-0.04437686693062334, 32'sd-0.05935394516069281, 32'sd0.1285448403772686, 32'sd0.02928284829553042, 32'sd-0.035355518690518825, 32'sd0.011163257145948405, 32'sd-0.07377504023134117, 32'sd-0.13753481283714972, 32'sd-0.06787376486018179, 32'sd-0.046722880332538394, 32'sd0.08535837868754548, 32'sd-0.004165455242815395, 32'sd0.07054908329717081, 32'sd0.03669549595600134, 32'sd0.09931965859924562, 32'sd8.843768724620681e-127, 32'sd-2.231830394698318e-126, 32'sd0.05236558322708531, 32'sd0.051554103888405145, 32'sd0.03612827189159458, 32'sd0.0013968931660181057, 32'sd0.04849489050743851, 32'sd0.028711240090148343, 32'sd-0.010488870008339611, 32'sd0.0028354432296487406, 32'sd-0.0029946232195463113, 32'sd-0.005206981663799705, 32'sd0.06971995365291837, 32'sd0.09865010468449442, 32'sd0.0374710001924969, 32'sd0.008154081006896923, 32'sd-0.007928679690574472, 32'sd0.0721087223026345, 32'sd-0.08661807433118175, 32'sd0.07774686560465595, 32'sd0.015474306796913116, 32'sd-0.13309989289098995, 32'sd0.01136762486705739, 32'sd-0.14383822719863545, 32'sd0.053119333346778354, 32'sd0.06140821421093544, 32'sd0.023418691264344284, 32'sd0.07116319672161762, 32'sd0.08250342585546185, 32'sd1.3502074392996326e-119, 32'sd0.04340891157117026, 32'sd-0.02387402283394307, 32'sd-0.05638217570274655, 32'sd-0.056546633575040535, 32'sd0.05380629950673428, 32'sd-0.07135922246471767, 32'sd0.04606749199253045, 32'sd-0.06297079806203883, 32'sd-0.06503144900011477, 32'sd0.08994605814663674, 32'sd-0.008869938765827689, 32'sd-0.03518490458652233, 32'sd0.012382519709783832, 32'sd0.10676302451939693, 32'sd0.09229545914221605, 32'sd-0.03154895063950735, 32'sd-0.16130073090941474, 32'sd-0.11244697633087822, 32'sd-0.020976864512797948, 32'sd-0.02781261760762945, 32'sd-0.04827080612819538, 32'sd-0.04182913490665971, 32'sd0.03146601832292977, 32'sd0.032819700286774445, 32'sd0.01435868849245195, 32'sd-0.05055686707679847, 32'sd0.013732341702392651, 32'sd1.3095069015520063e-122, 32'sd0.06002803823981637, 32'sd0.05038227395513999, 32'sd-0.023474024192463798, 32'sd-0.019473883448026027, 32'sd-0.04576066024291415, 32'sd-0.1539202744493198, 32'sd-0.1464005973903516, 32'sd-0.0853002048395739, 32'sd0.05116717506582148, 32'sd-0.05625116314004117, 32'sd-0.11019473948500556, 32'sd-0.051409249041632736, 32'sd-0.04166603525279373, 32'sd-0.021009310418555166, 32'sd0.009672454115138314, 32'sd0.014510775162951193, 32'sd-0.07216194623549797, 32'sd-0.09392033893054552, 32'sd-0.22154407716153143, 32'sd-0.04188354871631176, 32'sd-0.06046941634043615, 32'sd-0.049365823554576874, 32'sd0.0029181721149850715, 32'sd0.010722675457349713, 32'sd-0.10257841520704992, 32'sd-0.11955723450198075, 32'sd-0.04284311063955631, 32'sd0.03820882397356972, 32'sd0.018330497232984827, 32'sd0.08502046705484026, 32'sd-0.015831936360570002, 32'sd-0.008761540366336055, 32'sd0.09578551672729436, 32'sd-0.009808908755963783, 32'sd0.00011581120531055817, 32'sd0.05372385610407043, 32'sd-0.0541926365517503, 32'sd-0.03124156658821529, 32'sd-0.11295935914221927, 32'sd-0.03716211972981214, 32'sd0.0915795448902509, 32'sd0.014140425084619017, 32'sd0.06648431926445927, 32'sd0.19816582711767677, 32'sd0.032431335015256114, 32'sd-0.09221853647966584, 32'sd-0.01674494013949061, 32'sd-0.004235591546096198, 32'sd0.01377245034850178, 32'sd-0.08260241452010772, 32'sd0.023766966280668905, 32'sd0.030463891049062396, 32'sd0.023169551420755868, 32'sd0.04310734632808794, 32'sd0.019946468006177585, 32'sd0.05634304836463452, 32'sd0.046413978664122765, 32'sd-0.025535706676239948, 32'sd0.10407161793358558, 32'sd0.06295631326919854, 32'sd-0.022524084810553714, 32'sd-0.05467593723668376, 32'sd0.07958810077288357, 32'sd0.10043948700250752, 32'sd0.028717113262485376, 32'sd-0.12514115375414497, 32'sd-0.14913605133948069, 32'sd-0.12466306967925345, 32'sd-0.10264348438795375, 32'sd0.04027504152949894, 32'sd0.08877257650625213, 32'sd0.15624830366712542, 32'sd0.09386842871979445, 32'sd0.003208589645657213, 32'sd0.03156052032314793, 32'sd0.06168462152664476, 32'sd-0.03823179114559, 32'sd-0.12365470113906213, 32'sd-0.12263307182279626, 32'sd0.0004935472681210832, 32'sd0.09897695304313477, 32'sd0.07562719932382196, 32'sd0.04020159145544289, 32'sd-0.006821215753506105, 32'sd-0.01472921268672405, 32'sd0.14102344571312062, 32'sd-0.011999979286140135, 32'sd-0.03846290979040625, 32'sd0.00695611221122496, 32'sd0.00022155403592676357, 32'sd-0.021564539787813142, 32'sd0.12216790102412911, 32'sd-0.04920885781349831, 32'sd-0.04387682632836687, 32'sd-0.01182222044347607, 32'sd-0.13462829548299632, 32'sd-0.07076507262107838, 32'sd0.10584219787129141, 32'sd0.012801711965575748, 32'sd0.03260393737182837, 32'sd0.0775068275594435, 32'sd-0.048754850036090355, 32'sd0.10979416423122093, 32'sd-0.09169600158434896, 32'sd0.03449412687080186, 32'sd-0.006016307893371603, 32'sd-0.04424759386767836, 32'sd-0.021059440531886017, 32'sd-0.027151623101794798, 32'sd0.06989511223422981, 32'sd-0.008605441242557986, 32'sd-0.028033792113866203, 32'sd0.09780735905470316, 32'sd0.018793922937116663, 32'sd0.056888768101695956, 32'sd-0.05174087179123138, 32'sd0.05861841804162223, 32'sd-0.06410197113316889, 32'sd0.06214039852814822, 32'sd0.002916272893684674, 32'sd-0.09090722471780699, 32'sd-0.05034623272370074, 32'sd-0.10335192315035437, 32'sd-0.1013962707176637, 32'sd0.08299502522432216, 32'sd0.068386785352636, 32'sd-0.04331523978556215, 32'sd-0.08602867942432642, 32'sd0.05561409684796691, 32'sd-0.041463602362269016, 32'sd0.08958182114137195, 32'sd-0.02621608290525309, 32'sd-0.014375193761393163, 32'sd0.004114108751109656, 32'sd0.03462642160466407, 32'sd0.01119183692335344, 32'sd0.05155966949277589, 32'sd0.015566062910289342, 32'sd0.08190122065358518, 32'sd-0.028416793888625017, 32'sd-0.028219076268696318, 32'sd0.0547061261801557, 32'sd-0.11531919989807994, 32'sd-0.09511614826173292, 32'sd-0.02051414042894808, 32'sd-0.04376122915430653, 32'sd0.05491075884281311, 32'sd0.06667615703620153, 32'sd-0.06264904598086997, 32'sd-0.03719384289384184, 32'sd-0.10716527946814632, 32'sd0.003382712550398496, 32'sd0.11975849999910991, 32'sd0.059457949877763816, 32'sd0.0772994496025147, 32'sd-0.004706967098969045, 32'sd0.0011767607007909008, 32'sd-0.05324370555579913, 32'sd0.08120344676489169, 32'sd0.08548624388696156, 32'sd0.07571359899475956, 32'sd0.06802378497860709, 32'sd0.0914226930006909, 32'sd-0.012247476221025937, 32'sd-0.11800851253101508, 32'sd0.03967491903675878, 32'sd0.02173199711447905, 32'sd0.1021102403378904, 32'sd0.06543900190519081, 32'sd0.05190733731269308, 32'sd-0.15096406804454954, 32'sd0.0010353095938896444, 32'sd-0.07952643615546223, 32'sd0.0264209747573517, 32'sd0.09088812469062624, 32'sd0.08450790510681642, 32'sd-0.03208859031833858, 32'sd-0.006511665306651922, 32'sd-0.06378220470644348, 32'sd0.13803835442093404, 32'sd0.19915563813210524, 32'sd0.18565387031601815, 32'sd0.040990255767441156, 32'sd0.10282678980203927, 32'sd-0.00398877694337175, 32'sd0.0632481224664205, 32'sd0.00247146881332936, 32'sd0.007016481557916537, 32'sd0.008524563563291883, 32'sd0.125018237071238, 32'sd0.11090783950078963, 32'sd0.2019576665526387, 32'sd0.13926580803179042, 32'sd0.004542812399525881, 32'sd-0.06834293373326852, 32'sd0.05039660233885183, 32'sd-0.08065135747525021, 32'sd0.026055491363723683, 32'sd-0.059327805877233936, 32'sd-0.11422681010032787, 32'sd0.06430387905165337, 32'sd0.12490374983176582, 32'sd0.11662753331244384, 32'sd0.07251853890874378, 32'sd-0.056796304518359896, 32'sd-0.027725892689592208, 32'sd0.14276431352644903, 32'sd0.1767540344486664, 32'sd0.10480929715697267, 32'sd0.0991391036301391, 32'sd0.08554517924077958, 32'sd0.15273073805112894, 32'sd0.08061540696178703, 32'sd0.07843323092559348, 32'sd-0.1126063731636604, 32'sd0.014567909822636683, 32'sd-0.06874364148029902, 32'sd-0.0541816869493039, 32'sd0.096173174600714, 32'sd0.10666865131839778, 32'sd-0.08780317576144601, 32'sd0.02759640698438889, 32'sd0.007966761255264373, 32'sd0.1275241725719335, 32'sd-0.022484845654270166, 32'sd-0.02215034977079944, 32'sd-0.0691817414877323, 32'sd-0.14853813142929623, 32'sd0.05046035349257501, 32'sd-0.05040573013051246, 32'sd0.0455169489887214, 32'sd0.03828930732842927, 32'sd0.03871248221382781, 32'sd-0.007717846472930429, 32'sd0.07450852286003852, 32'sd0.19928737910993952, 32'sd0.20720388421447877, 32'sd0.1299758524219962, 32'sd-0.007782086895313886, 32'sd0.03596179544893114, 32'sd0.04824422438069201, 32'sd-0.09955674345388665, 32'sd-0.17713284388015446, 32'sd-0.04511271471100416, 32'sd-0.10334321992281419, 32'sd0.037353725448874844, 32'sd0.10287132700109097, 32'sd0.13003313763543656, 32'sd-0.06279592871772069, 32'sd0.03509347003841608, 32'sd0.05144345067596775, 32'sd0.1109534254665554, 32'sd0.07364510165312751, 32'sd0.033544076414355264, 32'sd0.012510080440683892, 32'sd-0.0476090047723513, 32'sd0.019571094535964006, 32'sd-0.023693917744363642, 32'sd-0.07298427403299584, 32'sd-0.028551604252209636, 32'sd-0.14162116248190398, 32'sd-0.05616225634205146, 32'sd0.12047194240262189, 32'sd0.1422919452827237, 32'sd-0.02133253895715878, 32'sd-0.018278376121797026, 32'sd0.0026344319528763148, 32'sd0.017900028984180905, 32'sd-0.026075540302669644, 32'sd0.06363238678710094, 32'sd-0.12121787394455137, 32'sd0.04182228805005682, 32'sd-0.03678562298632533, 32'sd-0.04671655734973578, 32'sd0.051913581370321205, 32'sd0.04075262390302914, 32'sd-0.03391311808102997, 32'sd0.10411451839761088, 32'sd0.012672259991582184, 32'sd0.04439562588161623, 32'sd0.061679144740645855, 32'sd0.08525462039750341, 32'sd-0.07150157752409966, 32'sd-0.0975418193992494, 32'sd-0.10190598477153144, 32'sd-0.21117208891685116, 32'sd-0.2356828139862029, 32'sd-0.19962593687538632, 32'sd-0.2738160744736449, 32'sd-0.05626031744904508, 32'sd0.024383639749775487, 32'sd-0.015171543188620013, 32'sd-0.05045287681321288, 32'sd-0.09489366883957544, 32'sd-0.18341309714555118, 32'sd0.005609466727088627, 32'sd0.02948021660221405, 32'sd0.09769485005725663, 32'sd-0.05235191238901677, 32'sd0.0980791438146084, 32'sd-0.0025008323399367833, 32'sd0.02853511379263492, 32'sd0.07818725093473751, 32'sd-0.015198205978723213, 32'sd-0.04486177796284506, 32'sd0.018997858157695897, 32'sd-0.022403497909713663, 32'sd-5.403801792770375e-118, 32'sd-0.016477437077422708, 32'sd-0.05012959402817485, 32'sd-0.010917448334723865, 32'sd0.05498429451463424, 32'sd0.005674735564153115, 32'sd-0.11529946193223428, 32'sd-0.18519367916492452, 32'sd-0.16730041306239524, 32'sd-0.18515426851046082, 32'sd-0.1865975474843951, 32'sd-0.07526149605600067, 32'sd-0.0801551490015558, 32'sd-0.1009300823037784, 32'sd-0.04429130771803485, 32'sd-0.06538675559316544, 32'sd-0.016400305584191643, 32'sd-0.11035521660369046, 32'sd-0.08480211291890291, 32'sd0.018239304157835545, 32'sd-0.025762645174319372, 32'sd0.05000115194330093, 32'sd0.009264516083520566, 32'sd-0.07249902620543382, 32'sd0.04755684563310755, 32'sd-0.03222871496331096, 32'sd0.030454902674390275, 32'sd0.023731321451572085, 32'sd-0.007450823616843703, 32'sd0.032400878503697335, 32'sd-0.05775422017997935, 32'sd0.09371987010859498, 32'sd-0.02765473926740168, 32'sd0.06836888194800132, 32'sd0.08393893496686734, 32'sd-0.07706867825135208, 32'sd-0.15078357165500647, 32'sd-0.05936703628126809, 32'sd-0.07082439045834467, 32'sd-0.08511216648181119, 32'sd-0.08468718687966029, 32'sd-0.04314754420273189, 32'sd-0.09931440536405861, 32'sd0.0034181628696292495, 32'sd-0.025888664905770763, 32'sd0.015281456360129774, 32'sd-0.009191642656899446, 32'sd0.06889114493627035, 32'sd-0.02987735392443078, 32'sd0.024942809238063433, 32'sd-0.08821914178769445, 32'sd-0.11841199179968315, 32'sd-0.029300222241189475, 32'sd-0.02723487234046844, 32'sd-0.045149166141537654, 32'sd0.02722125460253831, 32'sd0.035930282848677705, 32'sd0.02306479833665598, 32'sd0.04499859317206299, 32'sd0.12775645588059242, 32'sd0.06388979915896581, 32'sd0.051264465709013565, 32'sd0.08786658347445953, 32'sd0.07162976081307476, 32'sd0.043407867390096756, 32'sd0.09375395296543639, 32'sd-0.040179195676721687, 32'sd-0.08338561361662823, 32'sd-0.062381376668096296, 32'sd-0.029082225396399278, 32'sd-0.06367854393563444, 32'sd-0.10334964359415941, 32'sd-0.02426887540083552, 32'sd-0.020579054862140074, 32'sd0.11953345168855233, 32'sd0.028808190120745383, 32'sd-0.02572701043091282, 32'sd0.053251991952992996, 32'sd-0.1471657792631247, 32'sd-0.14527173438641935, 32'sd-0.09646035038889963, 32'sd-0.10132260426945806, 32'sd0.06903029880482815, 32'sd-0.008464090467596642, 32'sd1.3182768900461975e-122, 32'sd-0.06930095586969727, 32'sd0.01760346406360393, 32'sd0.01888058664068197, 32'sd0.05442557363003053, 32'sd-0.032019340028445184, 32'sd0.04565004597716374, 32'sd0.14010020000559117, 32'sd0.01338538826033417, 32'sd0.027744716495661906, 32'sd0.035393440417831115, 32'sd-0.016587468720423767, 32'sd-0.030839106599421188, 32'sd-0.10914825362961426, 32'sd0.06302399724427295, 32'sd0.05841793098093051, 32'sd0.12284915167758875, 32'sd0.09983069692621283, 32'sd0.11201781106175535, 32'sd-0.09025279198285849, 32'sd-0.00508813825195637, 32'sd-0.020438831001957775, 32'sd-0.1673852041362798, 32'sd-0.07377870472103053, 32'sd-0.12941136405848191, 32'sd-0.09808798531325745, 32'sd0.10237962760473412, 32'sd0.032436872808186995, 32'sd0.1294102744195115, 32'sd0.0339276426787877, 32'sd0.02289687344642153, 32'sd-0.0317119493515261, 32'sd0.008494328424279919, 32'sd-0.059662318183273035, 32'sd-0.03631201678653674, 32'sd0.00617646388729305, 32'sd-0.055540971598541135, 32'sd0.03610647050221891, 32'sd0.06876675689116256, 32'sd0.09691159065400795, 32'sd-0.004232119317526242, 32'sd0.008842381529434432, 32'sd0.10704803345691995, 32'sd-0.011339642605443737, 32'sd0.07473112486418576, 32'sd0.03481369721843148, 32'sd0.05546496900961279, 32'sd-0.01693708668720128, 32'sd0.08259972997240007, 32'sd-0.1499193671282167, 32'sd-0.02480279216940861, 32'sd-0.07090083781745458, 32'sd-0.10123313506248113, 32'sd-0.024804659072951384, 32'sd-0.016052133750199586, 32'sd-0.030358856702402175, 32'sd0.07969366397724845, 32'sd0.06503087217568974, 32'sd0.03711179291563931, 32'sd-0.025170677921447084, 32'sd0.08657123186473357, 32'sd-0.03148785655188331, 32'sd-0.0872294209992156, 32'sd0.01743556316841783, 32'sd0.0232481011657899, 32'sd-0.045295199496722706, 32'sd0.08790176730543864, 32'sd-0.014440175551339238, 32'sd-0.01597583642837484, 32'sd-0.014859444881817726, 32'sd0.016061562790404847, 32'sd-0.05543834233695307, 32'sd0.053776113780513064, 32'sd-0.0025098326598407754, 32'sd-0.07305513475482873, 32'sd-0.05608586341028097, 32'sd-0.11578191073039702, 32'sd-0.0935349662123766, 32'sd-0.09293416145642858, 32'sd0.03692994037774627, 32'sd-0.10059315991998694, 32'sd-0.021753330984549017, 32'sd0.10351386794848721, 32'sd0.024489184118622134, 32'sd2.3348986789779746e-119, 32'sd0.04370702586903926, 32'sd0.015155794348400827, 32'sd0.12585422466387286, 32'sd0.008830047711070642, 32'sd0.0034481730062757374, 32'sd-0.07626417990758665, 32'sd-0.03083533188987052, 32'sd0.04246169525714339, 32'sd0.0124322953500538, 32'sd0.1989741773842179, 32'sd0.18751705420036222, 32'sd-0.004220015147684186, 32'sd0.0042417424501165575, 32'sd0.023597382582014617, 32'sd-0.09390893681620772, 32'sd-0.027637057617679275, 32'sd0.06058816789337459, 32'sd-0.040435839610626925, 32'sd-0.08280818885670596, 32'sd0.05577541541311693, 32'sd-0.01835478110231073, 32'sd-0.05601846977722786, 32'sd0.002610943135695012, 32'sd0.04095677315391465, 32'sd0.011449354588831713, 32'sd0.03218953983512399, 32'sd1.4146567489672997e-118, 32'sd-1.6349421799794357e-123, 32'sd6.456549551901884e-116, 32'sd0.02533188931733582, 32'sd0.10233862515746321, 32'sd0.020071908862221353, 32'sd0.020598703482505497, 32'sd-0.016250169790594866, 32'sd0.02851470049122432, 32'sd-0.0027532696116765103, 32'sd0.20468429965264598, 32'sd0.12541721332037786, 32'sd-0.027697690636212788, 32'sd-0.07327821004932025, 32'sd0.07515077821706645, 32'sd0.11636493541788928, 32'sd-0.021652489332484735, 32'sd0.0905025792143538, 32'sd0.03684228666744032, 32'sd0.02066198982445268, 32'sd0.09669238822962332, 32'sd0.006690774259842456, 32'sd-0.07880713917759107, 32'sd-0.0019745304685801104, 32'sd-0.04604037221982053, 32'sd0.0022520745064776556, 32'sd0.06368400637414848, 32'sd0.01108633065026452, 32'sd-6.570459718871512e-115, 32'sd-1.7284317320010596e-125, 32'sd2.779755594405155e-114, 32'sd0.0745661125141198, 32'sd0.06143458786360052, 32'sd0.0286824379396701, 32'sd-0.03422055106222991, 32'sd0.037350347717193234, 32'sd-0.030850412325240634, 32'sd-0.04757395814689539, 32'sd0.12128328984122635, 32'sd0.029320972640557226, 32'sd-0.06229677526201741, 32'sd-0.02737444762340069, 32'sd-0.057906897557510564, 32'sd0.033792322610587074, 32'sd-0.06351623308579117, 32'sd-0.048987378995204674, 32'sd-0.08651624787948028, 32'sd-0.010565235424895575, 32'sd0.0072654915088456095, 32'sd0.033950600826994366, 32'sd-0.027140109411189346, 32'sd-0.03863192702708758, 32'sd0.04377743321900092, 32'sd0.04950040692538864, 32'sd-0.033577782819827325, 32'sd-0.010664378734506628, 32'sd-1.0375366076984047e-122, 32'sd9.249307907843046e-119, 32'sd2.232587270186013e-124, 32'sd-4.431643435991359e-120, 32'sd0.03355473123553707, 32'sd-0.046280405946787465, 32'sd0.011811369635203423, 32'sd-0.06209332268472281, 32'sd0.033269079004057615, 32'sd-0.0825962247910952, 32'sd0.014723576133216686, 32'sd-0.02770528172790072, 32'sd-0.0862479927676703, 32'sd-0.048730473056317634, 32'sd0.030499392695707322, 32'sd-0.0162801465960453, 32'sd-0.06645811014983469, 32'sd-0.03227977822373283, 32'sd0.04116719268576002, 32'sd-0.0027013175510767116, 32'sd-0.12867231993729353, 32'sd0.02359277218054878, 32'sd-0.09726418625527437, 32'sd-0.03122123298065607, 32'sd-0.023855025328829684, 32'sd0.04958317714558531, 32'sd-0.010586449131799756, 32'sd1.753572338482618e-122, 32'sd-6.21027764069772e-126, 32'sd1.508931409538217e-127, 32'sd-3.270060413454222e-122, 32'sd5.254253896677571e-119, 32'sd-1.2680348708918126e-120, 32'sd0.039051206595796875, 32'sd0.03839235689414469, 32'sd0.019299249445829184, 32'sd0.028680750391680988, 32'sd-0.010024915628476683, 32'sd-0.01632881275262323, 32'sd0.067758823421512, 32'sd-0.002298845345360616, 32'sd0.018887562573427236, 32'sd-0.04698882729478073, 32'sd-0.018756491749769517, 32'sd0.09562344069859785, 32'sd-0.018880077427085033, 32'sd0.04395179373014352, 32'sd-0.04435296047391477, 32'sd-0.03492701606632929, 32'sd0.007945034785166411, 32'sd-0.00280482427868056, 32'sd-0.06916784113767929, 32'sd0.03644165866088938, 32'sd4.866650824299879e-117, 32'sd6.142294370614981e-121, 32'sd-2.136607976744015e-122, 32'sd2.1846675090889244e-121},
        '{32'sd-6.260478264503677e-116, 32'sd-3.48201947028556e-115, 32'sd-4.555471851575646e-125, 32'sd-1.9190692548392325e-115, 32'sd4.4309474726682845e-122, 32'sd7.607239407970755e-121, 32'sd1.7377204274811111e-124, 32'sd7.505912088576645e-118, 32'sd2.5564452687171085e-126, 32'sd2.114965440285718e-117, 32'sd-1.1483323176477657e-118, 32'sd1.06734129306629e-115, 32'sd-0.016708955875569215, 32'sd-0.02381182294934761, 32'sd-0.008847874621968245, 32'sd-0.02386554131319704, 32'sd9.937830861499071e-126, 32'sd4.526574740689395e-123, 32'sd8.415243768919222e-126, 32'sd2.295473862691993e-119, 32'sd1.9304392436219044e-127, 32'sd-1.0520804530593604e-122, 32'sd4.6923322833256905e-123, 32'sd1.671901747935257e-122, 32'sd-1.4047700861514637e-125, 32'sd-6.292128418434152e-124, 32'sd2.5291199069838085e-123, 32'sd-2.256396571025814e-120, 32'sd3.6142728073977655e-129, 32'sd-2.8237993800668025e-124, 32'sd-1.3393082170867273e-122, 32'sd-4.269066393076538e-127, 32'sd-0.06018565174067595, 32'sd-0.09039655951943189, 32'sd-0.0786070287517709, 32'sd-0.0627573671003243, 32'sd-0.05259042048473827, 32'sd0.006115731396195432, 32'sd-0.009816801895374386, 32'sd-0.11264823194721461, 32'sd-0.034071871665729385, 32'sd-0.10572677246102065, 32'sd-0.03675115537698052, 32'sd-0.0995112095470745, 32'sd-0.015688123756503792, 32'sd-0.05779637845846863, 32'sd0.049792484436376995, 32'sd-0.03251556375815411, 32'sd-0.08780192114655742, 32'sd-0.06268558366070742, 32'sd-0.02984532199255513, 32'sd-0.053046094884966574, 32'sd4.358576221360476e-121, 32'sd-8.766140627961843e-126, 32'sd-4.326385941909544e-125, 32'sd1.0536017985540574e-122, 32'sd6.560886830276075e-127, 32'sd9.075542766138331e-119, 32'sd-0.02366194968719847, 32'sd-0.08216660101431843, 32'sd-0.0374739913731424, 32'sd-0.05038068292076244, 32'sd-0.019618046374390498, 32'sd0.049855756889531914, 32'sd0.010949149441471398, 32'sd0.023094653199510144, 32'sd0.020803729126680173, 32'sd-0.021042539620454142, 32'sd-0.081142617539335, 32'sd-0.13085220494005326, 32'sd-0.1952389420158229, 32'sd-0.024332691950868828, 32'sd-0.02958431892207645, 32'sd-0.08259360447894779, 32'sd0.046142636977136275, 32'sd0.14283138872061446, 32'sd0.009869547431116937, 32'sd-0.04935138415706799, 32'sd-0.03280497081518476, 32'sd-0.11242452274592567, 32'sd-0.06987532445992661, 32'sd0.0020574145642720315, 32'sd-2.8292671578387196e-125, 32'sd2.545594373523739e-126, 32'sd1.5564770191122312e-126, 32'sd7.87418587121111e-125, 32'sd-0.07825975835225316, 32'sd0.04347929607518509, 32'sd-0.10031198442836933, 32'sd0.05813669456377503, 32'sd0.059921143367965925, 32'sd-0.06219100240676863, 32'sd-0.08596288985177125, 32'sd0.006015687244604927, 32'sd0.022058589014406615, 32'sd-0.0738867290518971, 32'sd-0.09254554994899493, 32'sd-0.11203816998126745, 32'sd0.051654952403880385, 32'sd0.010068226892956712, 32'sd-0.019745179786159965, 32'sd0.14251318918271658, 32'sd0.06276682664209464, 32'sd0.04151668038267739, 32'sd0.11065887647818995, 32'sd-0.02530871401409068, 32'sd-0.05313369388542229, 32'sd-0.03603079637481708, 32'sd0.08023332802218848, 32'sd0.08102576277442383, 32'sd0.06209874311947834, 32'sd1.969545033104772e-117, 32'sd-4.664620991473124e-115, 32'sd-0.05248552785986366, 32'sd0.03967842788997917, 32'sd-0.0536660674623748, 32'sd-0.11955207016182841, 32'sd-0.02415811322404599, 32'sd-0.022221381844860236, 32'sd-0.13893858687475338, 32'sd-0.05486751189800841, 32'sd-0.09573306888893392, 32'sd0.028944782450734872, 32'sd-0.14236280818644043, 32'sd-0.08174270867076366, 32'sd-0.05700038076399789, 32'sd0.03474327628306729, 32'sd-0.057193513418168695, 32'sd0.04739330565446581, 32'sd-0.04897190958281819, 32'sd-0.014185929181915777, 32'sd0.034482337965888066, 32'sd-0.021343268664783425, 32'sd-0.035471195486772515, 32'sd0.06049333262743327, 32'sd0.025460575795201966, 32'sd0.07334601041583044, 32'sd-0.016655545003419942, 32'sd-0.016605526547149096, 32'sd0.047954708587136914, 32'sd-3.004006560385326e-122, 32'sd-0.0049259990918817526, 32'sd-0.0013530352159172095, 32'sd0.08056004757174416, 32'sd-0.14074591714116294, 32'sd0.007814840408993289, 32'sd-0.010668082405471301, 32'sd-0.054714667041571984, 32'sd-0.18767222759667745, 32'sd0.04081077089755008, 32'sd0.003424247300489676, 32'sd-0.055093007810174816, 32'sd0.0063592885797843805, 32'sd-0.12069039475358237, 32'sd-0.006438997326214914, 32'sd0.08258714534027507, 32'sd0.1223492106973245, 32'sd0.14386692144986804, 32'sd0.03824526850115028, 32'sd0.05386007253844483, 32'sd0.028033074546631887, 32'sd0.14182809144863498, 32'sd0.11556991077732102, 32'sd-0.003389388427137117, 32'sd0.02519401809725057, 32'sd-0.04062219836646509, 32'sd0.0003789703815562381, 32'sd0.037276082814009494, 32'sd3.550638614491288e-114, 32'sd0.04389566522790196, 32'sd0.03369538723848751, 32'sd0.07077150398546236, 32'sd-0.12328172253218397, 32'sd0.03511453979937602, 32'sd-0.07886017536191273, 32'sd-0.11811026261287538, 32'sd0.024563752063833467, 32'sd-0.03532984963659661, 32'sd-0.10866038907334614, 32'sd-0.10144577576309248, 32'sd-0.07214168896832103, 32'sd-0.05961110586368759, 32'sd-0.01414246129571756, 32'sd0.11252987982524933, 32'sd-0.01029361596919025, 32'sd0.011302883503278406, 32'sd-0.0243365081557505, 32'sd0.02511191070795119, 32'sd0.08323781122666778, 32'sd0.05005977565324068, 32'sd0.0583740324395243, 32'sd0.09251894286449547, 32'sd0.03941807096686623, 32'sd0.04500201635674624, 32'sd-0.017779291126504324, 32'sd-0.06489509509462765, 32'sd0.017285810634892932, 32'sd-0.016295051145820395, 32'sd-0.04208600421071428, 32'sd-0.02749320483319805, 32'sd-0.08962077402132834, 32'sd-0.055392698250497786, 32'sd-0.18951364063317203, 32'sd-0.01633190840206884, 32'sd-0.11916958346968157, 32'sd-0.06050132906541581, 32'sd-0.08952476091311032, 32'sd-0.010265806940900905, 32'sd-0.0499225160859855, 32'sd-0.020604969415478683, 32'sd0.07139542556315663, 32'sd0.08543695664287619, 32'sd0.061244527127636963, 32'sd0.045991841816282346, 32'sd-0.12333591756667321, 32'sd0.06030532313700261, 32'sd0.09364866338230238, 32'sd-0.06833593149669062, 32'sd-0.0727446994481704, 32'sd-0.05607438593590255, 32'sd0.00598976464473691, 32'sd-0.03464877057662013, 32'sd-0.027310053041198004, 32'sd0.05350517636913178, 32'sd-0.023013650744976227, 32'sd-0.02847063060771331, 32'sd-0.14480830661377944, 32'sd0.014123790756521287, 32'sd-0.1494574459512247, 32'sd-0.10782273517543917, 32'sd-0.16310183411349025, 32'sd-0.09100107951410578, 32'sd-0.02401913331266188, 32'sd-0.10568108433686055, 32'sd0.009342278066422861, 32'sd0.009455076972776548, 32'sd-0.030749418737426006, 32'sd0.05209681323369268, 32'sd0.009315543554106959, 32'sd-0.024563667618362223, 32'sd-0.09829835945326211, 32'sd-0.07664963180624373, 32'sd-0.06923872745987375, 32'sd-0.038414942926590555, 32'sd0.016310691024261012, 32'sd-0.015668116279220528, 32'sd-0.10315404461289306, 32'sd-0.11376455880734379, 32'sd-0.1600027204005576, 32'sd-0.10587706046957918, 32'sd-0.08437083412710078, 32'sd0.0002909056862569889, 32'sd-0.06196996886029888, 32'sd-0.12299327388181071, 32'sd0.0034532060806832165, 32'sd0.028829659737483602, 32'sd-0.09353502299934834, 32'sd-0.04048755499666088, 32'sd0.006826229831643905, 32'sd-0.0050733370571402585, 32'sd-0.1409023770915848, 32'sd-0.032231821211241574, 32'sd-0.052627561530556026, 32'sd0.12361345823450004, 32'sd-0.10106469031876851, 32'sd-0.10788988544426369, 32'sd-0.060331364006909735, 32'sd0.008727824952927, 32'sd-0.032780990401567185, 32'sd0.04118312120098245, 32'sd-0.03860376737654544, 32'sd-0.04335729918675266, 32'sd-0.16646887284298453, 32'sd0.04238839229672232, 32'sd-0.1367621743514862, 32'sd-0.05907889655484713, 32'sd-0.06994414878325726, 32'sd-0.07716699610906333, 32'sd-0.036199029647317665, 32'sd-0.054410760249811334, 32'sd-0.06843304634730923, 32'sd-0.06416795491175012, 32'sd-0.1209300262805342, 32'sd-0.02539200023018311, 32'sd0.08681911265006645, 32'sd0.042265277683889046, 32'sd-0.1670821632833856, 32'sd-0.02626137225627922, 32'sd-0.1417055421711823, 32'sd-0.10479260289242101, 32'sd-0.03866843353995294, 32'sd0.06140054790595373, 32'sd0.12763274172232486, 32'sd-0.05064424299851095, 32'sd0.1335726057738029, 32'sd0.08508568055133897, 32'sd-0.06406312157530546, 32'sd0.05593784476132015, 32'sd0.06162441219914905, 32'sd-0.0950757643842935, 32'sd-0.12826302470264356, 32'sd-0.16129098409280043, 32'sd-0.009809537047145336, 32'sd-0.15141828531578505, 32'sd-0.08868361652096622, 32'sd0.057829712783690014, 32'sd-0.036170597948840116, 32'sd-0.06206443432780026, 32'sd0.022942976420540058, 32'sd0.016509668328001707, 32'sd-0.031513483651440875, 32'sd0.03991932882914384, 32'sd0.08273978008430775, 32'sd-0.04987181343938478, 32'sd-0.028176258483417163, 32'sd-0.0800611525154015, 32'sd-0.1854021347553447, 32'sd-0.13601318304421112, 32'sd0.035161448103480555, 32'sd-0.036635775574078856, 32'sd0.0976204816173655, 32'sd0.09416697639563444, 32'sd0.2066158343821256, 32'sd0.041868680260169315, 32'sd0.08278802284731704, 32'sd0.03410084574032017, 32'sd-0.06510808853141965, 32'sd-0.07046508542984369, 32'sd-0.18131369679554735, 32'sd-0.12628936042307, 32'sd-0.17008432838905024, 32'sd-0.05299529401788398, 32'sd-0.07285501477907426, 32'sd-0.09315088063171463, 32'sd0.06349550317346764, 32'sd0.07080069091338458, 32'sd0.02716029854553213, 32'sd0.004131761992195342, 32'sd-0.16700354679545792, 32'sd-0.06612645798797216, 32'sd-0.16570266506729514, 32'sd0.027986482853822863, 32'sd0.07746508352982352, 32'sd-0.15473640211223544, 32'sd-0.12552033288822215, 32'sd-0.07212497280087064, 32'sd0.08584135470117858, 32'sd0.07448443480004288, 32'sd0.1268534222108652, 32'sd0.15903088306748644, 32'sd0.1431012393420052, 32'sd0.05698423717145789, 32'sd0.14243317324241714, 32'sd0.03180879687537042, 32'sd-0.03349628253795217, 32'sd-0.026434977489523084, 32'sd0.06604504604744134, 32'sd-0.1752113779070383, 32'sd-0.057358776334797947, 32'sd0.052037191792095906, 32'sd0.019764784807416124, 32'sd0.04186135846852365, 32'sd-0.0014671333627133767, 32'sd-0.036490080370267707, 32'sd-0.027134887082186306, 32'sd-0.0323172386732377, 32'sd-0.12062635882301206, 32'sd-0.02147883791831349, 32'sd-0.19943760366423055, 32'sd-0.044926756863814844, 32'sd0.03921374399589545, 32'sd0.02870986405191825, 32'sd-0.16069453487130841, 32'sd0.0922974884858116, 32'sd-0.0015254343637076723, 32'sd-0.0012826848556510976, 32'sd0.1521088526592785, 32'sd0.12455346855622239, 32'sd0.13563384251940477, 32'sd0.08521893676347889, 32'sd0.12744828485420906, 32'sd0.13055771574469227, 32'sd-0.008032703660577595, 32'sd-0.0012378469956892532, 32'sd-0.017506278788847484, 32'sd-0.13685531258142355, 32'sd-0.14490241820487657, 32'sd-0.10415930771098031, 32'sd-0.047152599654323016, 32'sd-0.02718566374061871, 32'sd0.003730341769220027, 32'sd-0.0611977361000751, 32'sd-0.06730708689500649, 32'sd-0.08849043471136148, 32'sd-0.016002090837488648, 32'sd-0.08759989962200848, 32'sd-0.15130252386366647, 32'sd-0.13166402917438783, 32'sd-0.05020636969536793, 32'sd-0.10497975438641453, 32'sd0.06442981690312287, 32'sd0.11557273162654454, 32'sd0.01047017505555225, 32'sd0.020522719320736776, 32'sd0.09743406311355428, 32'sd0.12808758579377663, 32'sd0.10450443866458922, 32'sd-0.03096193812646822, 32'sd0.09649973549532857, 32'sd0.1355548679532941, 32'sd-0.07588431141761774, 32'sd-0.03609926883438515, 32'sd-0.02644730713624219, 32'sd-0.04581207815045997, 32'sd-0.01774952104136048, 32'sd-0.16500630840412045, 32'sd-0.10769076576141662, 32'sd-0.019566790357648488, 32'sd-0.017471631202923048, 32'sd0.010468891853459554, 32'sd-0.05138253854134369, 32'sd-0.06272322994644852, 32'sd-0.02324505481831371, 32'sd-0.03711059176491723, 32'sd-0.05247766564952579, 32'sd-0.005999846100112434, 32'sd-0.06481668018589341, 32'sd0.005722281640892036, 32'sd0.006523517896484175, 32'sd-0.04630697766458511, 32'sd-0.1782921307442499, 32'sd-0.1493267982869957, 32'sd0.0576023192529311, 32'sd0.008571846161191643, 32'sd0.03807341017651379, 32'sd1.0809111903254542e-05, 32'sd0.07445137746581372, 32'sd0.09960099186774661, 32'sd-0.018903751277142684, 32'sd0.09313770462789038, 32'sd0.0896816259751308, 32'sd0.07828881528669125, 32'sd0.025995709564889627, 32'sd-0.07593881565056532, 32'sd-0.07225042693519823, 32'sd-0.09599741191131313, 32'sd-0.0963520215201522, 32'sd-0.049149983022757825, 32'sd0.011585667144116438, 32'sd-0.08117733974457325, 32'sd-0.04364024750509583, 32'sd0.08256871218770294, 32'sd-0.024506901656191668, 32'sd0.05196464993305711, 32'sd-0.13317481004217463, 32'sd-0.11617735711843548, 32'sd0.01617148346413763, 32'sd-0.05922882776848092, 32'sd-0.0180971528910267, 32'sd-0.04909835119668016, 32'sd0.008696508325025545, 32'sd0.0011713094098146878, 32'sd0.06010026356216752, 32'sd0.1801573485028927, 32'sd0.09777549533264154, 32'sd-0.04795494092820908, 32'sd0.002701409860378749, 32'sd0.11065518318081219, 32'sd0.02233531013063329, 32'sd-0.04896608166476388, 32'sd-0.010583988426832015, 32'sd0.06984572822161274, 32'sd-0.044792430114264405, 32'sd-0.09798300000937799, 32'sd-0.010248746553392796, 32'sd-0.0888311632622383, 32'sd3.344913293769098e-126, 32'sd-0.02694786973004859, 32'sd-0.05589482811886265, 32'sd-0.0067425684356792965, 32'sd0.054808167901512654, 32'sd0.009133294965325604, 32'sd-0.03394322469243494, 32'sd0.05740501335394652, 32'sd-0.04757673005891822, 32'sd-0.045091827175015496, 32'sd-0.06093475112554658, 32'sd-0.03429392934759526, 32'sd-0.023398921820792007, 32'sd-0.04759110608122136, 32'sd-0.007032061186592142, 32'sd0.08348515589348028, 32'sd6.835056127573063e-05, 32'sd0.16741287126948395, 32'sd0.09218326172540116, 32'sd-0.02132531121778052, 32'sd0.04225410637520663, 32'sd0.018140382898255435, 32'sd0.02113371693331654, 32'sd0.013955559220618656, 32'sd0.011996383625893893, 32'sd-0.07351181037149333, 32'sd0.06199911127677229, 32'sd0.01732449431457446, 32'sd-0.02774197937376189, 32'sd-0.07076683643138504, 32'sd0.0668592257083104, 32'sd0.02381375166019243, 32'sd-0.05951920931565367, 32'sd0.019108711780957122, 32'sd-0.06518956142712316, 32'sd0.007756198497657646, 32'sd0.0979573102679684, 32'sd-0.027703729459212307, 32'sd-0.04940994074282296, 32'sd0.03755380605688513, 32'sd-0.05107460619365622, 32'sd-0.03952686905134078, 32'sd-0.06606758337589656, 32'sd0.011053054408324676, 32'sd0.03754544855210715, 32'sd0.14253663645325748, 32'sd0.10407129597426296, 32'sd0.11286825939943361, 32'sd-0.045533166857378585, 32'sd-0.08586026746665992, 32'sd-0.11410945758745275, 32'sd-0.06901455350186521, 32'sd-0.057357976568144925, 32'sd-0.1304377466819682, 32'sd0.00538410807083923, 32'sd0.05251033473789326, 32'sd-0.03985466869537257, 32'sd-0.0701918348601334, 32'sd0.021678185671480072, 32'sd-0.022657923400472194, 32'sd0.02416101826700156, 32'sd-0.002924166140013625, 32'sd-0.06183953362438728, 32'sd0.11425519079579623, 32'sd0.053953587323022904, 32'sd-0.016628405972216723, 32'sd0.008891043224149929, 32'sd0.041061151718531363, 32'sd-0.04985119815958549, 32'sd-0.04962671023601153, 32'sd-0.08520802617631888, 32'sd-0.12074717987535645, 32'sd0.13745104469316263, 32'sd0.036380621716041804, 32'sd0.02968416551736537, 32'sd0.11110196890536489, 32'sd-0.07795693741135959, 32'sd-0.08171712503157942, 32'sd-0.04515135199902925, 32'sd-0.050148359558498536, 32'sd-0.07399697697121314, 32'sd-0.12689512434554823, 32'sd0.0716164712975613, 32'sd-0.04174724639123974, 32'sd-6.678747849800693e-126, 32'sd-0.021481070412687885, 32'sd-0.028450757491783007, 32'sd0.06367552460165009, 32'sd-0.06297084581671125, 32'sd-0.0528198127216323, 32'sd0.11637176069578344, 32'sd0.041973224772787, 32'sd-0.07796273275052032, 32'sd0.005743812105149694, 32'sd-0.04962891236023803, 32'sd-0.012785890159505833, 32'sd-0.06830795810205977, 32'sd0.018074289299744885, 32'sd-0.09265685517174904, 32'sd0.10457168179129461, 32'sd0.11682810656456269, 32'sd0.03748370902881762, 32'sd0.12201977757952875, 32'sd0.09742140763394108, 32'sd-0.0385737137379308, 32'sd-0.03430897775847611, 32'sd-0.025208201964261327, 32'sd-0.08585917747162292, 32'sd0.025553928387943594, 32'sd-0.024181041876696754, 32'sd0.0378442640918777, 32'sd-0.04191975855679901, 32'sd-0.04194223110665529, 32'sd-0.06579414495291491, 32'sd0.012726110032983875, 32'sd0.04847389933691667, 32'sd0.030211481576242705, 32'sd0.0918230280855021, 32'sd0.11654042475991183, 32'sd0.03447996249431408, 32'sd-0.10149725218651183, 32'sd0.07182966624402047, 32'sd-0.05594635825239592, 32'sd-0.06198219539656666, 32'sd-0.011518643907180345, 32'sd-0.06662240177955911, 32'sd0.026535541529492186, 32'sd-0.014535628645260801, 32'sd0.10354949773879836, 32'sd0.012026689371755585, 32'sd-0.055235367193921796, 32'sd-0.07207254261896338, 32'sd-0.09021326656949269, 32'sd-0.20724003810659028, 32'sd-0.15863136239121406, 32'sd0.02878706633481617, 32'sd-0.0671426067812076, 32'sd-0.050953295095092783, 32'sd0.03098501045002095, 32'sd0.0010789639682591775, 32'sd-0.056716405733735695, 32'sd-0.0906187430842708, 32'sd0.049805814817315754, 32'sd-0.0795192088282253, 32'sd-0.05228465036759376, 32'sd-0.059688652366363025, 32'sd-0.06163252106961405, 32'sd0.059519156149511115, 32'sd0.026248180161129352, 32'sd-0.05582277403530889, 32'sd-0.014383925305949813, 32'sd-0.004368802638783872, 32'sd0.04608911621982698, 32'sd0.08390693098907584, 32'sd0.10915887553794497, 32'sd0.10470327046109076, 32'sd0.08080245189094673, 32'sd-0.15382137623649528, 32'sd-0.01242375127781803, 32'sd-0.0880677311728305, 32'sd-0.16595530041902737, 32'sd-0.19471333200944999, 32'sd-0.0852487898074559, 32'sd0.0421490767214421, 32'sd0.009802246770746167, 32'sd-0.026157478536377374, 32'sd-0.0029547422424119315, 32'sd-0.07483998687211406, 32'sd-2.355826656237882e-120, 32'sd0.0036833460164797057, 32'sd-0.04117603614001085, 32'sd-0.03355732609544103, 32'sd-0.028219269529457598, 32'sd0.0007959715760415098, 32'sd-0.00291573964993868, 32'sd0.01569508028469286, 32'sd-0.007459842248866027, 32'sd-0.05710521889196314, 32'sd0.030924239053748907, 32'sd-0.011943384288419685, 32'sd0.0047104611042333095, 32'sd0.08407972514983404, 32'sd0.09254078329565424, 32'sd0.14837117826652707, 32'sd0.006719233815525141, 32'sd-0.12385997480190658, 32'sd0.08298389365652693, 32'sd-0.007772610894763139, 32'sd-0.1802770336213995, 32'sd-0.12769825051285932, 32'sd-0.06482953589667971, 32'sd-0.006131599688245362, 32'sd-0.054758716411489376, 32'sd-0.01855891116294266, 32'sd0.013698378097421676, 32'sd-5.88890043726825e-115, 32'sd2.2578184409265507e-117, 32'sd-1.090419577320322e-121, 32'sd0.003116674439303783, 32'sd-0.0590677168040843, 32'sd-0.0909218964363359, 32'sd0.13521124165838505, 32'sd0.07150211362118261, 32'sd-0.023227763251526454, 32'sd-0.054739883064375654, 32'sd0.04713903723369894, 32'sd0.014498150958334597, 32'sd0.031270303185939353, 32'sd0.033291101059308624, 32'sd-0.005202534613305296, 32'sd0.0022379114671422376, 32'sd0.028355226182710684, 32'sd0.13989871040657867, 32'sd-0.03541280123280736, 32'sd-0.03223745479635303, 32'sd-0.24391269538147928, 32'sd-0.06964074724448706, 32'sd0.01544991687295015, 32'sd0.12655645081960393, 32'sd0.11124970973953048, 32'sd0.0708204192289456, 32'sd-0.16214983029096605, 32'sd-0.05654654013833941, 32'sd-1.067709298228079e-115, 32'sd2.974643101164793e-121, 32'sd-1.7851145434967612e-119, 32'sd0.0400618111178891, 32'sd-0.06199810385185942, 32'sd-0.05625759078024505, 32'sd-0.031549549461815596, 32'sd-0.009362613211301645, 32'sd0.002921062000552748, 32'sd0.004254005849326429, 32'sd-0.011298492256462848, 32'sd-0.06367024469628331, 32'sd-0.006074934485048708, 32'sd-0.09213413539057574, 32'sd-0.18295920448773956, 32'sd-0.0714397457533774, 32'sd-0.034465138996192336, 32'sd-0.06577792296377266, 32'sd-0.17246673407021373, 32'sd-0.11717456450589891, 32'sd-0.16729115802056507, 32'sd-0.07119091299245248, 32'sd0.03912299735105886, 32'sd0.0659951968230302, 32'sd0.007825373444450116, 32'sd0.048968142749252645, 32'sd0.014417794404545386, 32'sd-0.0769957736079594, 32'sd-2.337460967825533e-124, 32'sd2.1329807058319313e-127, 32'sd9.483431591048235e-119, 32'sd-3.339652816837268e-120, 32'sd-0.004812867989724892, 32'sd-0.10513071281309877, 32'sd-0.07294064147894692, 32'sd0.03916272571066304, 32'sd0.08977512691217354, 32'sd0.053485337946172114, 32'sd-0.10434307928785319, 32'sd-0.015650217237116463, 32'sd0.0575770879860627, 32'sd-0.12598993860233995, 32'sd-0.11460858082458716, 32'sd-0.11756186144849737, 32'sd-0.03685097561660723, 32'sd0.10119465894982559, 32'sd0.012455605502583901, 32'sd-0.10452995832749186, 32'sd-0.09147545191714869, 32'sd-0.08448961093241093, 32'sd0.040557502481807464, 32'sd-0.09085904044479602, 32'sd-0.02677717063721739, 32'sd-0.029828528544593523, 32'sd-0.06944500758988909, 32'sd-3.3025862579539123e-121, 32'sd-7.772710339484377e-119, 32'sd3.5369781799855324e-115, 32'sd1.3376743564767698e-122, 32'sd-1.1335425812862193e-115, 32'sd3.583632231961789e-121, 32'sd-0.027750949638810286, 32'sd-0.026379762956805927, 32'sd-0.10864878396061692, 32'sd-0.007639254402056827, 32'sd0.057696725908058764, 32'sd-0.013416365993028556, 32'sd-0.07536763557440912, 32'sd-0.1261858961225178, 32'sd0.05891251870958356, 32'sd-0.09476831760395883, 32'sd0.017606574017182974, 32'sd0.07343022983814085, 32'sd0.07909609109439392, 32'sd0.019785448754312575, 32'sd-0.07371207375835036, 32'sd-0.09827671914816363, 32'sd-0.09223560521404191, 32'sd-0.03954263700280939, 32'sd0.006114023930720085, 32'sd-0.05863851801597061, 32'sd-2.456287222467194e-115, 32'sd6.890398507555217e-121, 32'sd3.250311229941848e-127, 32'sd-1.1435186186745982e-115},
        '{32'sd2.291319465277559e-126, 32'sd-4.7244629250748894e-120, 32'sd-3.380981608044037e-120, 32'sd-1.36043455259599e-122, 32'sd1.7334454970577556e-120, 32'sd4.2153343608155937e-119, 32'sd6.800857350598269e-126, 32'sd-4.951625827672881e-118, 32'sd7.127172132008672e-116, 32'sd-4.556596605939482e-118, 32'sd-1.647642959618235e-116, 32'sd-1.436062814600989e-118, 32'sd0.09744429255230357, 32'sd0.05935933302398422, 32'sd0.11999865243264253, 32'sd0.09883667110132993, 32'sd-3.178400791238163e-129, 32'sd1.1009820114158675e-123, 32'sd-5.36635077019181e-115, 32'sd1.1814857413755002e-122, 32'sd6.098160000481667e-121, 32'sd-1.0653236793545812e-123, 32'sd1.202244105025818e-115, 32'sd-1.8969328097943708e-114, 32'sd-3.2236448834757865e-120, 32'sd6.280193898371709e-126, 32'sd1.0238876568929482e-124, 32'sd1.3293538794386817e-115, 32'sd1.0391369671351225e-122, 32'sd1.7650895742334514e-117, 32'sd-5.744016406015823e-125, 32'sd-1.5852004130109974e-117, 32'sd0.1313378348053484, 32'sd0.12076293966849862, 32'sd-0.002949473468734782, 32'sd0.09374652500281007, 32'sd0.1025167086188785, 32'sd0.0633082931688171, 32'sd0.10828201953453233, 32'sd0.028007588845596423, 32'sd0.11977913974556496, 32'sd0.08434292768127287, 32'sd0.035591405634778146, 32'sd0.01938349614386038, 32'sd0.03459792824415345, 32'sd0.05321116990003816, 32'sd0.11650696901797748, 32'sd-0.0350958661616979, 32'sd0.07840083690427235, 32'sd0.03282369411918358, 32'sd0.16085011585047884, 32'sd0.11961820070160074, 32'sd-9.510574876196514e-120, 32'sd1.7483163473231172e-116, 32'sd1.8125645757700445e-117, 32'sd9.26592918433195e-116, 32'sd1.0264187617644661e-120, 32'sd1.0887200849125524e-121, 32'sd0.146070645842927, 32'sd-0.009700716373311793, 32'sd0.023901564388169316, 32'sd-0.01733038767485777, 32'sd-0.10676959521258816, 32'sd-0.047744786117210634, 32'sd0.008169451088889413, 32'sd-0.1278030914241963, 32'sd0.010021434244957134, 32'sd0.009913572016564186, 32'sd-0.0022451777536741627, 32'sd-0.056182146468319975, 32'sd-0.0007025588295081625, 32'sd0.07532089798173072, 32'sd-0.016761631424227826, 32'sd0.05388956692501737, 32'sd-0.03333786723362111, 32'sd0.02142204219165123, 32'sd-0.0036101229027521607, 32'sd-0.051171140367997844, 32'sd-0.003449311446424673, 32'sd0.052444611304228186, 32'sd-0.04378089257939378, 32'sd0.1570803784629342, 32'sd-3.175073197806326e-120, 32'sd-1.016114484584797e-122, 32'sd-8.689563172507701e-115, 32'sd4.130591646458485e-128, 32'sd0.08907436500365452, 32'sd0.02578966165135986, 32'sd-0.06546067026634851, 32'sd0.06074723135433033, 32'sd-0.005882868423973835, 32'sd-0.06648181531466528, 32'sd0.08475766608815827, 32'sd-0.09345303355431894, 32'sd0.026636514401233293, 32'sd0.026662038942476096, 32'sd0.04500151900115604, 32'sd0.04605247472367369, 32'sd0.05578162400517851, 32'sd0.12296572526606882, 32'sd0.02843052657219291, 32'sd-0.0027006705353308774, 32'sd0.05443389394218702, 32'sd0.03250922774195626, 32'sd0.09768588269361302, 32'sd-0.013227463355462918, 32'sd0.045526680290285594, 32'sd-0.07003701465408024, 32'sd0.023591242040901517, 32'sd0.09687493606565915, 32'sd-0.009593763725512239, 32'sd-1.5777745138523595e-123, 32'sd-3.907146077108114e-125, 32'sd0.12418323209473676, 32'sd-0.0549861238265622, 32'sd0.015256835705645629, 32'sd0.03976672810852996, 32'sd0.0434397485261327, 32'sd-0.028196458997281192, 32'sd-0.04330428147682436, 32'sd0.09740271965414571, 32'sd0.01877799144004002, 32'sd0.07259945425197217, 32'sd0.05330526290638094, 32'sd0.00460445510934688, 32'sd0.04125052684014918, 32'sd0.05593024039243289, 32'sd0.06377117812663524, 32'sd0.021414071847634254, 32'sd0.0075866027597722725, 32'sd0.0619595011256659, 32'sd0.010928560706675104, 32'sd0.08913901013719759, 32'sd0.021814239642757787, 32'sd0.05848761988206823, 32'sd0.06733523850529292, 32'sd0.07392106332653897, 32'sd-0.0633916719070141, 32'sd-0.06413118340818998, 32'sd0.06353146712565462, 32'sd-2.600439224690908e-124, 32'sd0.10355137942141904, 32'sd0.0645117411021084, 32'sd-0.011371429413465165, 32'sd-0.07012987728890013, 32'sd-0.004501649760607028, 32'sd0.013499392990953504, 32'sd-0.02717046449332271, 32'sd0.09484353067986533, 32'sd0.0876349768601306, 32'sd-0.08232277735421853, 32'sd-0.10127280413976349, 32'sd-0.016721887969236408, 32'sd-0.0570258431207952, 32'sd-0.008020090612052128, 32'sd-0.08376165188542696, 32'sd-0.03171509320694642, 32'sd0.04521364441360683, 32'sd-0.07693747336649161, 32'sd-0.01744098525158181, 32'sd-0.027025368804775136, 32'sd0.006312409788995373, 32'sd-0.04996269102057793, 32'sd-0.07832177988779374, 32'sd-0.031875736656436775, 32'sd0.013672448762560562, 32'sd-0.09121612244771522, 32'sd0.03784518222399004, 32'sd-1.8725625386656086e-116, 32'sd-0.016048033511206823, 32'sd0.00897671412257751, 32'sd-0.06515320885734259, 32'sd-0.0874677995160716, 32'sd0.050361264013593435, 32'sd-0.0019635694876558893, 32'sd-0.11218216672192101, 32'sd-0.13068166186119493, 32'sd-0.05509275320965246, 32'sd-0.09233909795155087, 32'sd-0.012702667339622376, 32'sd-0.09631826984816046, 32'sd-0.09293758846069512, 32'sd-0.06454761334655955, 32'sd-0.1614139955931928, 32'sd-0.12006944691760899, 32'sd-0.14540265678329267, 32'sd-0.033695231656403736, 32'sd-0.05919028822097695, 32'sd0.025459518667958526, 32'sd0.0757108152626163, 32'sd0.06350225780507787, 32'sd-0.019982913105350712, 32'sd-0.053602044586033, 32'sd0.007966011595800859, 32'sd-0.01892188121777004, 32'sd-0.012206575279328825, 32'sd0.13614081814112877, 32'sd0.08097094124009148, 32'sd-0.12161045053280566, 32'sd0.04001610255284694, 32'sd-0.09343869794095062, 32'sd-0.04149718325569324, 32'sd0.01087292792571607, 32'sd0.05825659180043593, 32'sd-0.022846109881197712, 32'sd-0.06887398993742715, 32'sd0.0033554170976261982, 32'sd-0.1411062190755519, 32'sd-0.02529142192663177, 32'sd-0.09576498283739554, 32'sd-0.1707952260944302, 32'sd-0.21060248837296922, 32'sd-0.10952314410758203, 32'sd-0.14055457072538163, 32'sd-0.13498585564165533, 32'sd-0.029381938595783415, 32'sd-0.1691617368285551, 32'sd-0.08035108032596103, 32'sd-0.011485665701530229, 32'sd0.00460908298443669, 32'sd-0.05114737516889069, 32'sd0.014815440432995328, 32'sd-0.09443163697113333, 32'sd0.020291588468682474, 32'sd-0.017187911005555646, 32'sd0.021152893211320824, 32'sd-0.10196239170747014, 32'sd0.002363719081222371, 32'sd-0.011002679397500324, 32'sd0.03403385642608537, 32'sd0.03679221207265443, 32'sd-0.01569151127457429, 32'sd0.03345473449741402, 32'sd0.030096064828138782, 32'sd0.09441499214927279, 32'sd-0.06908390488978215, 32'sd0.0651088596136246, 32'sd0.04613648295099243, 32'sd-0.11152026355410247, 32'sd0.048046814356517226, 32'sd0.0040758504708591, 32'sd-0.019506060856763756, 32'sd-0.06124022515570977, 32'sd-0.023353869806670733, 32'sd0.048102867391833955, 32'sd0.0298030610679789, 32'sd0.03185628389887181, 32'sd0.004157967900748342, 32'sd0.06048204465322142, 32'sd0.059369147856470905, 32'sd0.043526458050236916, 32'sd0.056481543993658595, 32'sd0.09109286660070451, 32'sd0.004186815701687048, 32'sd0.01484052932213176, 32'sd0.050358225158251696, 32'sd0.10728079615110622, 32'sd0.11856880045573803, 32'sd0.06648569850065282, 32'sd0.06680694792508983, 32'sd0.13177358738935677, 32'sd0.016978997517355005, 32'sd0.10250881655941443, 32'sd0.08105576038770775, 32'sd0.18688733046609982, 32'sd0.11311636093876201, 32'sd0.15023742495597853, 32'sd0.160487475137974, 32'sd0.19683005553632657, 32'sd0.16172580587575125, 32'sd0.040940077246069656, 32'sd0.0034957839364084435, 32'sd0.13244168711942045, 32'sd0.17580938359753928, 32'sd0.12962715407774128, 32'sd-0.001448947156747497, 32'sd0.07123786744585656, 32'sd0.004847064257002167, 32'sd0.002914640345813483, 32'sd-0.1282379999566303, 32'sd0.08809065168299811, 32'sd0.0922258435827807, 32'sd0.14073065266383705, 32'sd-0.07368109928198546, 32'sd0.05863365153788069, 32'sd0.012266436756062826, 32'sd0.005560271011938944, 32'sd-0.02475671808005025, 32'sd-0.09245891427544548, 32'sd0.08275938116697014, 32'sd0.11034910118896106, 32'sd0.27835888813580584, 32'sd0.14079204071260623, 32'sd0.2554777145321302, 32'sd0.17207394971967369, 32'sd0.1603954294160504, 32'sd0.15609775884025798, 32'sd0.026750777015444264, 32'sd0.17260926924695177, 32'sd0.1652236558699397, 32'sd0.17723718843665126, 32'sd0.24730019562132666, 32'sd0.11131997180510014, 32'sd0.08297744083403759, 32'sd0.15631439975358274, 32'sd0.01973229409248515, 32'sd0.006919328894444118, 32'sd0.06097182304246117, 32'sd0.04170480317475808, 32'sd0.0501926551369537, 32'sd0.01631734510079653, 32'sd0.15388779798653213, 32'sd0.04580488754166129, 32'sd-0.07134904517166991, 32'sd-0.03759590564922788, 32'sd0.008056337087325054, 32'sd0.019503496319104748, 32'sd0.02625847646172543, 32'sd0.08159148639270923, 32'sd0.20645868724779184, 32'sd0.16628334894348448, 32'sd0.08266785680714141, 32'sd0.17733724666143402, 32'sd0.16475259769986417, 32'sd-0.015584598242111539, 32'sd0.08782773336640433, 32'sd0.1672106461604365, 32'sd0.16391912498282693, 32'sd0.10346210522359196, 32'sd-0.025360939669666238, 32'sd0.08193561495870581, 32'sd0.08777335221164005, 32'sd0.13066993141117655, 32'sd0.0875106927618785, 32'sd-0.006157204860700987, 32'sd-0.09228661211676913, 32'sd0.13349691866891922, 32'sd-0.06007730651567841, 32'sd0.060156598503887854, 32'sd-0.07696540709420029, 32'sd-0.10619922585447089, 32'sd-0.1263124261246915, 32'sd-0.08729864453867421, 32'sd-0.02536299373258003, 32'sd0.06656994422293823, 32'sd0.039790951453424, 32'sd0.11282968046602858, 32'sd0.016607030882834106, 32'sd-0.04027108783494739, 32'sd-0.059251581025607965, 32'sd-0.05426900684268255, 32'sd-0.059057633940438364, 32'sd0.054111446408392175, 32'sd-0.053458283284698364, 32'sd-0.05138612667577368, 32'sd0.06600522816300552, 32'sd0.011019368575517524, 32'sd-0.05386581001894159, 32'sd-0.008214662694919557, 32'sd-0.10294033947703941, 32'sd-0.10934855928758831, 32'sd0.01656922399627065, 32'sd0.08670701866386851, 32'sd0.05577571652556842, 32'sd0.11157723050134856, 32'sd-0.0012176102617188018, 32'sd-0.026840490553549055, 32'sd-0.06312134672607189, 32'sd-0.16748336538502884, 32'sd0.01549070078592813, 32'sd-0.058988146851425415, 32'sd-0.007356185399123339, 32'sd-0.03900489513237268, 32'sd-0.05800276480104184, 32'sd0.011442864410131792, 32'sd0.025182241244637325, 32'sd-0.08842302973863955, 32'sd-0.2467097488638228, 32'sd-0.0990366450563361, 32'sd-0.2117353900887193, 32'sd0.03143067567101659, 32'sd-0.015224475953625492, 32'sd-0.12545425966736573, 32'sd-0.13859395968770763, 32'sd-0.12056421825247766, 32'sd-0.11293642508611991, 32'sd-0.20662361946806013, 32'sd-0.1308208434733432, 32'sd-0.15610958812538517, 32'sd-0.20761944706018115, 32'sd-0.09900133456545256, 32'sd0.10324546942859876, 32'sd0.12945567647758258, 32'sd0.009643616048737933, 32'sd0.05291371568132149, 32'sd-0.0929414648747363, 32'sd0.0075858970148855575, 32'sd-0.06017531862931651, 32'sd-0.017306805074439126, 32'sd-0.11110081113223555, 32'sd-0.0605137348250018, 32'sd-0.08753942589490465, 32'sd-0.03699609827001376, 32'sd-0.06142630667534301, 32'sd-0.06287540477335025, 32'sd-0.1999580818776232, 32'sd-0.2268102412005685, 32'sd-0.052003391985833924, 32'sd-0.04051341461824659, 32'sd-0.14280960197131437, 32'sd-0.06036521851881162, 32'sd0.021515665340781875, 32'sd-0.024255946263315547, 32'sd-0.08125476825400872, 32'sd-0.14932776207004048, 32'sd-0.12172880674783461, 32'sd-0.070339780875843, 32'sd0.12976194222857784, 32'sd-0.16230440492908696, 32'sd0.07988622531619581, 32'sd0.017711990488168003, 32'sd-0.037937914676485905, 32'sd-0.03671820804263026, 32'sd-0.06712633979580952, 32'sd0.053097816041924116, 32'sd0.06434651039698569, 32'sd0.013631513574913368, 32'sd-0.023499019237889537, 32'sd-0.09044357925471164, 32'sd-0.1102060870607913, 32'sd0.013345282431360248, 32'sd-0.1529982628508808, 32'sd-0.09604853382443206, 32'sd-0.1318406387012823, 32'sd-0.07656816911637737, 32'sd-0.048642082547482514, 32'sd-0.09580520759629785, 32'sd-0.10792800343662001, 32'sd-0.14623293931847076, 32'sd-0.019064879548636626, 32'sd0.02490893869915475, 32'sd0.05951533488802637, 32'sd0.07607438433074439, 32'sd0.06076508023871324, 32'sd0.06419387072538751, 32'sd0.011919181472926895, 32'sd0.07597595783079471, 32'sd0.017091862529495818, 32'sd0.086695950923021, 32'sd-0.06454112505560708, 32'sd-0.027165594957909642, 32'sd0.11872300884667945, 32'sd0.08365747897151563, 32'sd0.07983058121679266, 32'sd0.0804728341286977, 32'sd-0.007347386245530104, 32'sd-0.10619991211564589, 32'sd-0.0727507689574382, 32'sd-0.14782236296231654, 32'sd-0.1824568931466385, 32'sd-0.08954754411942979, 32'sd-0.07463312182176167, 32'sd-0.16053557534782653, 32'sd-0.011998708779955425, 32'sd-0.1002986857594643, 32'sd-0.046993935768039265, 32'sd0.03035915759245361, 32'sd-0.004084369256209403, 32'sd0.15168408261065758, 32'sd0.11909024382459119, 32'sd-0.08602602344494012, 32'sd-0.038322998646806716, 32'sd0.0677583520511308, 32'sd-0.05032895192343329, 32'sd0.03372581926078262, 32'sd0.02197347428787224, 32'sd6.753230697717071e-117, 32'sd0.027700160988443207, 32'sd-0.09537186725778059, 32'sd0.005591928853438809, 32'sd0.11591295267565054, 32'sd0.1136260707521711, 32'sd0.09507897622342282, 32'sd-0.0670194174224558, 32'sd-0.06277519139241201, 32'sd0.017760176213409924, 32'sd-0.016211070170776738, 32'sd0.025756416603176506, 32'sd-0.01816610307351238, 32'sd-0.1111315989584832, 32'sd0.0063906395692520926, 32'sd0.008195527633300774, 32'sd-0.010632328086319595, 32'sd-0.04281482306138087, 32'sd-0.007363845851626658, 32'sd-0.13332602603693508, 32'sd0.0917365944423625, 32'sd0.10355377068411556, 32'sd-0.1741805851378618, 32'sd-0.06341344248564929, 32'sd0.06105322346953769, 32'sd-0.01366564864040822, 32'sd0.0398770647029499, 32'sd-0.0021699902620410006, 32'sd0.021499933162144394, 32'sd0.04031157783536385, 32'sd-0.02080574960535237, 32'sd0.010330102921433472, 32'sd0.057787007308150985, 32'sd0.12393428193049807, 32'sd0.0030737341042108538, 32'sd-0.0044944062658666285, 32'sd0.06483345075201175, 32'sd0.004552461306049438, 32'sd0.11573947317713, 32'sd0.058706934827164235, 32'sd0.10209331756070188, 32'sd0.06494170736487126, 32'sd-0.05070030506232719, 32'sd-0.04737424304956596, 32'sd0.013223233273380916, 32'sd0.072025697950057, 32'sd0.03790921076001122, 32'sd-0.06319802783353612, 32'sd0.019708407524814214, 32'sd0.025242277035223987, 32'sd-0.09873207760158265, 32'sd-0.06343374229130712, 32'sd0.03084410669290226, 32'sd-0.04530019420239555, 32'sd0.04794290859819796, 32'sd-0.015639884016805713, 32'sd0.12800743726252947, 32'sd0.04606152942144264, 32'sd0.07952328833487139, 32'sd0.1129995583022765, 32'sd0.07079228586679538, 32'sd0.07208198125242514, 32'sd0.10439384755441757, 32'sd0.08957802897239686, 32'sd0.13849793919039902, 32'sd0.072744028340598, 32'sd-0.020023225542124663, 32'sd0.0601504637667186, 32'sd0.06621495832884454, 32'sd0.06769639915171334, 32'sd-0.00306669840584822, 32'sd0.023228361964621243, 32'sd0.020179193904071357, 32'sd0.002608991792520453, 32'sd-0.09346851606089006, 32'sd0.05700897617776956, 32'sd-0.0431389527737135, 32'sd-0.1029684725694904, 32'sd-0.23982223767126087, 32'sd-0.07041906025654349, 32'sd0.025809158197725723, 32'sd0.06786566721739329, 32'sd-0.05997817825441177, 32'sd-0.013502757667264158, 32'sd-4.170674554628426e-123, 32'sd-0.0004555043476526156, 32'sd-0.010884387062255144, 32'sd-0.008110794980820967, 32'sd-0.042545738416197465, 32'sd-0.01140976657872196, 32'sd0.016643599008349722, 32'sd-0.038319359034060474, 32'sd-0.0226632950317543, 32'sd0.08615877740045931, 32'sd0.11692159533806445, 32'sd0.03143440766215414, 32'sd0.004748755806601189, 32'sd0.05966957758163995, 32'sd0.09795873056336607, 32'sd-0.0665525391332624, 32'sd0.06339483478939749, 32'sd-0.05069270134292185, 32'sd-0.050605560796201834, 32'sd-0.0793011957697152, 32'sd-0.025852032094071723, 32'sd-0.16580512856495214, 32'sd-0.18446238076804436, 32'sd-0.07829000871169475, 32'sd-0.06258967943468433, 32'sd-0.020203548508444844, 32'sd-0.053219162665815646, 32'sd0.054231581467141896, 32'sd0.08820042511667651, 32'sd0.07721265953073224, 32'sd-0.13834753196478827, 32'sd-0.06197538159753523, 32'sd-0.05596074514503057, 32'sd-2.970373392533962e-05, 32'sd-0.016026794632292705, 32'sd-0.051060388849708725, 32'sd0.029806873832200296, 32'sd0.06692224614399407, 32'sd0.029115156939942065, 32'sd-0.009514465977698673, 32'sd0.05541770037539215, 32'sd-0.022492400360129113, 32'sd-0.061761633567020316, 32'sd0.01684961684441847, 32'sd-0.006286671900933919, 32'sd0.05034479019914787, 32'sd0.10413878757443415, 32'sd0.02122128330421535, 32'sd-0.15266030970837527, 32'sd-0.1568028332803012, 32'sd-0.1188404189778827, 32'sd0.01263662222439967, 32'sd-0.04787934650826812, 32'sd-0.013586942155740668, 32'sd-0.1367697602432347, 32'sd0.03527474478246375, 32'sd0.07583542813045521, 32'sd0.12420301234090533, 32'sd-0.0625370080989773, 32'sd-0.08743484011158344, 32'sd-0.0163937279384947, 32'sd0.07443330689123626, 32'sd-0.04731366499499845, 32'sd-0.02289835663408279, 32'sd-0.11383233332163353, 32'sd0.031245704880952685, 32'sd0.009097151380766135, 32'sd-0.0013631580979029322, 32'sd0.049397831976032806, 32'sd-0.030449887202719676, 32'sd-0.01445811386573933, 32'sd0.0026093318415543318, 32'sd0.041488759091108586, 32'sd0.011430593268018882, 32'sd0.03425911250388362, 32'sd-0.0407869774976433, 32'sd-0.16364702647883686, 32'sd-0.04114694468850635, 32'sd-0.10427791708875217, 32'sd0.0011369482686338062, 32'sd-0.06148791628005916, 32'sd-0.03585801481565893, 32'sd0.059743917564955604, 32'sd0.07900036876213903, 32'sd-5.270618719599323e-124, 32'sd0.14083357919699963, 32'sd0.049008826214109985, 32'sd-0.005940953344840969, 32'sd0.09309002200866655, 32'sd0.017194048060412078, 32'sd-0.03959905610209974, 32'sd-0.041477088001110725, 32'sd-0.014883154775269615, 32'sd0.01620308403608509, 32'sd0.03860092228788982, 32'sd-0.022520658605064837, 32'sd0.06672600027443344, 32'sd0.020945486478280567, 32'sd0.11590685106086017, 32'sd0.08941672839522805, 32'sd-0.026594943282581395, 32'sd-0.09284655083740001, 32'sd-0.013053319033891278, 32'sd0.02283876839123424, 32'sd-0.025558944652866924, 32'sd8.040102989199324e-05, 32'sd0.02254942524761993, 32'sd0.05032364667112379, 32'sd0.012854550866250005, 32'sd0.04928402012883458, 32'sd-0.04007839643754387, 32'sd1.1659288810674111e-125, 32'sd7.1720009836922e-117, 32'sd7.05032372307732e-117, 32'sd0.0552507679029302, 32'sd0.005167085026175963, 32'sd-0.01271567651232989, 32'sd0.03767788426486869, 32'sd-0.02690551522988738, 32'sd0.03362867750081336, 32'sd-0.00458848913174832, 32'sd-0.002587786748160035, 32'sd-0.03313782024118852, 32'sd-0.030447871196688934, 32'sd-0.035587355296084804, 32'sd0.04940415369336912, 32'sd0.044661734346325824, 32'sd0.03617252070391267, 32'sd-0.04177742016751377, 32'sd0.07468570410062639, 32'sd-0.031004651106202923, 32'sd-0.03912884326137733, 32'sd-0.080847454609297, 32'sd0.02155322588917464, 32'sd-0.020344799338618245, 32'sd-0.07747417401018514, 32'sd0.04831652713034987, 32'sd0.049372111268666745, 32'sd-0.09295602089524635, 32'sd-2.847344423888579e-121, 32'sd-3.968457206524661e-121, 32'sd1.0165003451356074e-122, 32'sd0.13517711599070825, 32'sd0.08728194339047901, 32'sd0.038613204784286585, 32'sd-0.08242384662024024, 32'sd0.016571514489737073, 32'sd-0.020343301232016223, 32'sd-0.04276852960240478, 32'sd-0.003400913303881814, 32'sd0.0705935788739892, 32'sd-0.10604099886273395, 32'sd-0.008811550771119581, 32'sd0.061463347749125874, 32'sd-0.007816416686881973, 32'sd-0.06626902205707053, 32'sd0.08348106439325775, 32'sd0.06237068901530865, 32'sd0.0769037668666186, 32'sd0.0660880396776634, 32'sd-0.01099137332518286, 32'sd-0.059879231634678266, 32'sd-0.02032760918206247, 32'sd-0.09270654800762906, 32'sd0.054574616172329296, 32'sd0.14497435430776331, 32'sd0.08286523530775355, 32'sd3.828889461799924e-117, 32'sd1.7029402781403025e-124, 32'sd1.2725449072138525e-115, 32'sd5.085776114322293e-122, 32'sd0.1427406274005879, 32'sd0.041822272906979256, 32'sd0.04708356216686924, 32'sd0.059358937154563224, 32'sd0.024145428497051136, 32'sd-0.03974947266221172, 32'sd-0.023828096223253534, 32'sd0.012490063141320017, 32'sd-0.03101465829271486, 32'sd0.05396565634912541, 32'sd0.005093630033023574, 32'sd0.1382782835496079, 32'sd0.042508619607012285, 32'sd0.023990253170243465, 32'sd0.021433002732921546, 32'sd0.039370177016869706, 32'sd0.025482120226798213, 32'sd0.03865279529912281, 32'sd0.02882437684180953, 32'sd0.005490565163473304, 32'sd0.0328638736367157, 32'sd-0.008695800430310922, 32'sd0.15274711642019195, 32'sd-1.286851182129199e-115, 32'sd-3.9981263116357245e-125, 32'sd2.9172763412940694e-121, 32'sd-2.229969991856235e-122, 32'sd-1.0397902091175598e-120, 32'sd4.917268015189417e-117, 32'sd0.14510306904470205, 32'sd0.07573988739914149, 32'sd0.0439606040865279, 32'sd0.06935163286273686, 32'sd0.06808654015447292, 32'sd0.034767649625605544, 32'sd0.0202890977335385, 32'sd0.02978928609383903, 32'sd0.01185428928616467, 32'sd0.04770657384544596, 32'sd0.028508758688784965, 32'sd0.02863113287618538, 32'sd0.08616421146932235, 32'sd0.0092063623672877, 32'sd0.016491607836744276, 32'sd-0.043383204205568945, 32'sd0.04167160521091337, 32'sd-0.010349712348352089, 32'sd-0.06848863126250014, 32'sd0.12094690322498317, 32'sd1.3623313094782615e-125, 32'sd-3.672175309436913e-119, 32'sd-2.653758703335465e-124, 32'sd-7.533180461314758e-119},
        '{32'sd-1.3712565329273077e-125, 32'sd-1.6561142284653656e-123, 32'sd1.1801249567895654e-116, 32'sd1.4033308138523405e-117, 32'sd-8.616638018944867e-117, 32'sd-5.123028194430295e-122, 32'sd-8.800206210774711e-127, 32'sd-8.872296289283679e-116, 32'sd3.366964539794472e-120, 32'sd7.334349257450567e-123, 32'sd-6.355616319443889e-117, 32'sd2.4636241886310912e-124, 32'sd0.100049400841088, 32'sd0.03594856740699592, 32'sd0.08851327253678985, 32'sd0.028944525090140526, 32'sd5.308216511858657e-125, 32'sd1.414879066077605e-115, 32'sd1.7994113506361643e-114, 32'sd-8.62461241921953e-117, 32'sd-5.067088963770997e-118, 32'sd3.3489718323315974e-116, 32'sd1.3794362531023037e-125, 32'sd-1.0823972324338416e-121, 32'sd-8.306582603937813e-116, 32'sd7.231462275490555e-126, 32'sd2.5333241579808766e-124, 32'sd-4.782517093698648e-118, 32'sd-5.541260213423861e-122, 32'sd8.925875239519307e-121, 32'sd-1.109221139756348e-122, 32'sd1.6968030320993726e-125, 32'sd0.03587045439274204, 32'sd0.08016138228315209, 32'sd-0.06640494454937963, 32'sd0.08647874995649488, 32'sd0.038639370727954196, 32'sd0.0012537148959490645, 32'sd0.09747846062534334, 32'sd-0.03816286308910841, 32'sd0.07217344458394698, 32'sd0.05146523523277081, 32'sd0.12121252379563471, 32'sd0.07984300734433801, 32'sd0.07913145412722829, 32'sd0.05352521657891227, 32'sd0.08905299492078814, 32'sd0.0070147365648888915, 32'sd0.05626049418460399, 32'sd-0.010612164774727298, 32'sd0.03610897849092521, 32'sd0.021359234503694292, 32'sd1.869689277305852e-126, 32'sd2.3477593278544074e-118, 32'sd-2.0088632185596684e-116, 32'sd1.11709393166447e-119, 32'sd-2.191246975005418e-118, 32'sd-8.551715541334808e-121, 32'sd0.021638061871613, 32'sd0.028010072593585428, 32'sd0.11458019400571152, 32'sd-0.006269875502698821, 32'sd-0.03473744883457586, 32'sd-0.008160051518552367, 32'sd0.05959249722400349, 32'sd0.059287377816228254, 32'sd0.09744002694993158, 32'sd0.0608179634593557, 32'sd0.022336428122790977, 32'sd0.13881502351434508, 32'sd0.052965091939165626, 32'sd0.04456323108804109, 32'sd0.061789411306963915, 32'sd0.035466627365365475, 32'sd0.014897845003330471, 32'sd-0.0585512174913633, 32'sd0.11463473063024245, 32'sd0.0936081267777511, 32'sd0.08241640873922335, 32'sd-0.08964599907939144, 32'sd0.06371414099508346, 32'sd0.09491150525024641, 32'sd1.1391893222889854e-119, 32'sd-3.579626206203854e-123, 32'sd-2.7866132027031367e-127, 32'sd2.3681248030887443e-116, 32'sd0.06604146511785038, 32'sd0.11204402626541408, 32'sd0.0040726518506552754, 32'sd0.08545959241397662, 32'sd0.07281132792125954, 32'sd-0.03689465743078876, 32'sd0.11174118124909013, 32'sd0.026649735180377422, 32'sd-0.04559985536408753, 32'sd0.16922967591912422, 32'sd0.16212354010285557, 32'sd0.11414174092268549, 32'sd-0.11608875086963287, 32'sd-0.11526157072162305, 32'sd0.04323601939757327, 32'sd0.07719969635278348, 32'sd-0.01842850798195472, 32'sd-0.014201798591740464, 32'sd-0.04905410361243746, 32'sd-0.02382099689486093, 32'sd0.04010254894059964, 32'sd-0.08635937211255643, 32'sd0.00019836560538062566, 32'sd-0.037620463177724855, 32'sd0.009058989661405021, 32'sd-3.271397058216924e-120, 32'sd3.941260748863339e-129, 32'sd-0.005143022401378624, 32'sd-0.029064083551412215, 32'sd-0.06876540809972995, 32'sd0.0599694416026255, 32'sd-0.011262416498776294, 32'sd-0.009480469049851104, 32'sd-0.003938528661662116, 32'sd0.05326634664387643, 32'sd-0.08459218386664234, 32'sd-0.021800813456530774, 32'sd0.017589730315747797, 32'sd0.08439552524829536, 32'sd0.004856497014752451, 32'sd-0.014822234816702215, 32'sd0.02958536196957151, 32'sd-0.039615344933151005, 32'sd-0.05549117714150694, 32'sd-0.04040830983670436, 32'sd0.05355725396450956, 32'sd0.036825417358490986, 32'sd-0.10394890961740642, 32'sd-0.07120311777115478, 32'sd0.05376196224348758, 32'sd0.05796924799306997, 32'sd0.05296210965811531, 32'sd-0.13678046410729552, 32'sd0.026600149810607085, 32'sd-1.3977279328900027e-124, 32'sd0.007767522103344352, 32'sd0.06129620962772534, 32'sd0.046751019319135764, 32'sd0.022163071518834513, 32'sd-0.02726326225158418, 32'sd-0.0005327394588027202, 32'sd-0.0032062689934600373, 32'sd0.033482944871237444, 32'sd-0.031127401116112324, 32'sd0.0343803023536467, 32'sd-0.039295557461103976, 32'sd0.060864455883346213, 32'sd0.00018734877668719838, 32'sd-0.050594187560733445, 32'sd0.004610662563105975, 32'sd-0.004019244094458758, 32'sd-0.03350551958806817, 32'sd-0.15480440997535835, 32'sd-0.16273154588698832, 32'sd-0.11092913227476019, 32'sd0.0017414508457007816, 32'sd-0.15100878199224868, 32'sd0.05337735447006309, 32'sd0.09556852314870833, 32'sd0.08455052686858767, 32'sd-0.025722685154324763, 32'sd0.047308628381676494, 32'sd-2.067975941301961e-127, 32'sd-0.03167271114446419, 32'sd0.044764290470790634, 32'sd0.08428435613753667, 32'sd0.0561593498542617, 32'sd-0.05924197711047132, 32'sd-0.01985061942023515, 32'sd0.10277721138566025, 32'sd0.06862944332243116, 32'sd0.04651801048078483, 32'sd0.02257791489425014, 32'sd0.046684609825942074, 32'sd0.0886607945848156, 32'sd-0.05566285689859691, 32'sd-0.08241259688843705, 32'sd-0.22739417624559982, 32'sd-0.09865925254690185, 32'sd0.011917134457307962, 32'sd-0.07823150461689436, 32'sd-0.01732180239688441, 32'sd-0.11866243620500673, 32'sd-0.08635521463496722, 32'sd-0.10794175385984169, 32'sd-0.01328823202080839, 32'sd0.04185351020625271, 32'sd0.03205319722195644, 32'sd0.005757490275724564, 32'sd-0.02716853955719416, 32'sd0.04313894076424454, 32'sd0.0820680700432791, 32'sd0.04936833054803915, 32'sd-0.040449401329597574, 32'sd0.08697005910358822, 32'sd0.031228151745921202, 32'sd-0.02692778959766604, 32'sd0.045799688154551065, 32'sd0.00980916738571653, 32'sd0.07061342745591999, 32'sd0.09983576965613075, 32'sd0.0034321307372535536, 32'sd-0.039752731757655306, 32'sd-0.0975271345227287, 32'sd-0.12696397942990054, 32'sd0.005176331632054691, 32'sd-0.021266214163823384, 32'sd-0.09905062994634373, 32'sd0.09351828031515873, 32'sd0.10382761856889823, 32'sd0.009405516706967586, 32'sd0.017685019628762597, 32'sd0.039029273915566286, 32'sd-0.09574736754742579, 32'sd-0.07850846355676637, 32'sd-0.10999689493895241, 32'sd0.005419756003107, 32'sd0.027166800338213747, 32'sd0.024801490146016396, 32'sd0.0611256452156609, 32'sd0.04237655592322664, 32'sd0.017455466106240124, 32'sd0.09086700449784059, 32'sd-0.08908935416726523, 32'sd0.06662058006194926, 32'sd0.13964654400484441, 32'sd0.039109348092019124, 32'sd0.1469057859012314, 32'sd0.1423738314307972, 32'sd0.1896665469966443, 32'sd0.010782260567028067, 32'sd-0.21439201399422392, 32'sd-0.13993674639870704, 32'sd0.01645259991250895, 32'sd0.09659563363415112, 32'sd-0.0828570160168648, 32'sd0.07784260229109996, 32'sd-0.055183765245339515, 32'sd0.0753096739465495, 32'sd0.06321906481193887, 32'sd0.11670154213874116, 32'sd-0.024642315300027612, 32'sd0.033544206132347515, 32'sd-0.014519298753084612, 32'sd-0.0803120602670079, 32'sd0.009640072033565605, 32'sd0.01565833530012756, 32'sd-0.057000677013858185, 32'sd-0.07240723191541876, 32'sd0.049137665024692044, 32'sd0.08355792373598625, 32'sd0.012227129753956616, 32'sd0.07080792608505691, 32'sd0.08596668397825515, 32'sd0.12909038213292848, 32'sd0.047764217040708656, 32'sd0.021778041807910185, 32'sd0.034310270352144005, 32'sd-0.1297028746994787, 32'sd-0.1922236960644948, 32'sd-0.09604413576695629, 32'sd-0.07429941440953726, 32'sd0.03878486700371896, 32'sd0.06080381207746072, 32'sd0.16289342755303943, 32'sd0.009479782557953627, 32'sd0.14473427424687282, 32'sd0.11780759232170308, 32'sd0.04023688995391059, 32'sd-0.005202282669374698, 32'sd0.08360605735023574, 32'sd0.10339356727069396, 32'sd-0.03506509375166293, 32'sd-0.09637091856514048, 32'sd0.09863661002397373, 32'sd-0.050076529424777604, 32'sd-0.0027001654830617, 32'sd-0.042113356541588785, 32'sd0.1659487969501018, 32'sd0.12086460676054983, 32'sd-0.00028631183205370467, 32'sd0.016346672018241228, 32'sd0.08662270400899869, 32'sd-0.035341380148835304, 32'sd0.06787109337412985, 32'sd0.053421710104326545, 32'sd-0.06232737131651852, 32'sd-0.06481326694735458, 32'sd-0.1259614055552601, 32'sd-0.0514968719707374, 32'sd0.10316989876455111, 32'sd3.3534539609721545e-05, 32'sd0.237270304484593, 32'sd0.12047230699570495, 32'sd0.04231415315511972, 32'sd-0.031649534142470286, 32'sd0.050785532620923765, 32'sd0.08840254431613138, 32'sd0.16108332214200805, 32'sd0.08789699297464243, 32'sd-0.024231878499455954, 32'sd0.008025411519790478, 32'sd-0.004064802481617343, 32'sd-0.03427280177802498, 32'sd0.09216765704643007, 32'sd0.09371165673307275, 32'sd-0.01974713891662095, 32'sd0.09878951247928752, 32'sd0.0879198176071904, 32'sd0.05124949949830239, 32'sd0.12158201799315264, 32'sd0.21633611282227772, 32'sd0.04203616372790205, 32'sd-0.0006050284549700995, 32'sd-0.09856319141887063, 32'sd-0.17002867909584357, 32'sd-0.15172019232054804, 32'sd0.0246550418215323, 32'sd0.08467654760567393, 32'sd0.09421754995859734, 32'sd0.14287671272313807, 32'sd-0.00450704176938427, 32'sd0.01942482587296051, 32'sd-0.07456254695625843, 32'sd0.10691074182005608, 32'sd0.0626759849138314, 32'sd0.13711625861779456, 32'sd0.033888687196218875, 32'sd-0.09404784513886484, 32'sd-0.06319714292840334, 32'sd0.07330976985216134, 32'sd0.03791977052688559, 32'sd0.06491961673857871, 32'sd-0.0818783154353201, 32'sd-0.023748704552338594, 32'sd0.08093219027998175, 32'sd-0.08690373621849964, 32'sd0.09057321142184196, 32'sd0.23222489026208507, 32'sd0.13510489600812345, 32'sd0.030405911172223094, 32'sd-0.05699560057293962, 32'sd-0.1424741718358898, 32'sd-0.09031077129128438, 32'sd-0.133152487839295, 32'sd-0.12281534038932967, 32'sd-0.07539442807160146, 32'sd0.09058382922742209, 32'sd0.0013227899747196882, 32'sd-0.026032876102621175, 32'sd0.019653366162270734, 32'sd0.015674844979490975, 32'sd0.015428031660744456, 32'sd0.03775104293679968, 32'sd0.1622331785870172, 32'sd0.0017607255428725196, 32'sd-0.08038787572821583, 32'sd-0.0033237003672492212, 32'sd0.029150115832511092, 32'sd-0.033178552673799995, 32'sd-0.07855588343285011, 32'sd-0.010302583291296784, 32'sd-0.014637158857926562, 32'sd0.10672597978872773, 32'sd0.1110106087287805, 32'sd0.15959695648075944, 32'sd0.10265709836079996, 32'sd0.14624375194245062, 32'sd0.11622500327255302, 32'sd-0.09656909518995112, 32'sd-0.18785847776211015, 32'sd-0.15258725133612414, 32'sd-0.18546899681828208, 32'sd-0.12211252139073966, 32'sd-0.07489457737194041, 32'sd0.09074359673558625, 32'sd0.04062389414739227, 32'sd0.004367264571563151, 32'sd0.04744629769170351, 32'sd0.08315947681405708, 32'sd-0.0030686988245107977, 32'sd0.08212407269419357, 32'sd0.03983458258044547, 32'sd0.020833317280489594, 32'sd0.028228164742623914, 32'sd0.05299470656302286, 32'sd-0.020919458514160993, 32'sd-0.007296190618306638, 32'sd0.0165026715333367, 32'sd0.04552804012989141, 32'sd-0.012859997589422339, 32'sd-0.018159487203721618, 32'sd0.06434314535211039, 32'sd0.1191576997594482, 32'sd0.039100731545338066, 32'sd0.041825311845034616, 32'sd-0.0028697931079261175, 32'sd0.0352591698552775, 32'sd-0.1049769095127965, 32'sd-0.16660213066277527, 32'sd-0.18337882909439948, 32'sd-0.1949322016801265, 32'sd0.16533637307242363, 32'sd0.14254741180328684, 32'sd0.1733680576963579, 32'sd0.03791415519748403, 32'sd0.07289223993151522, 32'sd0.11242233556767846, 32'sd0.09737088700083167, 32'sd0.0673738610758418, 32'sd-0.05166442236899953, 32'sd0.05034525563414478, 32'sd0.006114630947348745, 32'sd0.0402242137218466, 32'sd0.02835405664266943, 32'sd-0.05188058063887327, 32'sd-0.15593143543330326, 32'sd0.067050544806253, 32'sd-0.021097707501085153, 32'sd-0.023538858731235835, 32'sd0.0024011420344889896, 32'sd0.15221537177494238, 32'sd0.10052545771431967, 32'sd-0.013253955367021382, 32'sd-0.07434344142790615, 32'sd-0.034681765840680806, 32'sd-0.13068062076231304, 32'sd-0.08512880497925261, 32'sd-0.20052238485816226, 32'sd-0.011805147292058818, 32'sd0.03518041314908982, 32'sd0.10504368377776993, 32'sd0.06132954808269808, 32'sd0.049182140226097175, 32'sd0.06071341541893462, 32'sd-0.02635486035755185, 32'sd0.08041268934415813, 32'sd0.1037142001406538, 32'sd-0.09476965824522392, 32'sd0.09807941110808378, 32'sd-0.05621030130590258, 32'sd0.007229956806917818, 32'sd0.034387211977228944, 32'sd0.03661311410513663, 32'sd-0.07029674359184211, 32'sd0.05492149789640613, 32'sd0.03191969844810595, 32'sd0.0998551194130805, 32'sd0.05897774993573355, 32'sd0.09414977609419553, 32'sd0.10166474244024915, 32'sd-0.11475527044138978, 32'sd0.002054246799763032, 32'sd-0.03852952103538695, 32'sd-0.03367975882394517, 32'sd-0.14487281078964576, 32'sd-0.11679869539434705, 32'sd-0.004859947876013479, 32'sd0.06808366065827529, 32'sd0.26573764384031895, 32'sd0.12688524621848435, 32'sd0.03002860949130241, 32'sd0.07936373865298021, 32'sd0.05972078937757336, 32'sd-0.05489289153727521, 32'sd0.04989267423849923, 32'sd-0.029552301120166685, 32'sd0.038103254017062396, 32'sd0.024929047695231344, 32'sd-0.025804725855211385, 32'sd1.4791233907382385e-115, 32'sd0.0049671447585798376, 32'sd0.07155590264984985, 32'sd-0.006281925946856764, 32'sd0.027419475221863245, 32'sd0.031804718595044565, 32'sd0.016861654291993395, 32'sd0.06600105501100217, 32'sd0.03165412637447565, 32'sd0.06357549913632088, 32'sd-0.046230656538159824, 32'sd-0.06745860638037245, 32'sd-0.1521733814618994, 32'sd-0.20831985844084352, 32'sd0.044432885527869864, 32'sd0.009743578541679242, 32'sd0.23967646657112238, 32'sd0.1838037985694382, 32'sd0.10209904057541559, 32'sd-0.020223725237957083, 32'sd-0.12984147810699445, 32'sd-0.01154801320370904, 32'sd0.10589244988982542, 32'sd0.017987421846399298, 32'sd-0.010227421067263239, 32'sd-0.027978640335231515, 32'sd-0.03858075324134123, 32'sd-0.005643213456982571, 32'sd0.006836009569393638, 32'sd-0.0798314698174276, 32'sd0.09453932275825222, 32'sd-0.1309971418077066, 32'sd-0.01345932113500853, 32'sd0.008301461328104814, 32'sd-0.04556216921671308, 32'sd-0.009730895237632188, 32'sd-0.008477615276562914, 32'sd0.09925979923049273, 32'sd-0.01700419371099611, 32'sd-0.13610287188942571, 32'sd-0.26909877152421596, 32'sd-0.04725914568825826, 32'sd0.023361535437865708, 32'sd0.13320718067019574, 32'sd0.21012343018445473, 32'sd0.1374969731163937, 32'sd0.08398036970407596, 32'sd-0.10234832366968265, 32'sd-0.11834012483282644, 32'sd-0.07539955020168962, 32'sd0.041488430298767316, 32'sd-0.057169752286052, 32'sd0.08216031744711161, 32'sd0.08546188908746735, 32'sd0.027593584113651766, 32'sd0.03416305892212422, 32'sd0.042688193158715734, 32'sd0.08710533145643982, 32'sd-0.023913373971933855, 32'sd-0.0901256100620938, 32'sd-0.08174224593266953, 32'sd-0.026861588599723624, 32'sd0.0053036207625182215, 32'sd0.08728628204527042, 32'sd0.05368943924105128, 32'sd0.0655893148639192, 32'sd0.03402314624639419, 32'sd-0.09152049995570591, 32'sd-0.28839736133728583, 32'sd-0.20668401074828763, 32'sd0.02061714905437563, 32'sd0.15153571499413673, 32'sd0.21512030906568802, 32'sd0.08317781305719442, 32'sd0.07380147120146673, 32'sd0.07935732472395678, 32'sd0.033067341441323096, 32'sd-0.13485820812502308, 32'sd0.037269237438636645, 32'sd0.03995762602231808, 32'sd0.049693156284367684, 32'sd0.03582711105414193, 32'sd-0.012914099205583597, 32'sd-0.08974638357719422, 32'sd-1.104133890025985e-121, 32'sd-0.007499918029380765, 32'sd0.11063445346514411, 32'sd-0.02028491417922956, 32'sd-0.06997654456047508, 32'sd0.10063233768388746, 32'sd-0.03632251371862516, 32'sd-0.007545921085087512, 32'sd0.1098124312975856, 32'sd0.05757819011114307, 32'sd-0.05405838640421122, 32'sd-0.12382950987626176, 32'sd-0.11367375015100072, 32'sd-0.14246917192462877, 32'sd0.03807118496801879, 32'sd0.20606932342561313, 32'sd0.21719357021987143, 32'sd-0.04880880617654919, 32'sd0.06974854102891168, 32'sd0.030347474610130595, 32'sd-0.07446043026462999, 32'sd-0.1119750626553082, 32'sd-0.031495998720689686, 32'sd-0.09150491723220375, 32'sd0.06982792487799708, 32'sd0.07112905579229621, 32'sd-0.12452311759125749, 32'sd-0.01822673325105161, 32'sd0.035054692694188164, 32'sd0.019698622900804902, 32'sd-0.038065500471857944, 32'sd-0.09534392954843367, 32'sd-0.12659214633068055, 32'sd0.0925280143704681, 32'sd-0.06377922083933144, 32'sd-0.05685939730481868, 32'sd0.06260592884328398, 32'sd0.04394111992323426, 32'sd0.11523874243030398, 32'sd0.008903641715347533, 32'sd-0.107088260168313, 32'sd-0.05862716373443641, 32'sd0.05501201600427842, 32'sd0.16947313358090446, 32'sd0.13630176050744222, 32'sd0.1273878721714897, 32'sd-0.028377510063688584, 32'sd-0.041723973583933927, 32'sd-0.07028604230628444, 32'sd-0.07112841548329855, 32'sd0.006991598540936378, 32'sd-0.007988222173471657, 32'sd0.036261753290574156, 32'sd-0.03832609203278767, 32'sd-0.006055546610285397, 32'sd0.08362080896146182, 32'sd0.009559460691918814, 32'sd-0.014388020119317788, 32'sd-0.03595628834636046, 32'sd0.02036738497215601, 32'sd-0.07192855714572526, 32'sd0.08793125620717103, 32'sd0.039839611659343674, 32'sd0.02517621000147931, 32'sd-0.014115239749165934, 32'sd0.08928718528796085, 32'sd-0.08012949278214403, 32'sd-0.06074228921920811, 32'sd-0.16500203666225474, 32'sd-0.057320522153548104, 32'sd0.03718909061185394, 32'sd0.21206674183191174, 32'sd0.14836081490249112, 32'sd0.09692013260924605, 32'sd-0.11574313514532278, 32'sd0.01800342671900156, 32'sd0.031087699553629635, 32'sd0.009605141760464519, 32'sd0.003946071740713464, 32'sd-0.20026458356380963, 32'sd-0.06278309486203158, 32'sd-0.05487654746277896, 32'sd-0.09386378260234464, 32'sd-0.026902370985584498, 32'sd-2.581764529384762e-126, 32'sd0.06637631507153287, 32'sd-0.06721367229358685, 32'sd0.011208011337646007, 32'sd-0.056767556594749954, 32'sd0.003764235554305657, 32'sd0.0778658304782511, 32'sd0.057160830613768546, 32'sd0.14987825742392918, 32'sd0.017593597134934066, 32'sd-0.03494443787775422, 32'sd-0.21706583432792373, 32'sd-0.1415031363645248, 32'sd-0.02777072951259945, 32'sd0.1805868400915578, 32'sd0.1278739285253091, 32'sd0.15940086296511163, 32'sd0.1300045676648292, 32'sd-0.13624247664183275, 32'sd-0.09511381611096134, 32'sd-0.021770873915289524, 32'sd0.030344450667949333, 32'sd-0.10524208818145017, 32'sd0.020872479344694668, 32'sd-0.016693090940224475, 32'sd0.03581296573529429, 32'sd-0.0039152359497007, 32'sd9.212145202612831e-122, 32'sd-2.7715668790647398e-117, 32'sd-1.3068333789956855e-116, 32'sd0.03351742529492505, 32'sd-0.005767860092732752, 32'sd0.009051993731633701, 32'sd-0.04576287223259598, 32'sd-0.031309208386792915, 32'sd0.024743857733029, 32'sd0.05184408613279932, 32'sd0.09293397318228411, 32'sd-0.09003120309949238, 32'sd-0.19519360150576853, 32'sd-0.18219500918248813, 32'sd-0.09383858388623523, 32'sd-0.03193033707829954, 32'sd0.01848606612621632, 32'sd0.021805319718940716, 32'sd0.046858313532164055, 32'sd-0.020496406878592752, 32'sd-0.0011321384816151089, 32'sd0.11668099964566915, 32'sd-0.03236174893183755, 32'sd-0.04575881104347632, 32'sd-0.005683503660103599, 32'sd-0.10691720198562345, 32'sd0.0016461493110161319, 32'sd0.040725834658213014, 32'sd-1.8993030118737634e-124, 32'sd-1.0071836361088461e-118, 32'sd-4.797136264169181e-119, 32'sd-0.05144676814452969, 32'sd-0.018850121858089906, 32'sd-0.09728953263227676, 32'sd-0.014566799597471085, 32'sd0.07037184895518069, 32'sd0.07523992025068635, 32'sd-0.013282149779796248, 32'sd0.033721221367036945, 32'sd-0.13496523461033288, 32'sd-0.15745875018590325, 32'sd-0.0432753146020681, 32'sd-0.06396618847823239, 32'sd0.04424300992647582, 32'sd0.033733575516500414, 32'sd0.12289640860448768, 32'sd0.12741608916608593, 32'sd0.03032031662295318, 32'sd-0.023874320629185302, 32'sd0.03157487374978235, 32'sd0.1451755860151814, 32'sd-0.028407797680740542, 32'sd-0.052218731761683186, 32'sd0.05160982342772785, 32'sd0.05843408459039886, 32'sd-0.006882383794136196, 32'sd-2.2507105008871926e-122, 32'sd-8.625754126585027e-117, 32'sd-3.538720343765689e-122, 32'sd-3.152310635097309e-120, 32'sd0.018430914705346742, 32'sd-0.037237027033108425, 32'sd0.008825623703739191, 32'sd0.043248410314441356, 32'sd0.07484159346124351, 32'sd0.036880665785501754, 32'sd-0.030347940665907434, 32'sd-0.09966346691782667, 32'sd0.01064662313024579, 32'sd0.014650041761999136, 32'sd0.023809526417550676, 32'sd0.06890573489137329, 32'sd0.03919262382592622, 32'sd0.05248556357210149, 32'sd-0.03252460746175294, 32'sd-0.05296938730210005, 32'sd0.025698055777844123, 32'sd-0.09014724751410602, 32'sd0.07454907120482022, 32'sd0.08241715480488579, 32'sd0.04763202626747872, 32'sd-0.017132081684488064, 32'sd-0.017454965560980303, 32'sd-2.38969210602034e-123, 32'sd-2.711905510246925e-122, 32'sd-1.0512857975827621e-119, 32'sd1.7106630334461927e-124, 32'sd2.150510289397217e-119, 32'sd-1.066425591807054e-124, 32'sd0.08559758966695855, 32'sd0.05045596890215687, 32'sd0.01796448940436926, 32'sd0.06680955285028554, 32'sd0.01615063220627287, 32'sd0.01065548448279767, 32'sd-0.10528621438872383, 32'sd0.048361832327652746, 32'sd-0.05712724569411128, 32'sd0.06829973782509312, 32'sd0.04331903257297865, 32'sd-0.04754562168727294, 32'sd0.046718282110124944, 32'sd0.010755219058838613, 32'sd0.08311769269650783, 32'sd-0.021272028709392175, 32'sd-0.06877931195809009, 32'sd-0.0021386553968010978, 32'sd0.008598636530962024, 32'sd-0.07120087266503768, 32'sd5.103388580878198e-117, 32'sd-2.0243721299800324e-120, 32'sd-6.218330254873859e-124, 32'sd4.960040537018038e-118},
        '{32'sd-1.3416029004754395e-125, 32'sd2.4033741212878226e-118, 32'sd1.469552373332914e-121, 32'sd-4.509490364518907e-115, 32'sd7.33560326297239e-123, 32'sd8.022991240147913e-123, 32'sd1.4988135770110625e-127, 32'sd7.221358279529356e-120, 32'sd-2.4924259647686264e-121, 32'sd-8.717097594924414e-127, 32'sd-3.040664170010366e-115, 32'sd4.454866091537579e-124, 32'sd0.036060728912055764, 32'sd-0.04203196690132192, 32'sd0.004075097400314935, 32'sd-0.03595030401321841, 32'sd8.502022529735255e-129, 32'sd1.4470192048691876e-123, 32'sd-3.117211273695037e-116, 32'sd-6.217023392804148e-119, 32'sd-1.1372763425049858e-119, 32'sd-1.7431089272311738e-123, 32'sd-5.819303582561843e-121, 32'sd-6.556393051666626e-117, 32'sd-2.4753703181044298e-123, 32'sd1.3748175495163941e-123, 32'sd-8.224925132472116e-127, 32'sd-5.944548151002018e-126, 32'sd1.0620523006706616e-121, 32'sd7.192784796696529e-126, 32'sd-1.387401757419685e-122, 32'sd-5.119095700579489e-123, 32'sd-0.045450105860604086, 32'sd0.07996806091625676, 32'sd0.0628538007284979, 32'sd-0.10240613620322071, 32'sd0.053317004294641805, 32'sd0.02393157030808581, 32'sd0.01399284178894982, 32'sd0.06355953740598301, 32'sd-0.06949758548056703, 32'sd-0.0515165807471855, 32'sd0.03699490766696889, 32'sd0.06018282381356319, 32'sd-0.025870107449380623, 32'sd0.007699894328117684, 32'sd-0.011916154805030395, 32'sd-0.01592708935808416, 32'sd0.02016254810743657, 32'sd0.0509646665512383, 32'sd0.02884237068134612, 32'sd0.03901220836688472, 32'sd-1.6807662880330305e-125, 32'sd-2.6108823771801927e-119, 32'sd4.73434169556334e-125, 32'sd2.354380809836615e-123, 32'sd-3.38956057659186e-120, 32'sd-6.892078938299815e-126, 32'sd0.09601159071404197, 32'sd0.03218041932417454, 32'sd-0.04823090031200019, 32'sd0.0678807630295094, 32'sd0.020946293234439937, 32'sd-0.0515198094444157, 32'sd0.018337026649996934, 32'sd-0.021962650958348272, 32'sd-0.015625604251250147, 32'sd0.07527695091919, 32'sd0.11369304656622366, 32'sd0.1553527641114968, 32'sd-0.06935835935002319, 32'sd0.04788341465186006, 32'sd0.11296619722831952, 32'sd-0.09709480823219371, 32'sd-0.03465518317553977, 32'sd0.10274651105886726, 32'sd0.05919884159105816, 32'sd-0.0620743758020501, 32'sd0.019899278654867368, 32'sd0.025479281146994343, 32'sd0.0568990238034914, 32'sd0.026177008374441105, 32'sd1.2018201231687934e-122, 32'sd-2.4325456104757665e-121, 32'sd5.900152769587158e-115, 32'sd-8.636552554596308e-117, 32'sd0.09797917716807768, 32'sd-0.0280662102817485, 32'sd0.03262686391556432, 32'sd-0.019031298250899876, 32'sd0.07990444994613721, 32'sd-0.04197352517540853, 32'sd-0.010150976025334197, 32'sd0.04068213996712768, 32'sd0.13342809465741792, 32'sd0.05910399887234542, 32'sd0.2113472723913841, 32'sd0.15129813692730296, 32'sd0.027037566078817375, 32'sd0.04515076270930119, 32'sd0.11967302939097338, 32'sd-0.05021312418003206, 32'sd-0.11388099412690406, 32'sd-0.12801751372157835, 32'sd0.06809583092271436, 32'sd0.023240842646529675, 32'sd-0.017151603055576916, 32'sd-0.05217917985237709, 32'sd0.040965388570291736, 32'sd-0.028554464128170892, 32'sd0.043339750130647475, 32'sd-2.412827172180715e-124, 32'sd-6.103935231324637e-125, 32'sd0.054342268757503115, 32'sd-0.06174682084924303, 32'sd-0.04694481909946822, 32'sd-0.02763400300832109, 32'sd0.05809267088817864, 32'sd-0.052651842196048945, 32'sd-0.08371220086676338, 32'sd-0.05972191325404614, 32'sd0.165136655170625, 32'sd0.07600493231296826, 32'sd0.08736627498149982, 32'sd0.16630796527566702, 32'sd0.040079852081135264, 32'sd0.07429924700426183, 32'sd0.05418201209347102, 32'sd-0.04315694893569083, 32'sd0.03431495642783336, 32'sd-0.04092742922680013, 32'sd-0.1076289920415041, 32'sd-0.013241941951607623, 32'sd0.056002029394342706, 32'sd0.07167062265454985, 32'sd-0.09801814126692916, 32'sd-0.04898178945769353, 32'sd-0.09444637514566255, 32'sd-0.007542951887898947, 32'sd0.02826134736689936, 32'sd1.8252154399720342e-127, 32'sd0.02803667262377005, 32'sd0.0181337479693279, 32'sd-0.02076789277614354, 32'sd0.015230589146499638, 32'sd-0.053375485184156427, 32'sd0.03777088757519328, 32'sd-0.03733542434665336, 32'sd0.05189553455373798, 32'sd0.012716435085712177, 32'sd0.07289921415167026, 32'sd0.09158959803766792, 32'sd-0.007236960071051814, 32'sd0.06784304584532011, 32'sd0.15045013789078732, 32'sd0.08443902102124778, 32'sd0.0029968315203455936, 32'sd-0.010095519336829815, 32'sd0.07783366507963589, 32'sd0.025388811954132146, 32'sd-0.010677527968350892, 32'sd-0.030654714312972987, 32'sd0.05447053852340994, 32'sd-0.03719913490890636, 32'sd0.005440193565485347, 32'sd0.031927332954513915, 32'sd-0.08873671251420129, 32'sd0.010333051230365603, 32'sd-7.930651511204458e-116, 32'sd0.05571617637689071, 32'sd0.02897456900411987, 32'sd0.10479919926582447, 32'sd-0.04173355856957336, 32'sd-0.0012228220812367345, 32'sd-0.04748789174367608, 32'sd-0.07947548041753372, 32'sd0.037027517902698884, 32'sd-0.026441640122466713, 32'sd0.057012035090486066, 32'sd-0.04092557910375854, 32'sd0.06604346076805423, 32'sd0.04462413088767834, 32'sd0.051369010590599354, 32'sd0.13110046304350936, 32'sd0.11948192393453648, 32'sd-0.004520076383838318, 32'sd0.08528808041978182, 32'sd-0.02818638633745265, 32'sd-0.022028959643965337, 32'sd0.0193133491651324, 32'sd-0.03458674311401869, 32'sd-0.0937034482346898, 32'sd0.038635949372173926, 32'sd0.14048577522558944, 32'sd0.02810281700857367, 32'sd-0.03449404153109157, 32'sd0.06075337849863039, 32'sd0.06049763914780137, 32'sd0.060254411043475446, 32'sd0.10391735817825855, 32'sd-0.06283347427189684, 32'sd-0.008289135175575786, 32'sd-0.062263938924883605, 32'sd-0.060494555031561044, 32'sd-0.10051910497646921, 32'sd0.01644603777135838, 32'sd-0.004458219849410048, 32'sd0.09716289077690378, 32'sd0.08894280422285979, 32'sd0.05605540633061301, 32'sd0.04647131847833874, 32'sd0.0907479565241774, 32'sd0.1598768044545557, 32'sd0.16051364227519924, 32'sd0.011565875735142951, 32'sd0.1833544332173413, 32'sd0.061087276117957806, 32'sd-0.025853544434697714, 32'sd-0.031152341435623565, 32'sd0.013768299420283603, 32'sd0.05426218306450227, 32'sd-0.01501501594349423, 32'sd-0.03704336931192898, 32'sd0.034567790978895924, 32'sd0.058692952714516, 32'sd0.05821353534021222, 32'sd0.028921852775918546, 32'sd-0.09411831052521794, 32'sd-0.030356622620945888, 32'sd0.07168994107441544, 32'sd-0.05257687729428505, 32'sd-0.05279745769514906, 32'sd-0.013076999728763715, 32'sd-0.1042295250741095, 32'sd0.025845530101128843, 32'sd0.01945237172403317, 32'sd0.04554703320491677, 32'sd0.1307578326653115, 32'sd0.12187281805198569, 32'sd0.10544277541869068, 32'sd0.09068335296093322, 32'sd0.10943300321772378, 32'sd0.11674277160198078, 32'sd-0.0030588370243071154, 32'sd0.14409041717308824, 32'sd0.0973312541810098, 32'sd0.11043173715208088, 32'sd0.04556064031275965, 32'sd0.03293822714536602, 32'sd0.013709728952841092, 32'sd-0.00915141426635725, 32'sd-0.08385066460504136, 32'sd0.06469856097934604, 32'sd-0.07565738668505871, 32'sd-0.11413380313513258, 32'sd-0.002881171631032847, 32'sd0.004592768009548127, 32'sd-0.08312207007514985, 32'sd-0.12812950826999792, 32'sd-0.0042956044556450666, 32'sd-0.01900292093885441, 32'sd-0.022538688602129684, 32'sd-0.07561005352968841, 32'sd-0.0009578052330259738, 32'sd0.023170825193387368, 32'sd0.11466666944688923, 32'sd0.14843925172597533, 32'sd0.10399396292984459, 32'sd0.09020875242909503, 32'sd-0.09967752492292467, 32'sd-0.08655994705756397, 32'sd0.002450383190223098, 32'sd0.046297203526769845, 32'sd0.03531680520270105, 32'sd0.0374463356885398, 32'sd0.05286268030815042, 32'sd0.10387556134858628, 32'sd0.09887981665934674, 32'sd-0.024157064254893407, 32'sd0.04670582113332159, 32'sd-0.03740254840921299, 32'sd0.0007112713543858637, 32'sd-0.07389583333441109, 32'sd-0.17786808829213516, 32'sd-0.00219853986775377, 32'sd-0.067637297778731, 32'sd-0.05403705529266553, 32'sd-0.10058167020131677, 32'sd-0.04212834630172008, 32'sd0.06148857633170103, 32'sd-0.08582054917585506, 32'sd0.029953378539716115, 32'sd0.08460981686180279, 32'sd0.12553833664844355, 32'sd0.06650408283601597, 32'sd0.0067076736887332865, 32'sd0.03826205066508419, 32'sd-0.0438837345924828, 32'sd-0.1468014672735425, 32'sd-0.06697549056471733, 32'sd-0.022929826543691585, 32'sd-0.06820864014292613, 32'sd0.040954875938018005, 32'sd0.05627889606444948, 32'sd0.09927681302049045, 32'sd-0.15485753372722327, 32'sd-0.08214061865460028, 32'sd0.07389494668862737, 32'sd0.04457317680259066, 32'sd0.02932697482786686, 32'sd-0.019492584399282913, 32'sd0.0744064278508835, 32'sd0.022806450537229555, 32'sd-0.07237991390576816, 32'sd0.04326234145862143, 32'sd-0.006021693189979193, 32'sd-0.09184614476569053, 32'sd-0.12863247978727885, 32'sd0.09986029071534432, 32'sd0.08209169966447864, 32'sd0.18081243273902992, 32'sd0.14592464739872452, 32'sd0.0127387665328929, 32'sd-0.031264572012397955, 32'sd0.009887856323139975, 32'sd-0.09063194426963882, 32'sd0.09709751534841131, 32'sd-0.016621799021478444, 32'sd-0.08316653724646522, 32'sd-0.16799881922687748, 32'sd-0.08532761724573129, 32'sd-0.07515635897447788, 32'sd0.00021863524991544458, 32'sd-0.09668182836866532, 32'sd-0.006458827639381775, 32'sd0.05590237355740281, 32'sd-0.002642529820875546, 32'sd-0.016261941024458493, 32'sd-0.04762351084858044, 32'sd0.05048593666353765, 32'sd0.06372300079328125, 32'sd-0.001975060537585895, 32'sd0.08580585012275746, 32'sd0.04183674524166829, 32'sd0.04175428727388205, 32'sd0.014521108946487917, 32'sd-0.016140513609274196, 32'sd0.06515014255210193, 32'sd0.15397778692916844, 32'sd0.1499842861983141, 32'sd0.035565647143743696, 32'sd0.008272852971248842, 32'sd0.01402774691377386, 32'sd-0.04237724544046594, 32'sd0.08016451080412647, 32'sd0.061805770613080534, 32'sd-0.07041283098349346, 32'sd-0.057081136356086394, 32'sd-0.050382413522884625, 32'sd0.013905664091858026, 32'sd-0.06629332456019087, 32'sd-0.07820343857583387, 32'sd-0.05429686588539907, 32'sd0.11241951478849418, 32'sd0.04788560387510597, 32'sd-0.002632554224363482, 32'sd0.01227697641980057, 32'sd0.1479300326302539, 32'sd0.13183893302885333, 32'sd-0.07591068965332372, 32'sd0.005341269626132739, 32'sd0.05223274778787993, 32'sd0.1051367519304189, 32'sd-0.05757682913962418, 32'sd0.04409313246235999, 32'sd0.04423825733049296, 32'sd0.011594899452788868, 32'sd0.0513181056665954, 32'sd0.03606449116294014, 32'sd-0.01047067505950927, 32'sd0.12744366364953819, 32'sd0.08049135147028608, 32'sd0.16789441816623996, 32'sd0.07521672661291656, 32'sd-0.05371039034778494, 32'sd-0.07336787578585577, 32'sd-0.07298364176046185, 32'sd0.0017556141065188542, 32'sd-0.04087227543192629, 32'sd-0.05012869250706366, 32'sd-0.029515843011549008, 32'sd0.07538622395278102, 32'sd0.06565327397651752, 32'sd-0.007658373763053619, 32'sd-0.09748368962748781, 32'sd-0.0273592903203939, 32'sd0.07295215447075216, 32'sd-0.13520853086333265, 32'sd-0.03349758945002998, 32'sd-0.02516120974942931, 32'sd-0.015542201163650895, 32'sd-0.034095130674703544, 32'sd-0.11869642297716086, 32'sd-0.10848553271486586, 32'sd0.056856249778715603, 32'sd-0.0076096807135506124, 32'sd0.07226741234999909, 32'sd-0.02368809780639007, 32'sd-0.012004921134160743, 32'sd-0.05102036039622538, 32'sd0.08532398273001718, 32'sd0.10273308310940545, 32'sd0.046922603007017304, 32'sd-0.02988546299533725, 32'sd-0.029791445734625985, 32'sd0.0950042414754995, 32'sd0.03848265169500004, 32'sd-0.04164261586757268, 32'sd-0.06735851544415318, 32'sd0.06404921848311662, 32'sd0.07035720462383951, 32'sd0.025058240110890383, 32'sd0.040798211397988074, 32'sd-0.025676257959493406, 32'sd0.08523259846923759, 32'sd-0.14954661245205159, 32'sd-0.18160284591530332, 32'sd-0.20081110013329082, 32'sd-0.27933252691744764, 32'sd-0.3540873650873, 32'sd-0.2416966046203812, 32'sd-0.06250145086173944, 32'sd0.04617664339154822, 32'sd-0.11954394617463723, 32'sd-0.03948750383407903, 32'sd-0.06942882475903384, 32'sd-0.017468039157603994, 32'sd-0.03214509456581718, 32'sd0.11130492756424373, 32'sd0.000527857396470217, 32'sd0.0965877535262935, 32'sd0.13688231967980347, 32'sd0.14979006418843802, 32'sd0.00037404424934441233, 32'sd0.011643309750649896, 32'sd0.11872659056348098, 32'sd0.008336785317360026, 32'sd0.028105359737319986, 32'sd0.05202247340481292, 32'sd0.06889806854121908, 32'sd0.0209240977938954, 32'sd0.04703706730279218, 32'sd0.07461222944939645, 32'sd-0.05327474570884705, 32'sd-0.06855391518358267, 32'sd-0.02103450322541313, 32'sd-0.30220358865557956, 32'sd-0.26421987840173466, 32'sd-0.1896312092995249, 32'sd-0.1532680521847218, 32'sd-0.08065443601539653, 32'sd-0.12060959447977876, 32'sd-0.043234641812512194, 32'sd-0.03989993413095607, 32'sd-0.007490007629444944, 32'sd0.06707502608519725, 32'sd0.11533324041597827, 32'sd0.06081133101664204, 32'sd0.1476175523156519, 32'sd0.18663575756598907, 32'sd0.17791721457082055, 32'sd-0.014413613275715716, 32'sd-0.009373075692716226, 32'sd-0.15363379507070263, 32'sd-0.026832379161370733, 32'sd0.052602657439520015, 32'sd-3.239143731173666e-116, 32'sd0.01067743888293548, 32'sd-0.03340560373745715, 32'sd-0.031490741038887334, 32'sd0.08825661306459771, 32'sd0.07819915718414659, 32'sd-0.04865837713391752, 32'sd0.0717254647790216, 32'sd-0.003927545382188453, 32'sd-0.11048992484137968, 32'sd-0.14496153622867897, 32'sd-0.05945640725180276, 32'sd-0.11327836041170468, 32'sd-0.07197983612413054, 32'sd-0.0202975866108413, 32'sd-0.06742789265231662, 32'sd-0.08093161363140237, 32'sd0.08189929224598597, 32'sd0.06444912520443682, 32'sd0.008111235890969105, 32'sd0.15606703540935946, 32'sd0.1467955828947477, 32'sd-0.006579893941668596, 32'sd-0.09992584367361386, 32'sd-0.036124931386745635, 32'sd-0.15027177327630212, 32'sd0.032614215482801, 32'sd-0.020857916753467428, 32'sd0.026919872990212267, 32'sd-0.0004134434763954267, 32'sd-0.009220209273310647, 32'sd0.030077528423099038, 32'sd0.1279971635754824, 32'sd0.09681869098527106, 32'sd0.13920135438741305, 32'sd0.11982029197347034, 32'sd0.1223399356011008, 32'sd0.055577402747499435, 32'sd-0.01927471885261425, 32'sd0.07900175554707055, 32'sd-0.11593692099004102, 32'sd-0.12983287561246543, 32'sd-0.13814687641536938, 32'sd-0.05401686082073204, 32'sd0.023617920012734103, 32'sd0.05483992746924171, 32'sd-0.047157694893322374, 32'sd-0.01095745321142196, 32'sd0.07256330148062644, 32'sd0.044161744812563214, 32'sd-0.03269485966153907, 32'sd-0.0771944682476363, 32'sd-0.050025658984686215, 32'sd-0.012549320053493289, 32'sd-0.09433911821607695, 32'sd0.011893225099933815, 32'sd0.028957210661799942, 32'sd-0.014761708038975101, 32'sd-0.01915375462925863, 32'sd0.05676475157721873, 32'sd-0.0026644364563714984, 32'sd0.06752824438277856, 32'sd0.035114204016686794, 32'sd0.009990627048355662, 32'sd0.08079238884740386, 32'sd0.1618513355615694, 32'sd0.06884880340162888, 32'sd0.14112772835297516, 32'sd0.07799292520085632, 32'sd0.11703749680138845, 32'sd0.11226277938941967, 32'sd0.13183230542509275, 32'sd0.12296078425415888, 32'sd0.02499965537709576, 32'sd0.08778382124463363, 32'sd0.07033184311110478, 32'sd-0.010911874750667704, 32'sd0.021753080363438097, 32'sd-0.001620775628086252, 32'sd-0.030309837060406127, 32'sd0.011906835372329084, 32'sd-0.06379568053477093, 32'sd-0.0907374871760275, 32'sd0.05983440182813504, 32'sd9.923901897415181e-122, 32'sd-0.06924325166296177, 32'sd-0.1253002729210682, 32'sd0.0893164219041862, 32'sd0.02984592101627537, 32'sd-0.04575003748961813, 32'sd-0.01807752911041353, 32'sd0.033186302398288806, 32'sd0.17240040493872644, 32'sd0.21140283256303122, 32'sd0.19060448666012023, 32'sd0.1539446187200657, 32'sd0.24710266634409575, 32'sd0.21610631756303594, 32'sd0.00269197001798018, 32'sd0.04363408309501657, 32'sd0.0036687094462824303, 32'sd0.12839048338648726, 32'sd0.02483326506197388, 32'sd-0.018917166153966228, 32'sd0.04221368359943615, 32'sd0.05567118491195578, 32'sd0.0023220357911652354, 32'sd-0.0074923313328375965, 32'sd0.04256314701671324, 32'sd-0.003666678943003739, 32'sd0.001191388802880843, 32'sd0.06079754647487054, 32'sd0.08650615282337966, 32'sd0.02598852469792147, 32'sd0.02048819331835907, 32'sd-0.020637844845126, 32'sd0.07295611209267167, 32'sd-0.005726538046523171, 32'sd-0.06825913515578504, 32'sd0.006739929540817819, 32'sd0.10833612799847099, 32'sd0.09614609020031956, 32'sd0.03136162913278823, 32'sd0.12158813040234633, 32'sd0.14232214508085786, 32'sd0.12412496849112993, 32'sd0.13926880845794956, 32'sd0.007941457305819338, 32'sd-0.11638074978002072, 32'sd0.04589836915507611, 32'sd-0.07473482123636563, 32'sd-0.09679877505731643, 32'sd0.03325937124517259, 32'sd-0.08010857110679921, 32'sd0.039647374480889216, 32'sd0.03644807607088621, 32'sd-0.11208499678624813, 32'sd0.04634382389575673, 32'sd0.027055613668193527, 32'sd0.10523570292712929, 32'sd0.042942039620345665, 32'sd0.058590188576105214, 32'sd-0.07856842084862292, 32'sd-0.006062829727156729, 32'sd0.013698958181824088, 32'sd-0.036541247825315946, 32'sd0.06429851557124372, 32'sd-0.004332504742452172, 32'sd-0.05167733489681488, 32'sd-0.051806485663407904, 32'sd-0.01986890566933877, 32'sd0.05084049736053264, 32'sd0.10103565788317921, 32'sd0.1220718211007543, 32'sd0.05902888196938855, 32'sd0.1134735328707696, 32'sd0.03626319891896055, 32'sd0.034676126809522534, 32'sd-0.04595240733034551, 32'sd-0.06531146343120085, 32'sd-0.012971969763978805, 32'sd-0.09141652991184392, 32'sd-0.017519924467168227, 32'sd0.022716580583211354, 32'sd0.0035291670648979977, 32'sd0.1233893889386805, 32'sd0.08631129610226998, 32'sd0.05223912684610407, 32'sd4.195709368891713e-123, 32'sd0.09898147330242424, 32'sd0.06826149866409555, 32'sd-0.09220471039062528, 32'sd-0.11063923955371101, 32'sd-0.052128263015304384, 32'sd0.07560215117341322, 32'sd0.02578128668620032, 32'sd0.07483054946441581, 32'sd0.08032192936616117, 32'sd0.08142267754890162, 32'sd0.13121641847640478, 32'sd0.03175058539609598, 32'sd-0.019174740639510055, 32'sd0.03356060260239129, 32'sd0.12490250557696844, 32'sd0.12309308968799822, 32'sd0.11013217419230241, 32'sd0.030954082584775725, 32'sd-0.05676421982898002, 32'sd-0.033083802162024875, 32'sd-0.08189704633033938, 32'sd-0.05210434364096712, 32'sd0.012650526060958654, 32'sd0.056287763175817886, 32'sd-0.04937986267881704, 32'sd0.12162373944395406, 32'sd-2.1677717823005273e-124, 32'sd-2.5834766824538363e-116, 32'sd8.01379372003124e-128, 32'sd0.03264416253122671, 32'sd-0.02179027432084607, 32'sd-0.09409041527412977, 32'sd0.00655232345374614, 32'sd0.003351130790521348, 32'sd0.15952471774461136, 32'sd0.0812745744035781, 32'sd0.06132598465687932, 32'sd0.08052235750581933, 32'sd0.06510699357164375, 32'sd0.11932204200708706, 32'sd0.08333841467841425, 32'sd0.12490442992415987, 32'sd0.030932709111333008, 32'sd-0.02707751343961494, 32'sd0.10466295465927077, 32'sd0.03913400145214315, 32'sd-0.018757847579803578, 32'sd0.013027515318711769, 32'sd0.015133857296773821, 32'sd0.024686418642274045, 32'sd0.012165352225826532, 32'sd0.1335111594724522, 32'sd0.05680768146883099, 32'sd0.04753764449945139, 32'sd-1.369583127730918e-123, 32'sd-3.2041550090530126e-119, 32'sd2.966353725292154e-120, 32'sd0.09745453921839295, 32'sd0.03266057549822164, 32'sd-0.0507073306092849, 32'sd0.010957124085045681, 32'sd-0.028420768313205353, 32'sd0.06595238076110176, 32'sd0.12111038833318816, 32'sd0.12720929299554481, 32'sd-0.037318239443632696, 32'sd-0.11256104071517896, 32'sd0.10824606597288186, 32'sd0.07408374523219546, 32'sd0.07545543688812399, 32'sd0.009135711106703144, 32'sd0.02207625998190008, 32'sd-0.23069799991154208, 32'sd-0.15717146598778495, 32'sd-0.02150640261268957, 32'sd-0.012640056266388068, 32'sd-0.017095331840637284, 32'sd-0.023226466281486453, 32'sd0.05068758700582037, 32'sd0.0712780524058916, 32'sd0.09307326411109558, 32'sd-0.054349363594221975, 32'sd-4.092874627353764e-123, 32'sd-1.4699812775185212e-123, 32'sd-4.817499531251764e-115, 32'sd5.5029488209948755e-126, 32'sd0.0697652934101861, 32'sd0.054420429112099086, 32'sd0.0320823525594039, 32'sd0.0638452291363018, 32'sd-0.04848148193048384, 32'sd0.009060576120246324, 32'sd0.004331903636099017, 32'sd0.08745849420320163, 32'sd-0.02186993084914157, 32'sd-0.020649254404571594, 32'sd-0.08392076824111017, 32'sd0.009114595511809305, 32'sd0.06919049505742318, 32'sd0.03631099275393209, 32'sd0.0628165994851485, 32'sd-0.07805443298670327, 32'sd-0.023196790377120788, 32'sd0.014647557215281402, 32'sd-0.04404226047366468, 32'sd-0.006822829897473537, 32'sd-0.03271097165666614, 32'sd0.016318276876741578, 32'sd0.03506026295010212, 32'sd3.904908911162299e-124, 32'sd-2.0753304371469924e-123, 32'sd1.6869600176364911e-125, 32'sd4.805845691596117e-124, 32'sd-1.0390508119430538e-115, 32'sd-6.422447252341212e-121, 32'sd0.017284528759755925, 32'sd0.08715680956231481, 32'sd0.01924317740681617, 32'sd0.06622797378691526, 32'sd0.056373625563068505, 32'sd0.02124813531752506, 32'sd0.06721522152830892, 32'sd0.007076086386985924, 32'sd0.018667675593581352, 32'sd0.06124502143042143, 32'sd0.049785056693059805, 32'sd-0.01269373623283151, 32'sd-0.02286359590933297, 32'sd0.041421984595008766, 32'sd8.716708963330786e-05, 32'sd-0.005473259734719321, 32'sd0.041967316102494275, 32'sd0.010944264080292167, 32'sd0.09067202141126282, 32'sd0.029898268389126636, 32'sd1.6941394765240515e-127, 32'sd1.6085908525516036e-115, 32'sd1.62776324575974e-115, 32'sd4.098567120366012e-122},
        '{32'sd3.2387937067146247e-121, 32'sd3.4561045333127844e-120, 32'sd-1.535528511504571e-123, 32'sd1.8768730380130967e-127, 32'sd-4.607049987958228e-127, 32'sd-9.295357312339751e-127, 32'sd4.32112116305068e-125, 32'sd1.0537072971521046e-122, 32'sd2.4472674666012083e-115, 32'sd-5.9134585872195355e-120, 32'sd3.8652466537485427e-115, 32'sd-6.65768077087128e-126, 32'sd0.08295827309054424, 32'sd0.07642488844763606, 32'sd0.16575432315644908, 32'sd0.1093635155209059, 32'sd-8.53272109886607e-125, 32'sd-3.1318031836394375e-120, 32'sd9.44918615174367e-128, 32'sd2.205939283984983e-121, 32'sd1.7715478747165815e-124, 32'sd1.0090066440937667e-121, 32'sd3.506165353186944e-114, 32'sd-4.121631401614865e-127, 32'sd-1.2806185000887293e-122, 32'sd3.8802546464385e-124, 32'sd-1.7203785477440932e-122, 32'sd1.652466409148875e-126, 32'sd3.849124198920079e-129, 32'sd-8.130468971863467e-124, 32'sd3.406177163057053e-119, 32'sd5.706395919132159e-120, 32'sd-0.00015999414734407366, 32'sd0.045697776886362465, 32'sd-0.005969016981987799, 32'sd-0.08180612711206499, 32'sd0.021539739322777942, 32'sd-0.02662291490888234, 32'sd0.12925997712191473, 32'sd0.05611232653836552, 32'sd0.0884763983971158, 32'sd0.07003979254601281, 32'sd-0.02113870921543306, 32'sd0.12682214978150927, 32'sd0.0834852336867526, 32'sd0.08950985223018447, 32'sd0.1311032916782217, 32'sd0.058549520764114585, 32'sd0.011466464293237987, 32'sd0.06365387816180919, 32'sd0.06654811588937615, 32'sd0.07533702023944094, 32'sd6.3672667169266585e-124, 32'sd6.390374756784941e-122, 32'sd-3.305525674736148e-122, 32'sd-9.961687823345775e-121, 32'sd-4.150849006071284e-121, 32'sd-2.519863383105126e-125, 32'sd0.13214223712192902, 32'sd0.08342612632762642, 32'sd0.08477677132707047, 32'sd-0.07067347467122341, 32'sd0.04535803912320376, 32'sd-0.008917177689167426, 32'sd-0.035210809546107585, 32'sd0.1342072808974388, 32'sd-0.0023378142620811347, 32'sd0.11902256890455558, 32'sd-0.05204909463993919, 32'sd-0.14436002671763085, 32'sd0.007561724611824228, 32'sd0.11326039185302915, 32'sd-0.042796728033455154, 32'sd0.03454813979648516, 32'sd0.018590511719362723, 32'sd0.002337894918437741, 32'sd-0.008973007420418589, 32'sd-0.016881118368940507, 32'sd0.08552297190491141, 32'sd0.05551907997327253, 32'sd0.02181216225764755, 32'sd0.12438821552244576, 32'sd1.0557652896296646e-115, 32'sd-7.307568258381333e-128, 32'sd5.790897831310095e-126, 32'sd7.427956095852599e-115, 32'sd-0.026816393460566326, 32'sd0.08089366994911484, 32'sd-0.02872284433714369, 32'sd0.005216255572811046, 32'sd0.01735060920236402, 32'sd-0.031870337760813765, 32'sd0.06374894456507808, 32'sd0.13480987887791213, 32'sd-0.06601068543626287, 32'sd0.008517402255766318, 32'sd-0.10516533183270767, 32'sd-0.030866107236875436, 32'sd-0.046881811093205925, 32'sd0.035207874673265166, 32'sd0.02931906333509085, 32'sd0.11696213496072348, 32'sd0.07025973132080834, 32'sd0.011701976576327922, 32'sd0.05078404205024496, 32'sd-0.012350159895163615, 32'sd0.09058558180235537, 32'sd0.020613902371137433, 32'sd-0.004360110237968532, 32'sd0.036088605019164624, 32'sd0.05815736555877196, 32'sd1.0552353061543882e-121, 32'sd-6.743015773261758e-119, 32'sd0.06084429723227113, 32'sd0.04165968399064299, 32'sd-0.04372367053272109, 32'sd-0.007761195105887132, 32'sd0.014557115756591367, 32'sd-0.03481578006745966, 32'sd0.0398846504819046, 32'sd0.09038196521861232, 32'sd0.09618073313592053, 32'sd0.06008178323032172, 32'sd0.007048854188691697, 32'sd-0.03698028162993047, 32'sd-0.1322059110646733, 32'sd-0.17975421672441755, 32'sd-0.051593693216631785, 32'sd-0.1437973036310106, 32'sd0.05356696669089951, 32'sd0.03348947229769325, 32'sd0.01619330727258211, 32'sd0.01753698236851188, 32'sd-0.07173118323819636, 32'sd-0.07164656775014182, 32'sd0.014126655564434216, 32'sd-0.02605045949120656, 32'sd-0.08055186458580824, 32'sd-0.06953223395751419, 32'sd0.07184356126349056, 32'sd-3.9577677198069465e-117, 32'sd0.07854345446222893, 32'sd0.10963169170291141, 32'sd0.03036305014309486, 32'sd0.01890022891259845, 32'sd-0.08452135390940832, 32'sd-0.04406028136447945, 32'sd0.11904786820885815, 32'sd0.0777034786213171, 32'sd0.05746907808893039, 32'sd0.06550879410427618, 32'sd0.011524581183388564, 32'sd-0.10399212605914909, 32'sd0.012431857121068212, 32'sd-0.12285242629806369, 32'sd-0.030281244705516693, 32'sd-0.1425560719418459, 32'sd-0.11054018300489067, 32'sd-0.06377233971313927, 32'sd-0.03699636207298875, 32'sd-0.0792360490093042, 32'sd-0.21593772694574281, 32'sd-0.12083533966024455, 32'sd-0.032393138842884237, 32'sd-0.042778957252168535, 32'sd-0.04784152522872672, 32'sd-0.037372368838912366, 32'sd0.014332802378059088, 32'sd-5.824775165936797e-124, 32'sd0.018235824620849907, 32'sd0.05804092803154208, 32'sd-0.07346713711996934, 32'sd-0.002376908332843994, 32'sd0.0065500534022088774, 32'sd0.008188757314196571, 32'sd0.009404378780092268, 32'sd-0.04268210813728456, 32'sd0.07788321427360358, 32'sd-0.05344781612849911, 32'sd-0.046894231947965034, 32'sd-0.014802555027196313, 32'sd0.04393877102530263, 32'sd0.0766874292200218, 32'sd0.0212572417922864, 32'sd0.03079904700974558, 32'sd0.10220783231390741, 32'sd0.05465047329322517, 32'sd0.03099775947946398, 32'sd-0.03732532109429501, 32'sd-0.06470039302290904, 32'sd-0.03027943024159385, 32'sd-0.16483133097232225, 32'sd-0.054785718057284175, 32'sd-0.09042025607368549, 32'sd-0.031436279300953086, 32'sd-0.005135640286460033, 32'sd0.08287578287549971, 32'sd0.060588554633612846, 32'sd0.025016821998357367, 32'sd0.07116986374171674, 32'sd0.06069171017562243, 32'sd0.09425136680741521, 32'sd0.007370736027675033, 32'sd-0.0625795632497322, 32'sd-0.0013358675091001385, 32'sd-0.015464155481025789, 32'sd-0.16381519033566516, 32'sd-0.08433015081190791, 32'sd0.04153747249679178, 32'sd0.15579342781818112, 32'sd-0.010103669190141693, 32'sd-0.12048665621971719, 32'sd-0.14534953590082259, 32'sd0.05114078992922362, 32'sd-0.07474826738573499, 32'sd-0.0278923214077536, 32'sd-0.06073696706025943, 32'sd-0.13560484304624054, 32'sd-0.08958572556490528, 32'sd0.056567025100901, 32'sd0.02113436682619365, 32'sd-0.05963439220574884, 32'sd0.05807609187977645, 32'sd-0.0494897563067802, 32'sd0.04522320363391745, 32'sd0.04446628703502226, 32'sd0.05579222423575211, 32'sd0.01895558888707572, 32'sd-0.07705628632398677, 32'sd0.0445348913741688, 32'sd-0.018999314935418714, 32'sd0.03995566623266353, 32'sd-0.004505013028967263, 32'sd-0.09617553761470897, 32'sd-0.014087525085359293, 32'sd0.03408151664570855, 32'sd0.04018832269923831, 32'sd0.013471913507703425, 32'sd0.11738800266133842, 32'sd-0.14761214599079495, 32'sd-0.10656849486463785, 32'sd-0.14740610779393246, 32'sd0.01217553231639831, 32'sd-0.04704276341157205, 32'sd-0.1136317949109099, 32'sd-0.1675758743327339, 32'sd-0.1229087143976766, 32'sd0.010566708515090733, 32'sd0.030643034496333814, 32'sd0.01199852030641297, 32'sd0.023162668035555792, 32'sd0.060122211173506294, 32'sd0.11532980840101893, 32'sd0.1461048414086495, 32'sd-0.037366034710961886, 32'sd0.050419023388264386, 32'sd-0.0030396761607045636, 32'sd0.18703269645802081, 32'sd0.14830242989841055, 32'sd0.0356057829036182, 32'sd-0.03102428236154685, 32'sd-0.05284549601378347, 32'sd0.07116208098423218, 32'sd0.11315256243435379, 32'sd0.16385356584409327, 32'sd0.08898847962373804, 32'sd0.1286163983255536, 32'sd-0.016997254384977404, 32'sd-0.20075297544335502, 32'sd-0.13627500031964124, 32'sd0.028425026913010566, 32'sd-0.07420372757123912, 32'sd-0.11393125815070361, 32'sd-0.10984005505544706, 32'sd-0.058525981432247146, 32'sd-0.002850539884458296, 32'sd0.038021297751130105, 32'sd-0.04253078157895329, 32'sd-0.026064597700343483, 32'sd-0.003270347400348508, 32'sd0.03514056083033896, 32'sd0.07171772183668507, 32'sd0.06749664690514055, 32'sd0.025425939519984682, 32'sd0.0032257721801464793, 32'sd0.15293869234249252, 32'sd0.096300414510776, 32'sd0.04081820421313577, 32'sd-0.027968068907342367, 32'sd0.028694790283721208, 32'sd-0.10277878043740091, 32'sd0.08760898073318069, 32'sd0.10915043783543006, 32'sd0.13876257656815277, 32'sd-0.0003757128198201673, 32'sd-0.039574442984694626, 32'sd-0.018993210304683154, 32'sd-0.1535562740545161, 32'sd-0.024879760121897673, 32'sd0.1091110768298915, 32'sd0.03618467333678904, 32'sd-0.0952654873556125, 32'sd-0.15369053434836807, 32'sd-0.025737073613057267, 32'sd0.1538860163174365, 32'sd0.024013247813197754, 32'sd-0.02992593842036784, 32'sd0.024512275199592325, 32'sd0.005499379377866346, 32'sd-0.055597241182871245, 32'sd0.024217597915321333, 32'sd0.09358104697705101, 32'sd0.0035904785828797174, 32'sd-0.0330089950850478, 32'sd-0.020458145202889032, 32'sd0.14591047667173096, 32'sd-0.014253533315924903, 32'sd-0.11096105730891749, 32'sd-0.10913416384727975, 32'sd-0.029818504685253846, 32'sd0.06761701296634133, 32'sd-0.04047935736493026, 32'sd0.0700220940669663, 32'sd0.07362381697329466, 32'sd0.09220834461641612, 32'sd0.0039575470038633095, 32'sd0.05793612735639098, 32'sd0.12224376370480548, 32'sd0.10930285744754745, 32'sd-0.1147385304803071, 32'sd-0.08827230147491472, 32'sd-0.0018353087156460792, 32'sd-0.09234027951323774, 32'sd-0.07408088944247371, 32'sd-0.07453414863534776, 32'sd-0.05133105785669151, 32'sd0.05118967906334072, 32'sd-0.08119967818227018, 32'sd-0.01620916398613167, 32'sd-0.04109772891518559, 32'sd-0.03326581970120236, 32'sd-0.002167734621160846, 32'sd-0.12539544044020995, 32'sd0.039732104284108845, 32'sd-0.0014325013874874556, 32'sd-0.1822692802100049, 32'sd-0.028251675537857592, 32'sd0.02339296293902422, 32'sd-0.002731111898663249, 32'sd-0.06776051753896907, 32'sd0.016864345217522322, 32'sd0.11986858775450782, 32'sd0.15183986545295727, 32'sd-0.046050370121611686, 32'sd0.04090367051036698, 32'sd0.05057677982744276, 32'sd-0.01483161804068272, 32'sd0.07936758928677982, 32'sd-0.09992618166436427, 32'sd-0.044781861678571046, 32'sd-0.055839605104827474, 32'sd0.10479652745675071, 32'sd0.044250120950441826, 32'sd0.0024708790256534703, 32'sd0.00640375649146254, 32'sd-0.013414842866560986, 32'sd0.031565058526501245, 32'sd-0.11149450706072711, 32'sd-0.010084981764577252, 32'sd-0.02375937054778394, 32'sd-0.030083462047230898, 32'sd-0.060878423264245744, 32'sd-0.08963588407198604, 32'sd-0.044549643627887686, 32'sd0.00539458845719606, 32'sd0.0989385820930262, 32'sd0.09960315496865967, 32'sd0.18938844306938654, 32'sd0.15388212859286815, 32'sd0.03875052853801405, 32'sd0.0759219664253658, 32'sd-0.07064988613431152, 32'sd-0.010862598213666615, 32'sd0.0433862862963524, 32'sd0.06561596726989573, 32'sd0.034489093831171665, 32'sd0.015342547557623902, 32'sd-0.009033212408527365, 32'sd0.17159484681803097, 32'sd0.0902953004988042, 32'sd-0.05729513338224146, 32'sd-0.10259474630986398, 32'sd0.0614764941051703, 32'sd0.0036824534644719267, 32'sd-0.09444910247782941, 32'sd0.04103944623177603, 32'sd0.003566282340318299, 32'sd-0.014464404224760495, 32'sd0.011350885553691981, 32'sd0.07533728106177383, 32'sd0.03258135053680548, 32'sd0.02120563863000627, 32'sd0.14351283462002212, 32'sd0.09627364831917676, 32'sd0.09051713298757683, 32'sd0.04080485736586885, 32'sd0.061141621571545283, 32'sd0.08108740639364768, 32'sd0.1212311735768356, 32'sd0.03564266044979866, 32'sd0.15179968656786974, 32'sd0.15113779249276835, 32'sd0.10323096773823323, 32'sd0.10327988947300583, 32'sd0.10531461972425457, 32'sd0.043036895426582934, 32'sd-0.031789827199263786, 32'sd-0.0041812183566052276, 32'sd-0.05472005072868138, 32'sd0.15545357258488682, 32'sd-0.021886901206426335, 32'sd0.024770656589103695, 32'sd0.028314374380075783, 32'sd0.01683113991698816, 32'sd-0.003294121265056993, 32'sd-0.06266428904466216, 32'sd-0.008902076660240097, 32'sd-0.05416731232434308, 32'sd0.055210158289572805, 32'sd0.10203706315117704, 32'sd0.13326195783996822, 32'sd0.17629751743600275, 32'sd0.050084686510375356, 32'sd0.0408898084385801, 32'sd-0.008290172897264502, 32'sd0.16172355783113163, 32'sd-0.042160927912479544, 32'sd0.1102777030254716, 32'sd0.1666588195379464, 32'sd0.10695494695997428, 32'sd0.05340852347671347, 32'sd0.11927075302495908, 32'sd-0.027042413379625357, 32'sd-0.009906656720732206, 32'sd0.11310000923645182, 32'sd0.038353474591491174, 32'sd0.08519998156704232, 32'sd0.0025440782947545207, 32'sd0.05956065138656451, 32'sd0.02552777251866767, 32'sd0.018217120347925053, 32'sd0.0023452665329144334, 32'sd0.03575401242078343, 32'sd-0.05625249844860549, 32'sd0.030563390163381218, 32'sd0.05795962544610337, 32'sd0.13916489816530023, 32'sd0.0025046966602621915, 32'sd0.041124295731225245, 32'sd0.20134748107296532, 32'sd0.012177879657108495, 32'sd0.031854111985675934, 32'sd0.0775498977750722, 32'sd0.0613269420671536, 32'sd-0.049535839099915865, 32'sd0.03880231142027021, 32'sd0.13446807536618946, 32'sd-0.00930764612051732, 32'sd0.035752437246816746, 32'sd0.1405077540091727, 32'sd0.038760227964198965, 32'sd0.08305415449613919, 32'sd-0.026330554232527992, 32'sd0.0014931693371653832, 32'sd-0.09617448285115236, 32'sd0.02162522092849276, 32'sd-1.0034801647336387e-126, 32'sd0.023903694344562836, 32'sd-0.10421713917269182, 32'sd-0.09529238127529499, 32'sd0.06439485399680596, 32'sd0.05617859979814287, 32'sd-0.05025994211904137, 32'sd-0.06221792380145921, 32'sd-0.04507712654509468, 32'sd0.025184545483105208, 32'sd0.10927856907354078, 32'sd0.06312853538812396, 32'sd-0.058393173729564825, 32'sd0.02201096936610788, 32'sd0.07695338791761115, 32'sd0.0640244522741717, 32'sd-0.06111676104688507, 32'sd-0.06488915160606247, 32'sd-0.007747205016488857, 32'sd0.1146987046956126, 32'sd0.11669893281511204, 32'sd0.059746368247117126, 32'sd0.0173669159953608, 32'sd0.11819303519989492, 32'sd0.04653186947555076, 32'sd0.09118825902882524, 32'sd-0.07482477878544175, 32'sd-0.024918427454111748, 32'sd-0.0344069416514604, 32'sd-0.03620970319359505, 32'sd-0.07102353823396661, 32'sd-0.028025764673743007, 32'sd0.03332577210918367, 32'sd-0.08246947331176244, 32'sd-0.12627127554987663, 32'sd-0.1006859022237935, 32'sd-0.045371346373867825, 32'sd0.03334333683827131, 32'sd0.0009083922690699811, 32'sd-0.11732730476368645, 32'sd-0.07990600601350957, 32'sd0.009583384160163149, 32'sd-0.012601156250447438, 32'sd-0.14397343789516961, 32'sd-0.23966165351781446, 32'sd-0.09689280312196993, 32'sd-0.05336376876621756, 32'sd0.0032014442056809513, 32'sd-0.10392084823640893, 32'sd-0.0710144492176033, 32'sd-0.005146777852489199, 32'sd0.04669230679517875, 32'sd0.03546564780930457, 32'sd-0.006324405837563043, 32'sd-0.00256997605765055, 32'sd-0.03088597837426139, 32'sd0.013096173674650107, 32'sd0.04552413367848948, 32'sd0.013694393386972814, 32'sd-0.07595252138036546, 32'sd-0.037014359930531884, 32'sd-0.0670187540375545, 32'sd-0.0570664579408895, 32'sd-0.07970739958363718, 32'sd-0.12879231689088208, 32'sd-0.07901082250049891, 32'sd-0.10151007756269768, 32'sd-0.009935643680951177, 32'sd-0.12762408122845395, 32'sd-0.08368319567645947, 32'sd0.024126718144266635, 32'sd-0.0692206360335399, 32'sd-0.1009016004096539, 32'sd-0.03470875272587165, 32'sd-0.1533296836932818, 32'sd-0.07618838778823776, 32'sd-0.13927669155323694, 32'sd-0.1398427852331746, 32'sd-0.07721832245497795, 32'sd-0.058551819873662675, 32'sd0.004731389019688612, 32'sd-0.04090829840885101, 32'sd-0.02559409857564476, 32'sd0.06375965265286995, 32'sd-2.0368793071592288e-120, 32'sd0.0005248592180918315, 32'sd-0.01803801321557583, 32'sd-0.05009653834881748, 32'sd-0.022367409919152273, 32'sd-0.008083189667424943, 32'sd-0.16074220162980643, 32'sd-0.14300497531042222, 32'sd-0.1678219514236713, 32'sd-0.16708778238068753, 32'sd-0.14858023032115622, 32'sd-0.07622219012470717, 32'sd0.045770255420473666, 32'sd-0.14563793609747724, 32'sd0.013304304507229447, 32'sd-0.1295872697573821, 32'sd-0.012889798023968098, 32'sd-0.14098932055569308, 32'sd-0.20913757546511363, 32'sd-0.1656106637433292, 32'sd-0.11554310386773867, 32'sd-0.14322057592072, 32'sd-0.040937061704061396, 32'sd-0.0904578321505804, 32'sd0.052552774293297834, 32'sd0.01815863734826584, 32'sd-0.0829944490810265, 32'sd0.04249701567555684, 32'sd0.028441048027694118, 32'sd-0.040178954884806405, 32'sd-0.10324521874936246, 32'sd-0.05192208424239561, 32'sd0.022036058804456415, 32'sd-0.04637797845137946, 32'sd-0.07119345997918983, 32'sd-0.11294149333214035, 32'sd-0.10576173839100632, 32'sd-0.1382118629531187, 32'sd-0.04403496297092157, 32'sd-0.09871413308962824, 32'sd-0.03662561895375518, 32'sd-0.19774033490451687, 32'sd-0.2144739110297467, 32'sd-0.1214557717689126, 32'sd-0.06783343400734769, 32'sd-0.13408928555867844, 32'sd-0.2195320434237487, 32'sd-0.18264585929272364, 32'sd-0.1840399410946135, 32'sd-0.11941313667663273, 32'sd-0.062176648144507136, 32'sd-0.11251418517430563, 32'sd-0.005974141504986117, 32'sd-0.026030239553040395, 32'sd-0.037144661893656054, 32'sd-0.015745711923783805, 32'sd-0.05260656448812678, 32'sd0.038346636861898584, 32'sd-0.0770730248795699, 32'sd0.06186028215976863, 32'sd-0.04299117784772028, 32'sd0.004265606774848247, 32'sd-0.0009317783890406218, 32'sd0.00785460849460194, 32'sd-0.06363897528558284, 32'sd-0.09691322502439537, 32'sd-0.00800771467443671, 32'sd-0.15664322647384196, 32'sd-0.09558248999207826, 32'sd-0.07341779539278613, 32'sd-0.10082648061205145, 32'sd-0.11816811980029478, 32'sd-0.049934523862306644, 32'sd-0.08276755756596614, 32'sd-0.12082490379470236, 32'sd-0.09464467997131144, 32'sd-0.02619339334441269, 32'sd-0.19140049260816208, 32'sd-0.0054440357339661325, 32'sd-0.028774174129297826, 32'sd-0.032959467410877276, 32'sd-0.051762858000999966, 32'sd-0.0026714926134055587, 32'sd0.013544122599806564, 32'sd-4.932031603955018e-115, 32'sd0.06529180589450684, 32'sd-0.05350359386086511, 32'sd-0.05532107179905098, 32'sd-0.0637463568157838, 32'sd-0.1613933205712976, 32'sd0.07052225596534661, 32'sd-0.03188693469190532, 32'sd-0.03178102039762289, 32'sd0.009786527285155644, 32'sd-0.051823932124013275, 32'sd-0.1963164167779365, 32'sd-0.08261658974936645, 32'sd-0.04157776269238646, 32'sd0.03717329284809662, 32'sd-0.08447894067448679, 32'sd-0.11400389680895459, 32'sd0.012444884793009705, 32'sd-0.04257081338796093, 32'sd-0.051793057803961075, 32'sd-0.1340264479223927, 32'sd-0.20150338669510914, 32'sd-0.06531723750693345, 32'sd0.06253915477072697, 32'sd0.05082931694106608, 32'sd-0.0026310469648961484, 32'sd-0.0702998487855534, 32'sd5.110634372370736e-123, 32'sd1.9212948990145694e-120, 32'sd-3.89146667846938e-123, 32'sd0.08238933339606717, 32'sd0.052470719399223174, 32'sd-0.10373900344741474, 32'sd-0.018518379118121986, 32'sd-0.0862509155534167, 32'sd0.03587026193992134, 32'sd0.0973602479659628, 32'sd-0.011672010886867683, 32'sd-0.07780923610092023, 32'sd-0.08198734443888585, 32'sd-0.015802220595789052, 32'sd-0.06578482669443501, 32'sd-0.014517781345495398, 32'sd0.060899099607844155, 32'sd-0.04847191617563918, 32'sd0.05444335995154497, 32'sd-0.0234843255501218, 32'sd0.04856246229652797, 32'sd0.06391606088002101, 32'sd-0.056981980937668306, 32'sd-0.10329841482450562, 32'sd0.07058054790489471, 32'sd-0.01365974636646109, 32'sd-0.10699549782220227, 32'sd0.09030031202511624, 32'sd1.6889818218479682e-121, 32'sd3.5589899815269783e-116, 32'sd-4.207251975646901e-125, 32'sd0.0288596630449165, 32'sd-0.007466345915915001, 32'sd-0.0031122578307117947, 32'sd-0.062430260906594655, 32'sd-0.011225049891540731, 32'sd0.06407498163224443, 32'sd0.04566985279373566, 32'sd-0.07131242541586681, 32'sd-0.07544622915507182, 32'sd-0.03673205323361506, 32'sd0.01235586664110754, 32'sd0.041536472468048403, 32'sd0.08745664885871357, 32'sd0.042817232646166915, 32'sd0.16146035050630198, 32'sd0.14349544833265326, 32'sd0.024293634363716777, 32'sd-0.04353519450929917, 32'sd0.08599871974576993, 32'sd0.05878207308833762, 32'sd-0.09434666459238412, 32'sd-0.1089695109216649, 32'sd-0.05040753803487946, 32'sd0.08066914738215525, 32'sd0.10344166901323498, 32'sd3.381964903830092e-120, 32'sd-8.583703320374748e-118, 32'sd1.5697670154661164e-124, 32'sd-6.909119638479803e-117, 32'sd0.11164446925139589, 32'sd0.06339178042527685, 32'sd-0.06853409497860463, 32'sd0.05201016972462453, 32'sd0.09309190818049151, 32'sd0.004403733207541575, 32'sd0.047080490596453646, 32'sd0.04437025917152987, 32'sd0.003974014436208555, 32'sd-0.005858260045681144, 32'sd0.0745980151087248, 32'sd0.1693939441862819, 32'sd-0.021802347674961652, 32'sd0.06526898967158345, 32'sd-0.05247725576934026, 32'sd-0.019396614337821427, 32'sd0.010411221452570342, 32'sd0.02183875685622898, 32'sd-0.01580797538125382, 32'sd0.03295735683948413, 32'sd0.05533671625048036, 32'sd0.028477969084221115, 32'sd0.07613928582528716, 32'sd-1.837989928503083e-121, 32'sd8.637972669257134e-117, 32'sd1.1044692564208074e-123, 32'sd5.405974419104024e-118, 32'sd2.3771029418960943e-128, 32'sd-4.860497623260267e-128, 32'sd0.13097656236913768, 32'sd0.06991897331653046, 32'sd0.08648821122983807, 32'sd0.04093668121443401, 32'sd0.01820884884349691, 32'sd0.05406176682399717, 32'sd0.08364548798343235, 32'sd0.08614301416350724, 32'sd-0.034078914541305544, 32'sd0.11609181989331252, 32'sd-0.025058772418387165, 32'sd0.1209067100393074, 32'sd0.005036837393679498, 32'sd0.1127320772243168, 32'sd0.03534291420077989, 32'sd0.012171776891900432, 32'sd-0.03653578043306507, 32'sd0.05016569400375195, 32'sd-0.021426294073375568, 32'sd0.17288833350377852, 32'sd-7.380840950409551e-117, 32'sd-1.3214998176936565e-118, 32'sd9.865092993595429e-121, 32'sd2.1172757554004627e-117},
        '{32'sd3.6857838000572277e-118, 32'sd5.985341660737281e-124, 32'sd-9.955686929891293e-122, 32'sd-1.3663113409326587e-123, 32'sd9.785644399972107e-125, 32'sd-5.251377377130258e-116, 32'sd7.308436105904065e-119, 32'sd7.792245344726268e-127, 32'sd-1.549819152644037e-123, 32'sd1.338186926638624e-128, 32'sd7.912123272560294e-118, 32'sd-3.049322958661182e-116, 32'sd-0.024280955401150817, 32'sd0.023549513000194974, 32'sd0.12274499966603657, 32'sd0.01433549620715614, 32'sd-1.73722118645691e-125, 32'sd1.8434085522944235e-116, 32'sd3.827286426702999e-117, 32'sd-2.579634216916931e-126, 32'sd1.0345543378916173e-121, 32'sd1.814812527512018e-116, 32'sd-4.379662610257958e-123, 32'sd3.496302402135884e-116, 32'sd9.382811246188365e-116, 32'sd-1.2091249390239629e-122, 32'sd1.0770809735357501e-122, 32'sd1.4058508671473327e-123, 32'sd1.3190117443729077e-122, 32'sd-7.478627149111245e-126, 32'sd-2.290449650080423e-121, 32'sd2.8166894104297282e-123, 32'sd0.04701843622713209, 32'sd-0.09182447428333049, 32'sd-0.009667439968513797, 32'sd-0.02303397960863846, 32'sd-0.024663797309173882, 32'sd0.013605604949178467, 32'sd-0.004588464381175541, 32'sd0.03753523337802995, 32'sd-0.00856769012840482, 32'sd-0.04481475479166874, 32'sd0.08434736526402793, 32'sd0.04907165588951692, 32'sd0.05821930260809442, 32'sd0.005804712725991096, 32'sd-0.07606562835736116, 32'sd0.05803158150630028, 32'sd-0.013073112946150687, 32'sd0.14656975465762787, 32'sd0.1023187605594387, 32'sd0.052659532599653204, 32'sd1.3414547670109462e-122, 32'sd-1.228733857818258e-121, 32'sd9.398328165637459e-116, 32'sd-1.8115791085572855e-124, 32'sd-1.5424370958397132e-123, 32'sd1.1719513203946817e-125, 32'sd0.07489630428819966, 32'sd0.05277975051140797, 32'sd-0.0074520550393085555, 32'sd-0.01548492127506595, 32'sd-0.0663905429060089, 32'sd-0.10650817113357407, 32'sd0.02363832034882049, 32'sd0.0867989017535188, 32'sd0.05784521504363546, 32'sd0.02882245783592832, 32'sd0.024794451962383522, 32'sd0.060374670079398444, 32'sd0.020668259478816474, 32'sd0.0151532536307374, 32'sd0.10200276405168372, 32'sd-0.07640803465801822, 32'sd-0.11567396956873541, 32'sd0.028496469125194678, 32'sd-0.018475404639226093, 32'sd-0.008754415179872818, 32'sd0.008218375500325498, 32'sd0.022852540469256572, 32'sd0.030916163937438422, 32'sd0.10624667958851779, 32'sd-2.983131152864126e-120, 32'sd-9.82388650721402e-121, 32'sd-7.335769603904561e-126, 32'sd-2.61490555766447e-126, 32'sd-0.020701702351195506, 32'sd0.00977581443824073, 32'sd-0.014039725964486768, 32'sd0.004336410723002976, 32'sd-0.012496499096202216, 32'sd0.08946238573718909, 32'sd0.08871636566992613, 32'sd-0.008215617151668398, 32'sd0.1031499239705495, 32'sd0.07435691239883724, 32'sd0.014876118911359535, 32'sd0.06596405806046055, 32'sd-0.11782863323763702, 32'sd-0.09558216116528766, 32'sd-0.02664772336730128, 32'sd-0.09703366938495467, 32'sd-0.0908250209819781, 32'sd-0.07798166605877535, 32'sd-0.01593636993150547, 32'sd0.0016949840412586819, 32'sd0.001148073817103978, 32'sd0.04377540057667142, 32'sd0.013929508503950224, 32'sd0.031730435342535036, 32'sd0.07411404879154981, 32'sd6.880203873918201e-122, 32'sd6.119978404549707e-118, 32'sd0.05475231660574604, 32'sd0.08477331616536612, 32'sd0.10820029488520148, 32'sd-0.0009155749773686678, 32'sd0.04015608536574591, 32'sd0.01101829668569373, 32'sd0.07173774366924818, 32'sd0.007951122199559553, 32'sd-0.0769014834121, 32'sd0.0767388989263398, 32'sd0.05152089024761498, 32'sd0.09318760660705379, 32'sd0.03532285411052876, 32'sd0.09592517126306235, 32'sd-0.019257624955268535, 32'sd-0.059776632820004505, 32'sd-0.15470360223857738, 32'sd-0.2236540340921608, 32'sd-0.1700263760845825, 32'sd-0.1568171685166035, 32'sd0.006288381292205706, 32'sd0.015193467842326948, 32'sd-0.022235947356554327, 32'sd0.02085341054134747, 32'sd-0.08692481687827346, 32'sd-0.0008059743561951474, 32'sd0.04861890642083025, 32'sd2.0473681049876526e-119, 32'sd0.09135188613858496, 32'sd-0.014462739702378088, 32'sd-0.04744384315396397, 32'sd-0.03436050929640463, 32'sd0.13569335778094627, 32'sd0.13024506323492305, 32'sd-0.004746430051137911, 32'sd-0.0001364025811169127, 32'sd0.04809188455085133, 32'sd0.07497302106122089, 32'sd0.0643394078744287, 32'sd0.14214478085308635, 32'sd0.050205356000634395, 32'sd0.013546103370632046, 32'sd0.07413386151885905, 32'sd-0.06717111626123544, 32'sd-0.16335879918347107, 32'sd-0.12667825911121977, 32'sd-0.09535829253298603, 32'sd-0.18936318152519838, 32'sd-0.07559430105347968, 32'sd-0.04059682409966104, 32'sd-0.0407135662053447, 32'sd-0.10838880605122829, 32'sd-0.020669382204556472, 32'sd-0.10193297029499382, 32'sd0.07964035631445099, 32'sd-4.141139371607207e-124, 32'sd0.08635589967577649, 32'sd0.01920898829316711, 32'sd0.05089749668373787, 32'sd-0.12131327094349455, 32'sd0.004103647878469937, 32'sd0.03770669621641751, 32'sd0.025196406365162488, 32'sd0.04067084482394789, 32'sd-0.06561628690915276, 32'sd0.006926611941593227, 32'sd-0.025849526175178102, 32'sd0.021081325461937445, 32'sd-0.015193440196650825, 32'sd-0.00027302466503810566, 32'sd-0.016820573477461527, 32'sd0.0597465034676944, 32'sd-0.05117881511754811, 32'sd-0.07846942357038324, 32'sd-0.12628622812897908, 32'sd-0.20345541809706827, 32'sd-0.17544315437094068, 32'sd-0.24013852826821264, 32'sd-0.1322409200554589, 32'sd-0.052588401780645236, 32'sd0.12108143287064733, 32'sd-0.015739609838351223, 32'sd-0.003980703453553593, 32'sd0.11634969194308377, 32'sd-0.029744233314728773, 32'sd0.04416938990532309, 32'sd0.08018990538711655, 32'sd-0.08084125869376502, 32'sd-0.09430085370366267, 32'sd-0.014076200169658467, 32'sd-0.021230498843434878, 32'sd0.015997385235483556, 32'sd0.0634321105514987, 32'sd0.07092664792067752, 32'sd0.010435874944754453, 32'sd0.04622803605830431, 32'sd0.04796192226005909, 32'sd0.07699421158731441, 32'sd-0.08155205323325979, 32'sd0.07258198971301595, 32'sd-0.14124417281702095, 32'sd-0.13722444200341644, 32'sd-0.3015345314701387, 32'sd-0.1482408699779081, 32'sd-0.17088825599930163, 32'sd-0.09406792638341961, 32'sd-0.13754703071940877, 32'sd0.08414723580462732, 32'sd0.12321043731462004, 32'sd-0.038923082108988434, 32'sd-0.05026450053311773, 32'sd0.003022275567265462, 32'sd-0.008765586148495352, 32'sd0.04729362194429485, 32'sd0.03432631547922477, 32'sd-0.044198613348325436, 32'sd-0.11248094304629352, 32'sd-0.006919230856235845, 32'sd-0.10416814683353842, 32'sd-0.06062339661395003, 32'sd-0.027214018253147537, 32'sd0.05534219283678046, 32'sd-0.034917111241105823, 32'sd0.10441136581755005, 32'sd0.04274077036422803, 32'sd0.09693537141355604, 32'sd0.12841073588172575, 32'sd0.05596581013867594, 32'sd0.054259702455218065, 32'sd-0.020067100665753835, 32'sd-0.07847753996783685, 32'sd-0.1861698525063069, 32'sd-0.10538755322193852, 32'sd-0.0031072432202163044, 32'sd-0.09969850610739013, 32'sd0.04338490493851518, 32'sd-0.12949143949546074, 32'sd0.011339689856805675, 32'sd0.009335175365811906, 32'sd0.05697589774513563, 32'sd0.04676282311828587, 32'sd-0.016343938643492144, 32'sd-0.08180751125883945, 32'sd-0.041268211385290306, 32'sd0.15320794505566718, 32'sd-0.05776719524221968, 32'sd0.05950122553242754, 32'sd-0.07955897204730111, 32'sd0.06959059980125348, 32'sd0.11502306529439496, 32'sd0.014692439635017106, 32'sd0.09884477338105113, 32'sd0.2549701121749687, 32'sd0.241585284706282, 32'sd0.22668489250306137, 32'sd0.2713926512638182, 32'sd0.07994485285666063, 32'sd-0.04047571280720252, 32'sd-0.14537143596210123, 32'sd-0.17836230207355305, 32'sd-0.13837992021047021, 32'sd0.08415185053219983, 32'sd0.060839336322136846, 32'sd0.14161465958585281, 32'sd-0.15467214919100614, 32'sd-0.03801390719077383, 32'sd-0.03443083951880581, 32'sd-0.03812567449794755, 32'sd-0.08459166754947381, 32'sd-0.0018117572603955992, 32'sd-0.11461817333308215, 32'sd-0.01264527434128302, 32'sd0.1178218793242719, 32'sd-0.004284674394967146, 32'sd0.015113545803578465, 32'sd-0.07110495190872254, 32'sd-0.021197612883063457, 32'sd0.17571745937268374, 32'sd0.18897437059605762, 32'sd0.2622263768031128, 32'sd0.2178347556251215, 32'sd0.17626154270266473, 32'sd0.12788957124532746, 32'sd0.1380868099385653, 32'sd0.06081341752846772, 32'sd-0.0035016839174019754, 32'sd-0.20456443734587462, 32'sd-0.24073973447205554, 32'sd-0.03611855254820098, 32'sd0.13985365448220294, 32'sd0.14383956806142872, 32'sd0.062440107403499874, 32'sd-0.1426063552131076, 32'sd0.006272736523505305, 32'sd0.05501699608301536, 32'sd0.07548631217201644, 32'sd0.06560517724348199, 32'sd0.026474903310481603, 32'sd0.006924857359155809, 32'sd-0.08345345283752058, 32'sd-0.05847255838263068, 32'sd-0.039747463670758536, 32'sd0.08374394924607288, 32'sd0.009330104634173893, 32'sd0.021368696025951504, 32'sd0.22085404888163115, 32'sd0.10871458189583313, 32'sd0.03082627366707684, 32'sd0.12679074605415833, 32'sd0.07038989141640313, 32'sd0.04603389291629651, 32'sd-0.07437218713678832, 32'sd0.20499258162092449, 32'sd0.1889944867069044, 32'sd-0.07984547622660827, 32'sd-0.21057369319659625, 32'sd-0.22035114637875935, 32'sd-0.04107794380610519, 32'sd0.162657972191775, 32'sd0.0782389988372405, 32'sd-0.037992601357379585, 32'sd0.013884932480830215, 32'sd-0.011173026383206957, 32'sd0.013994457495339487, 32'sd0.08036977127343739, 32'sd0.005993532743019517, 32'sd0.05283924997038535, 32'sd-0.019915245504960592, 32'sd0.02652178268889687, 32'sd-0.003294322419931618, 32'sd-0.14998484202973436, 32'sd-0.14151956950062838, 32'sd0.012513822774137673, 32'sd0.006515512362643675, 32'sd-0.10664574537785756, 32'sd-0.05725482169841819, 32'sd0.03656988707147589, 32'sd0.06101584390940207, 32'sd0.03356059206733331, 32'sd0.05666791484961681, 32'sd0.20922974128562719, 32'sd0.0314888905276246, 32'sd-0.17893889031230717, 32'sd-0.27834319343784686, 32'sd-0.2283363323363463, 32'sd-0.07969224968640276, 32'sd-0.011882866801276756, 32'sd0.012088725891600215, 32'sd0.021705241284808573, 32'sd0.03326614938005242, 32'sd0.060729818076403014, 32'sd0.06929687336856613, 32'sd0.05576266671639005, 32'sd-0.03285023267531259, 32'sd-0.1100352442889891, 32'sd-0.025336479399447522, 32'sd-0.17986522036699584, 32'sd-0.036406751888368824, 32'sd-0.09206298923626173, 32'sd-0.0864186918986662, 32'sd-0.0734253847629753, 32'sd-0.045578998794399764, 32'sd-0.009573211402049926, 32'sd-0.1337614160335483, 32'sd-0.07541030387673787, 32'sd0.06457352137817758, 32'sd0.02687875739479233, 32'sd0.06144805125514232, 32'sd0.13995127519335313, 32'sd-0.07548593978611585, 32'sd-0.1746513386892681, 32'sd-0.1795756390323663, 32'sd-0.11726835085246051, 32'sd0.013952541096552709, 32'sd0.03919262138226784, 32'sd0.1572589641866257, 32'sd0.01799168588730708, 32'sd0.07572836459069873, 32'sd0.006473558049355287, 32'sd0.03141792254180371, 32'sd-0.05705709683052832, 32'sd-0.01541698984050126, 32'sd-0.08035298643188026, 32'sd0.05044484177673525, 32'sd-0.08688665700637571, 32'sd-0.1711248384666617, 32'sd-0.09196283076602059, 32'sd-0.11222680671027811, 32'sd-0.06978778205518851, 32'sd0.019934137996455235, 32'sd-0.06286049532025996, 32'sd-0.04105520693563586, 32'sd-0.08325153120175868, 32'sd0.009973664878844416, 32'sd-0.07688378814138652, 32'sd0.10305642861600268, 32'sd0.04734353042489805, 32'sd0.006204997636278477, 32'sd-0.140400846075747, 32'sd-0.1672468491068541, 32'sd-0.005881611389938425, 32'sd-0.07001865704543267, 32'sd0.10196647240636265, 32'sd0.015938852571898216, 32'sd-0.06565540855771904, 32'sd0.0008636848089114451, 32'sd0.017301305375246923, 32'sd0.018107998063578844, 32'sd-0.07656773607164191, 32'sd-0.024404545263340394, 32'sd-0.03741697054246117, 32'sd0.09171931460016738, 32'sd-0.023368473121445982, 32'sd-0.08841255363762719, 32'sd-0.1469986788720148, 32'sd-0.07958084206642652, 32'sd-0.027897300986169406, 32'sd-0.11624951017717505, 32'sd-0.05489569119422119, 32'sd-0.019184358836628855, 32'sd0.03759866370943122, 32'sd-0.04754966413260615, 32'sd0.02429545287243695, 32'sd-0.016240395499274387, 32'sd0.05953357502675224, 32'sd-0.13163148270760155, 32'sd-0.10549712633779358, 32'sd-0.07095812662095524, 32'sd-0.10569368385419023, 32'sd-0.07230559739734214, 32'sd0.009002569723509907, 32'sd0.056840047324040424, 32'sd-0.11788488774262491, 32'sd-0.053451067974669565, 32'sd0.0930611012989523, 32'sd0.08627306387798449, 32'sd0.1333244427041039, 32'sd-0.005425030466647699, 32'sd-0.0005543090616517901, 32'sd0.01325554861948168, 32'sd-0.040818137361598256, 32'sd0.03812452100867457, 32'sd-0.024111113534717205, 32'sd-0.0641082204043959, 32'sd0.06983629757336761, 32'sd0.007504048458463253, 32'sd-0.001195858680596752, 32'sd0.10461018128868821, 32'sd0.05143046164445131, 32'sd0.008212973701807071, 32'sd-0.037155007072791346, 32'sd0.050601100733931384, 32'sd-0.03702336237730689, 32'sd-0.06997520462032657, 32'sd-0.054895984984417924, 32'sd-0.08079693817444349, 32'sd0.011061497197189546, 32'sd0.008659290549262403, 32'sd0.006067559924686429, 32'sd0.11409569291408304, 32'sd-0.03183221624147664, 32'sd-0.014861529969461768, 32'sd0.0925299520442231, 32'sd-1.3317448070437422e-127, 32'sd0.01809051669380048, 32'sd0.05174717317141287, 32'sd0.06765259087277156, 32'sd0.027892390956059714, 32'sd0.05616172315016061, 32'sd0.04469982233134456, 32'sd-0.09919670756604144, 32'sd-0.030432739207445644, 32'sd0.11023900840405318, 32'sd-0.040623404330958714, 32'sd0.04249402338682927, 32'sd-0.03581495580740073, 32'sd-0.03257229604087954, 32'sd0.007705129838434225, 32'sd-0.015955278021524306, 32'sd0.003806011094668615, 32'sd-0.06278168212392121, 32'sd-0.0005997891612189517, 32'sd0.028256157560887958, 32'sd-0.0016512002694773092, 32'sd-0.04623924118738968, 32'sd-0.06489141060693322, 32'sd0.09012753127553692, 32'sd0.008929089673619292, 32'sd0.12050554093165788, 32'sd0.08164190284198537, 32'sd0.007109917866425079, 32'sd-0.022999550105635393, 32'sd0.019113873395786123, 32'sd0.00015067048246598133, 32'sd-0.04692139884180896, 32'sd0.003311371993969328, 32'sd0.04161240779490336, 32'sd0.05850341643959095, 32'sd0.007109529998693456, 32'sd-0.0703905434477639, 32'sd-0.05300778376374021, 32'sd-0.023401738589733056, 32'sd0.0493297379826105, 32'sd-0.06398225476690879, 32'sd0.06356568714876698, 32'sd-0.0014280429001042728, 32'sd-0.0009312026116212835, 32'sd-0.0008002259137075176, 32'sd-0.010706176942233315, 32'sd-0.0012596168903819302, 32'sd0.05233982081012342, 32'sd-0.002686483406381915, 32'sd-0.0007431212356826284, 32'sd0.1426036572712372, 32'sd0.16544731037394453, 32'sd0.05583231444445328, 32'sd0.042757224906308504, 32'sd0.09437946378100286, 32'sd-0.03484226279750893, 32'sd0.022413751372380577, 32'sd0.0536052955884732, 32'sd-0.0634944459017414, 32'sd-0.09647287328127482, 32'sd0.01663960620078141, 32'sd0.0431902136620193, 32'sd0.05439010539230484, 32'sd0.14520421452136098, 32'sd-0.014731537754298866, 32'sd-0.1231140177172218, 32'sd0.03447898727657253, 32'sd-0.09466593826290662, 32'sd-0.0138787184978088, 32'sd0.0827902234231424, 32'sd0.059783888024833344, 32'sd0.0017550685006847103, 32'sd0.08348451512115095, 32'sd-0.021437430236515644, 32'sd0.015394345706586881, 32'sd0.04015631088156422, 32'sd0.07362812870148427, 32'sd0.032126906013209396, 32'sd0.1325987441384278, 32'sd0.1314898547524843, 32'sd-0.0045298201519221185, 32'sd-0.0015561636285638682, 32'sd0.05183163654169396, 32'sd-0.07851592252240007, 32'sd4.164589377515839e-115, 32'sd0.02443965076797503, 32'sd0.007583965576097922, 32'sd-0.09808355592969474, 32'sd-0.031784826189472884, 32'sd0.10128489821929336, 32'sd-0.023862035633216122, 32'sd-0.008280731432585915, 32'sd-0.09279224057185054, 32'sd-0.10641946474206247, 32'sd-0.00825309215547621, 32'sd0.011987140509654319, 32'sd0.11219877445347308, 32'sd0.09999109696865326, 32'sd-0.009417084415361165, 32'sd0.004451415402962036, 32'sd0.11683543796520528, 32'sd0.009555169785294911, 32'sd0.04930205670254005, 32'sd-0.06672172689164813, 32'sd0.05047126304571785, 32'sd0.06669241217885814, 32'sd0.14607494785230876, 32'sd-0.0022574884127065623, 32'sd0.009256503984836833, 32'sd-0.04877446738148952, 32'sd0.005657912211648113, 32'sd0.06530169318850376, 32'sd0.09775658467723344, 32'sd0.03963648863459088, 32'sd-0.039480557676713636, 32'sd-0.029082912516050715, 32'sd0.04204747953225794, 32'sd-0.02614280947986948, 32'sd0.13354326216030782, 32'sd-0.06353249338767718, 32'sd-0.03702786052636971, 32'sd-0.0025510630487637844, 32'sd0.0540204705190055, 32'sd-0.055115415888438705, 32'sd0.019139547026731898, 32'sd0.03053066649374842, 32'sd0.03546567271933386, 32'sd0.027784516963035286, 32'sd-0.028046214049315378, 32'sd-0.07376285347781249, 32'sd0.06649214747348234, 32'sd-0.060768077396462075, 32'sd-0.02376301956609863, 32'sd0.10679282403205363, 32'sd0.029300325990017466, 32'sd0.06362678486435736, 32'sd-0.07947614396129614, 32'sd-0.07625874042297857, 32'sd-0.02835300006990394, 32'sd0.07597605631335703, 32'sd0.04273924404466747, 32'sd0.002354970635105414, 32'sd0.044647292848183806, 32'sd0.09912358373660715, 32'sd0.11816427694155529, 32'sd-0.02995823314916449, 32'sd-0.04269596987347953, 32'sd0.019286020145527365, 32'sd0.07561064434709498, 32'sd-0.02538881694696177, 32'sd0.006856902134715176, 32'sd-0.08240709899300415, 32'sd0.03908229113218427, 32'sd0.009835136063578586, 32'sd0.07172468528126875, 32'sd-0.017610858982987646, 32'sd-0.02304931813657769, 32'sd-0.07788612082303456, 32'sd-0.04267092432580592, 32'sd-0.10494587355903792, 32'sd0.07359218540016627, 32'sd0.09572223523207697, 32'sd0.1319620570364074, 32'sd0.10552102058694804, 32'sd0.06834955947402044, 32'sd-0.047891174555842506, 32'sd-0.08737365798718827, 32'sd0.10508450584310823, 32'sd-2.754865837651332e-118, 32'sd0.07810133539183983, 32'sd0.0579417592698703, 32'sd0.019799965648815532, 32'sd-0.02685708705937438, 32'sd0.017425962879291657, 32'sd-0.01488362823935695, 32'sd-0.05237161147589818, 32'sd-0.020559906013044176, 32'sd-0.03385473117078874, 32'sd-0.05437575849683429, 32'sd-0.07420370134367764, 32'sd0.06549721519701467, 32'sd0.0692395383596009, 32'sd-0.0050707900251440174, 32'sd0.15572962485286526, 32'sd-0.05033468944074206, 32'sd0.04930427259889543, 32'sd0.021879361261310543, 32'sd-0.04478429153700116, 32'sd0.10785659069464924, 32'sd0.09067832649766543, 32'sd0.002668962775294076, 32'sd0.05875060900954338, 32'sd0.055050585714525375, 32'sd0.060943808968817306, 32'sd-0.06725764811576777, 32'sd-1.0447250494636279e-122, 32'sd3.2697581698324865e-119, 32'sd-2.39778456239581e-124, 32'sd0.07222935226176523, 32'sd0.09171981978723037, 32'sd0.015068317263998349, 32'sd0.018025764153119083, 32'sd-0.04153565197719983, 32'sd-0.10415176721761535, 32'sd-0.04463245279145286, 32'sd-0.1432172817354676, 32'sd-0.164196606861431, 32'sd-0.07085817458350915, 32'sd0.06398307238434105, 32'sd-0.027439420725379804, 32'sd-0.04677639753667928, 32'sd0.058700837663348604, 32'sd0.01495327265298917, 32'sd-0.0024991716611578517, 32'sd0.10333232713596577, 32'sd0.03516208833973211, 32'sd0.0029379994360320305, 32'sd0.05885566475826195, 32'sd-0.035229305716102145, 32'sd0.15528161119858522, 32'sd-0.008559621209282314, 32'sd0.03182069461654654, 32'sd0.04208889168497349, 32'sd1.5123563423554708e-124, 32'sd3.369585500187543e-125, 32'sd6.069804113538472e-124, 32'sd0.053053777130142796, 32'sd-0.009673073834862853, 32'sd-0.0852555445062686, 32'sd0.059556749149684306, 32'sd0.05059890320747449, 32'sd0.1498776375330809, 32'sd0.08703884677519552, 32'sd-0.16569718914523096, 32'sd-0.146422439812081, 32'sd-0.15128498016777012, 32'sd-0.05909972427248766, 32'sd0.008388005755953921, 32'sd-0.048831365508689134, 32'sd0.06024425861479107, 32'sd0.07355149256615866, 32'sd0.06492779358797572, 32'sd0.008322670139957659, 32'sd-0.06504334589012346, 32'sd0.007913160636412533, 32'sd-0.0701744974651273, 32'sd-0.030904675244184637, 32'sd-0.03927363195755659, 32'sd-0.08272238587803381, 32'sd0.022022263204803768, 32'sd-0.0055065863752297006, 32'sd1.9172957983169672e-122, 32'sd1.384219939409065e-115, 32'sd6.897282789283032e-124, 32'sd2.8418265630275887e-116, 32'sd0.07018317790493574, 32'sd-0.07197320092267116, 32'sd0.08665626332988371, 32'sd0.05062688193367011, 32'sd0.042042287884055424, 32'sd0.030992751111111227, 32'sd-0.05788307745055325, 32'sd0.09419676838134368, 32'sd-0.07430765708634651, 32'sd0.15115677283027149, 32'sd0.1151238563304514, 32'sd-0.009926252503157405, 32'sd-0.024217544232807735, 32'sd-0.08373513156051599, 32'sd-0.020276443062410124, 32'sd-0.11038075531688214, 32'sd0.06585655770360199, 32'sd-0.013446754597575286, 32'sd0.06147282741672402, 32'sd0.01747756979146766, 32'sd0.017035044142271565, 32'sd0.08308934956381514, 32'sd0.07564289052749541, 32'sd4.9207062966995215e-118, 32'sd-6.7373381884488e-126, 32'sd2.916666142544628e-120, 32'sd1.8938564334847027e-122, 32'sd1.4980869331957467e-119, 32'sd-3.198417339170594e-116, 32'sd0.13662163951909864, 32'sd-0.01522042471835825, 32'sd0.09776623852387736, 32'sd0.03942850440044705, 32'sd0.0660283937607311, 32'sd0.01598810582914146, 32'sd0.012441127913562748, 32'sd-0.037660678332848675, 32'sd0.10413724633360033, 32'sd0.05640063061958567, 32'sd-0.015700306238580063, 32'sd0.0007284544781208668, 32'sd0.03512204465870242, 32'sd0.07813672478999296, 32'sd0.04497031592624485, 32'sd0.0317317932263529, 32'sd0.02690137433923709, 32'sd0.08044230043462901, 32'sd0.06223989463362932, 32'sd0.16987435379355706, 32'sd2.5260040990056605e-118, 32'sd3.3155083195679256e-126, 32'sd-1.0612851339749058e-121, 32'sd2.0404527663431947e-116},
        '{32'sd-3.691596025398718e-126, 32'sd3.247544060013283e-116, 32'sd-1.1120358595883032e-121, 32'sd1.2794627006674137e-118, 32'sd-3.611158827267956e-119, 32'sd-2.260851355179342e-127, 32'sd-2.8133482698625406e-122, 32'sd-1.665380521543552e-124, 32'sd-7.519231978482965e-115, 32'sd-2.5682676323723394e-124, 32'sd-2.6665864317610886e-119, 32'sd7.442853115361979e-128, 32'sd0.03422289751889902, 32'sd0.10339777126910078, 32'sd-0.018882948123389896, 32'sd0.045433188224192164, 32'sd-4.0693430464433445e-127, 32'sd3.0206671734684557e-125, 32'sd-2.753079010940175e-125, 32'sd5.483322128559259e-124, 32'sd6.37871526734636e-126, 32'sd-2.5961544390360393e-120, 32'sd-1.0331297619188674e-115, 32'sd-3.8411981098992785e-119, 32'sd1.8233589323402028e-119, 32'sd-2.9555699602263235e-123, 32'sd5.18208238893261e-120, 32'sd1.4937340406065322e-115, 32'sd8.42572234549031e-127, 32'sd-3.599171181679904e-116, 32'sd-2.168521162533651e-118, 32'sd-8.449688658790043e-117, 32'sd-0.0027006633110682756, 32'sd0.04231042709517362, 32'sd-0.032765276981675355, 32'sd-0.046450948529211104, 32'sd0.02355661597712818, 32'sd0.06732493474628702, 32'sd-0.0034612577475612544, 32'sd0.007751332165743295, 32'sd-0.11461860101463243, 32'sd0.013675936920749017, 32'sd0.053143826501780574, 32'sd0.032249247024900014, 32'sd-0.021849280129157746, 32'sd0.11774269608885533, 32'sd0.12175731986040915, 32'sd0.004507573494491608, 32'sd-0.017418949032051365, 32'sd0.012125649030933102, 32'sd0.06645665285352612, 32'sd-0.002052032485127951, 32'sd-8.525875049717169e-117, 32'sd-1.2115622229033698e-127, 32'sd-4.3285150537197325e-125, 32'sd-3.295445837360441e-118, 32'sd2.6158542637574524e-114, 32'sd-1.005592272020524e-115, 32'sd0.03449427032821496, 32'sd0.07871673803974666, 32'sd-0.034172124454468995, 32'sd0.0035302063852418897, 32'sd-0.004147388467027172, 32'sd0.035947192702080986, 32'sd-0.06432877307724899, 32'sd-0.08116548423653024, 32'sd0.04491964764294262, 32'sd-0.08216501412292665, 32'sd-0.010530358659264095, 32'sd0.07072544750534236, 32'sd-0.1096751723516081, 32'sd0.013071632476069352, 32'sd0.06717007178720603, 32'sd0.11208233044741328, 32'sd0.07588506218131866, 32'sd-0.006884170498383836, 32'sd0.06644942681526468, 32'sd0.026486526832067005, 32'sd0.012540390875301783, 32'sd-0.02774327187707049, 32'sd0.010662141443598432, 32'sd0.04318332512128386, 32'sd7.314932680407195e-120, 32'sd2.5041842654258447e-119, 32'sd-6.224254351895555e-126, 32'sd-1.6506762778695435e-123, 32'sd0.030331714377228026, 32'sd-0.040797358959050435, 32'sd0.06757611084400619, 32'sd0.031010695917090624, 32'sd-0.004642283041588308, 32'sd-0.06854865631900113, 32'sd-0.10373170024777723, 32'sd-0.06084240771637418, 32'sd-0.12079564018364823, 32'sd-0.10256570253801282, 32'sd-0.15485257892540905, 32'sd-0.10824915646748179, 32'sd-0.10451666116373459, 32'sd0.12494902540035048, 32'sd0.06944633590222395, 32'sd0.0579913652594024, 32'sd0.0436823782610117, 32'sd-0.08171638192264273, 32'sd0.03783515873437488, 32'sd-0.02059205553423879, 32'sd-0.038271142817589004, 32'sd0.043498985768600784, 32'sd-0.04388317127721306, 32'sd0.05205973828102503, 32'sd-0.06998429984371751, 32'sd-3.0205043183457756e-123, 32'sd-7.392541329497035e-123, 32'sd0.007385467805150003, 32'sd-0.03791360161113988, 32'sd-0.025425692723591943, 32'sd-0.004474136584133408, 32'sd-0.09496701173979664, 32'sd-0.08185066816079141, 32'sd-0.021948452132208973, 32'sd-0.03843258710476169, 32'sd0.07954296333904014, 32'sd-0.0758988867494828, 32'sd0.013832799875550954, 32'sd-0.008642529456431037, 32'sd-0.05988720858000298, 32'sd-0.07643322848834674, 32'sd-0.04088179587971139, 32'sd0.11910941500513657, 32'sd-0.04080224357704162, 32'sd-0.08523918037020724, 32'sd-0.02402520851186853, 32'sd0.09257022122334095, 32'sd0.10783546645278226, 32'sd0.028624227078082983, 32'sd-0.021863206594889984, 32'sd0.03031872688119023, 32'sd-0.018441247264484182, 32'sd-0.02313468625978355, 32'sd0.017947341339493723, 32'sd-2.1200732024568227e-114, 32'sd-0.007423536906792104, 32'sd0.036683988261966845, 32'sd0.015026939910998927, 32'sd0.01564157140754466, 32'sd0.038953360800673326, 32'sd0.008275329225566612, 32'sd0.03148961270987287, 32'sd0.028759596303513126, 32'sd-0.05481715739531787, 32'sd0.0006429537303038249, 32'sd0.00922587256857676, 32'sd-0.12719602603973773, 32'sd-0.026741676393637153, 32'sd0.008429759688853991, 32'sd0.05511440707086109, 32'sd0.033863797269377785, 32'sd0.05623559425625759, 32'sd0.1067574970551071, 32'sd0.17671771509278802, 32'sd-0.01495542920669392, 32'sd-0.06400913071063138, 32'sd0.055787407506903045, 32'sd-0.14597299315852955, 32'sd0.022717650544382444, 32'sd0.079126603391574, 32'sd0.07916677630976482, 32'sd0.031548458934113115, 32'sd6.771990620327682e-125, 32'sd0.006146198433552238, 32'sd-0.03487671503923443, 32'sd0.07634212954076448, 32'sd-0.04795621998863697, 32'sd0.012341062916871313, 32'sd-0.034973248707861865, 32'sd0.012955151026770563, 32'sd0.01704637912956551, 32'sd0.057693909976175586, 32'sd-0.0598023836021764, 32'sd-0.0855034758272284, 32'sd-0.08599317390010265, 32'sd-0.12232400079140276, 32'sd-0.1310834970351543, 32'sd0.03274984464774971, 32'sd-0.001599033637780074, 32'sd0.05870881935257975, 32'sd-0.060318582225513784, 32'sd5.031540020736189e-05, 32'sd0.01657741637469054, 32'sd-0.04032249389379923, 32'sd0.022107922489541704, 32'sd-0.04107985839275657, 32'sd-0.04332560812880245, 32'sd-0.15373513822742554, 32'sd-0.006093533989826526, 32'sd-0.0867104573838907, 32'sd0.0449899113489754, 32'sd0.03203985516050649, 32'sd0.07603673750003183, 32'sd-0.05660289312084307, 32'sd-0.01265263855580187, 32'sd0.030112843851772337, 32'sd-0.006420847193018004, 32'sd0.0819394670209371, 32'sd-0.04106101393482158, 32'sd0.07364595023651996, 32'sd-0.07110175905464043, 32'sd0.0019381512937918992, 32'sd0.09519081242728675, 32'sd-0.010501725441529832, 32'sd0.01094706033297814, 32'sd0.06070663485290041, 32'sd0.18176609923417547, 32'sd0.10593580031215892, 32'sd-0.01942217546570766, 32'sd-0.061130776974695496, 32'sd-0.13923938669966446, 32'sd0.057891842713763, 32'sd-0.03544612178445664, 32'sd0.10617491430669883, 32'sd0.06665715576259161, 32'sd-0.010040102305782745, 32'sd-0.021075680907685218, 32'sd0.08861835115341705, 32'sd0.004158510902748696, 32'sd0.028127878999640754, 32'sd0.0574130206743456, 32'sd-0.09276661982264779, 32'sd0.01786992933159678, 32'sd-0.09409175947097329, 32'sd0.04234621162496072, 32'sd-0.011093195366658842, 32'sd-0.07266913309918809, 32'sd-0.10085272110759694, 32'sd0.06585836721851161, 32'sd0.04121008869420988, 32'sd-0.08841684055987709, 32'sd-0.06904800007766494, 32'sd-0.08744980835830404, 32'sd0.06872472987167313, 32'sd0.024124257802411654, 32'sd0.08835472683791126, 32'sd-0.024831601913215214, 32'sd-0.052210160801982604, 32'sd-0.05066166792343123, 32'sd-0.03280023658286199, 32'sd0.029600030280542988, 32'sd0.05910372883590988, 32'sd-0.04977869917434123, 32'sd0.03939455542573146, 32'sd0.12129292353994332, 32'sd-0.05165967663714944, 32'sd0.024631974996483088, 32'sd-0.014946997965472735, 32'sd0.11565020719595943, 32'sd0.04879757426320254, 32'sd-0.015337535202910308, 32'sd0.031948791044589975, 32'sd-0.03066500555723915, 32'sd0.015114435052908584, 32'sd-0.06738431375650925, 32'sd0.050144246936626176, 32'sd-0.05712403385442289, 32'sd-0.03166343790543674, 32'sd-0.10938421447555385, 32'sd-0.06496525209837768, 32'sd-0.05762138928896786, 32'sd-0.17410178304509097, 32'sd-0.08450878039213207, 32'sd0.04446393048834647, 32'sd-0.035712946219544045, 32'sd0.10137666905297643, 32'sd0.18749816340529102, 32'sd-0.043862542566606766, 32'sd-0.023216735964574416, 32'sd0.010317838202927193, 32'sd-0.0029344714097391434, 32'sd0.14742483443909665, 32'sd-0.038169226945612734, 32'sd0.04892087359971389, 32'sd0.05500866285367133, 32'sd0.08733940729678408, 32'sd0.06889598108100355, 32'sd-0.03526124664062683, 32'sd-0.04158488418040325, 32'sd0.011772429456005602, 32'sd-0.0018008889503767164, 32'sd-0.03584372488507679, 32'sd-0.08054950217484033, 32'sd0.0233749013105694, 32'sd0.03911453447067372, 32'sd0.030141667109722478, 32'sd-0.05278965454179091, 32'sd-0.08891947654126738, 32'sd-0.15592174778521375, 32'sd-0.1444071488984405, 32'sd-0.09765928204572284, 32'sd0.018067286052274693, 32'sd0.06348119706081205, 32'sd0.09456043887909452, 32'sd0.08576119494370738, 32'sd0.033901043384440915, 32'sd-0.0679186590639139, 32'sd-0.023486893013828718, 32'sd0.07312444909331012, 32'sd0.13687504687518523, 32'sd-0.009590475348107575, 32'sd-0.072906299603582, 32'sd0.04610824135118995, 32'sd0.008124928075075526, 32'sd0.004733944183468903, 32'sd0.11329084894828578, 32'sd-0.04162417523479408, 32'sd-0.035373954081935034, 32'sd0.0657975732501734, 32'sd0.06876717537629352, 32'sd-0.04500413573807466, 32'sd-0.09388162814432709, 32'sd0.05081415035875366, 32'sd-0.10512757690302804, 32'sd0.008583018740646367, 32'sd0.06317992192539866, 32'sd-0.056231196886847155, 32'sd-0.27527947906035116, 32'sd-0.18138164926544878, 32'sd-0.10162102520184899, 32'sd0.21340248941587964, 32'sd0.11430469101553382, 32'sd0.08029603464340224, 32'sd0.009182433128708952, 32'sd0.020712780763605956, 32'sd-0.00039733745260869813, 32'sd0.05174520066892251, 32'sd0.03174562315096038, 32'sd-0.042457273309687, 32'sd-0.00965978699217889, 32'sd0.013920880411485868, 32'sd0.09816671405570687, 32'sd0.02053032456199385, 32'sd-0.006353777274236903, 32'sd-0.08297127733618052, 32'sd-0.09973769253178154, 32'sd-0.06296386177285793, 32'sd-0.029184822863798653, 32'sd-0.051604086242920816, 32'sd-0.08223867868143549, 32'sd0.02689538225195245, 32'sd-0.03595501423476409, 32'sd-0.007017850219681806, 32'sd0.025636143421682092, 32'sd-0.07091485110108142, 32'sd-0.31784698919718246, 32'sd-0.12996315027314537, 32'sd-0.203737538144192, 32'sd0.07751672620691727, 32'sd0.08052870105449793, 32'sd0.10947661130536794, 32'sd-0.0060937903584499156, 32'sd-0.0596289006982442, 32'sd-0.10866166423414135, 32'sd-0.054170545313898255, 32'sd-0.02663653063268858, 32'sd-0.08354572875118639, 32'sd0.03479288308935882, 32'sd0.040573231501271366, 32'sd0.021741709127390804, 32'sd0.043998658575435494, 32'sd-0.048155526411652286, 32'sd-0.06628116698820898, 32'sd0.020660193276613975, 32'sd0.1547792313370699, 32'sd0.1534078352112051, 32'sd-0.041770640039197775, 32'sd0.07679495258300341, 32'sd-0.025001366069057944, 32'sd0.08663181435158543, 32'sd0.16311495668392073, 32'sd-0.08961938318334806, 32'sd-0.1637924735997743, 32'sd-0.22237859592218454, 32'sd-0.1811784405651894, 32'sd-0.03080711771176585, 32'sd-0.015290901848115544, 32'sd-0.04939653238457378, 32'sd-0.04490387915932631, 32'sd-0.017030231717271048, 32'sd-0.06300326063596898, 32'sd-0.019391666251353395, 32'sd-0.06049731114083462, 32'sd-0.028236329203061055, 32'sd0.02122269089638687, 32'sd0.08503600492151182, 32'sd-0.038152347731087694, 32'sd-0.03409107867511467, 32'sd0.06714402718199745, 32'sd-0.07622043305612258, 32'sd-0.04524606298613877, 32'sd0.034976859517109, 32'sd0.14345767401650167, 32'sd0.20081922779581726, 32'sd0.06181753743837276, 32'sd0.06390400976092364, 32'sd0.018976472340615537, 32'sd-0.001824927077616855, 32'sd0.04471891440408798, 32'sd-0.178973978307265, 32'sd-0.16072836472576796, 32'sd-0.184366738414742, 32'sd-0.2679175894788967, 32'sd-0.045953692972516745, 32'sd0.017042883821461543, 32'sd-0.10484640287395103, 32'sd-0.040406028190901305, 32'sd0.05411686646705082, 32'sd0.03268976066358848, 32'sd-0.008589809749958517, 32'sd-0.050666715967926115, 32'sd0.03801146018045336, 32'sd0.11313112414400435, 32'sd0.11594822569069801, 32'sd0.046076602701841586, 32'sd0.029903646315464383, 32'sd0.06866614508878231, 32'sd-0.07359772728440808, 32'sd0.009821206961787397, 32'sd0.05792066481146878, 32'sd0.1490941723588451, 32'sd0.06341640929432381, 32'sd0.030504825112418216, 32'sd0.15075612355404244, 32'sd0.1852356880678397, 32'sd0.07482066749774459, 32'sd0.023664733372575568, 32'sd-0.26060152456154395, 32'sd-0.13500166426747726, 32'sd-0.1097018062457674, 32'sd-0.055391558979182395, 32'sd0.09855396968022831, 32'sd0.037128631493289335, 32'sd0.0032913268734235594, 32'sd-0.03259901499184726, 32'sd0.01696452343116356, 32'sd-0.0411869842928625, 32'sd-0.05835206461575448, 32'sd0.1062504184333586, 32'sd-0.021803047678652755, 32'sd-0.005230618816470498, 32'sd0.0451377179727443, 32'sd0.009088451304505711, 32'sd0.003873945375370057, 32'sd-0.04419141674021022, 32'sd-0.08596258327883158, 32'sd0.0272096465323861, 32'sd0.031999876424017484, 32'sd0.026114239883173813, 32'sd-0.02297583192555948, 32'sd0.1495927131345375, 32'sd0.18882759812195904, 32'sd0.14444752130060243, 32'sd0.010899987452613238, 32'sd-0.053610816025075156, 32'sd-0.22572729042017897, 32'sd-0.10581712308977075, 32'sd0.00025938198450951714, 32'sd0.14687852109092792, 32'sd0.11070487371667286, 32'sd0.1857707384293334, 32'sd0.10808254525783033, 32'sd0.041626474715865495, 32'sd0.16994772728620416, 32'sd0.10298733739269436, 32'sd-0.038050654536824886, 32'sd0.005144585916344238, 32'sd-0.07546644048030567, 32'sd0.05117983499486324, 32'sd0.02503204233535085, 32'sd8.332427767608914e-116, 32'sd0.007240302463705168, 32'sd0.05021108009500004, 32'sd-0.04246953383794569, 32'sd-0.022262453981896368, 32'sd-0.01737414031702121, 32'sd0.0897692827077636, 32'sd0.06640022016415267, 32'sd0.12928377521055995, 32'sd0.08175917229537547, 32'sd0.04960036570607179, 32'sd0.003165372656009589, 32'sd-0.14327721148986644, 32'sd-0.0202481755953933, 32'sd0.10226813293966651, 32'sd0.10014915410332494, 32'sd0.2120774900995315, 32'sd0.11952977619437768, 32'sd0.043742944903344, 32'sd0.042324056032265654, 32'sd-0.033068364006011396, 32'sd0.135572772813919, 32'sd-0.020802225665551576, 32'sd0.05119891491049716, 32'sd0.061914629306383875, 32'sd-0.030659262586670656, 32'sd-0.029582332236297516, 32'sd0.10850722177120348, 32'sd0.03771289455570311, 32'sd0.00473083625149346, 32'sd-0.08868125156304159, 32'sd0.008081518801673643, 32'sd0.07616366132857803, 32'sd-0.004764324134286225, 32'sd0.021938949600251608, 32'sd0.1730462424361641, 32'sd0.20823850211871972, 32'sd0.2631027371226471, 32'sd0.03302837642269768, 32'sd-0.045009795544142445, 32'sd-0.062248253837702966, 32'sd-0.02126372331557947, 32'sd0.07458351879566816, 32'sd0.13635889145517627, 32'sd0.027690037783437715, 32'sd0.0005615442070481967, 32'sd0.16080845627851373, 32'sd0.0872020725031401, 32'sd0.166892233218392, 32'sd0.07526124045732395, 32'sd0.07622118585112929, 32'sd0.10710416247028852, 32'sd0.04548979625826522, 32'sd-0.016197201502617307, 32'sd0.03686979720325159, 32'sd0.07015482926631396, 32'sd-0.0149274970022066, 32'sd0.05312131398310348, 32'sd0.02843941010270655, 32'sd-0.02075702889772954, 32'sd0.001968788005278779, 32'sd0.02212669616201039, 32'sd0.0448913878443547, 32'sd0.07017636357397077, 32'sd0.12724412306711555, 32'sd0.05343157122157292, 32'sd0.027734563807514694, 32'sd-0.13896057680015186, 32'sd-0.16128571200912908, 32'sd0.0049061709446603895, 32'sd0.17582895345575955, 32'sd0.1494618331722781, 32'sd0.027738366768939288, 32'sd-0.019502001680365873, 32'sd-0.00826424742803067, 32'sd0.011298487770703471, 32'sd-0.0280454998851529, 32'sd0.10773750096358041, 32'sd-0.015282513170621181, 32'sd-0.014302492129089343, 32'sd-0.07330752331540236, 32'sd-0.030808438322666484, 32'sd0.0007134231849988426, 32'sd0.08338702856929849, 32'sd3.9025670474605493e-119, 32'sd0.07317791679174622, 32'sd0.07849045292418382, 32'sd0.02784788162879389, 32'sd0.031050675002443122, 32'sd-0.07175974661266118, 32'sd-0.04831792017980298, 32'sd0.11190685480178025, 32'sd0.0032181165825787613, 32'sd-0.03497077144401149, 32'sd0.04496972738412731, 32'sd0.0038475438053000625, 32'sd-0.09757024842948342, 32'sd-0.011632734841070988, 32'sd0.042840636076953126, 32'sd-0.023760180812890833, 32'sd-0.019526201687907235, 32'sd0.03440781485236294, 32'sd-0.019143476897073547, 32'sd-0.04032183640619908, 32'sd-0.03965913398495268, 32'sd0.019400919425715948, 32'sd0.03343505344719256, 32'sd-0.024044053742490742, 32'sd-0.007733433959506963, 32'sd-0.03043950820144615, 32'sd0.02730348874204821, 32'sd0.04564917266242634, 32'sd-0.039561250072575216, 32'sd-0.11162872020821939, 32'sd-0.038938908176236554, 32'sd0.03198041618574213, 32'sd0.10083002054102413, 32'sd0.07629752489400923, 32'sd0.025411769320357415, 32'sd0.08118786823998017, 32'sd-0.024453868025412415, 32'sd0.028920299069890517, 32'sd-0.028196251086484693, 32'sd-0.031276927115917126, 32'sd0.025075689306090863, 32'sd-0.08994030168622753, 32'sd-0.001817614957273712, 32'sd-0.006437005015378145, 32'sd-0.1905885047599342, 32'sd-0.06708496528520866, 32'sd-0.05946560766538111, 32'sd0.11136443019165876, 32'sd0.06744369294177623, 32'sd-0.002337272642098607, 32'sd0.12069777992964263, 32'sd0.0037742680830736932, 32'sd-0.038795767127192106, 32'sd-0.08052060345480609, 32'sd-0.07986223932695842, 32'sd0.029506858102719743, 32'sd0.03678301751989534, 32'sd-0.04638873016154172, 32'sd0.008811282810328615, 32'sd0.03913623282616355, 32'sd0.023790329872010157, 32'sd0.07391707518242192, 32'sd0.15352741138675136, 32'sd0.023168539078650664, 32'sd0.06778629343038967, 32'sd0.05980140387515106, 32'sd-0.07792929127179885, 32'sd-0.01213962159809279, 32'sd0.06507270457150006, 32'sd-0.10570135326869627, 32'sd-0.04433138247214175, 32'sd-0.19173288094197682, 32'sd-0.17805654456059142, 32'sd-0.11795718014466114, 32'sd0.008304986246041096, 32'sd0.09737601804022647, 32'sd-0.013150891226913698, 32'sd-0.03784770649942177, 32'sd0.012155489083473879, 32'sd-0.05801690729217164, 32'sd0.04929894688650756, 32'sd-0.08782169206680956, 32'sd-0.06532588744940757, 32'sd0.010655668359791062, 32'sd-7.065725805362786e-115, 32'sd0.04126020553077785, 32'sd0.03369579593656744, 32'sd0.048680035035910875, 32'sd-0.008718787562145738, 32'sd-0.05626411906716759, 32'sd-0.0618869250765195, 32'sd0.05709384098669437, 32'sd-0.04608524997334435, 32'sd-0.05810005974326581, 32'sd0.0019374239658565943, 32'sd0.1371933803154219, 32'sd0.033281190696892934, 32'sd-0.019471155226690354, 32'sd-0.058687601980274395, 32'sd-0.14145132137255895, 32'sd-0.18571569173170296, 32'sd-0.16696011983933515, 32'sd0.0291626960058291, 32'sd-0.0017321967782272585, 32'sd0.041868187541591675, 32'sd-0.05687657543761125, 32'sd-0.06651765337840894, 32'sd0.017619700287276503, 32'sd-0.02358947121575507, 32'sd0.014053994124140419, 32'sd-0.006039999498257295, 32'sd-2.616936875698102e-126, 32'sd-6.258575612010148e-124, 32'sd4.699378534944703e-124, 32'sd-0.0928821838552699, 32'sd-0.0010404012522715108, 32'sd0.0369118382109747, 32'sd-0.011685022729258232, 32'sd-0.020177458534697802, 32'sd0.014244532904460101, 32'sd-0.09358246076978197, 32'sd0.07258574727341924, 32'sd7.977139101482142e-06, 32'sd0.03386670592804795, 32'sd0.009621049633937407, 32'sd0.010564456861690054, 32'sd-0.09358822338024507, 32'sd-0.13132795163322325, 32'sd-0.1598968539751927, 32'sd-0.19415485868580662, 32'sd-0.1831301812532942, 32'sd-0.04929076650949126, 32'sd0.0047714284510591, 32'sd0.0020410445790397564, 32'sd-0.01575733797981145, 32'sd0.0021817838920960763, 32'sd0.005043819063699696, 32'sd0.09726148834155844, 32'sd-0.04431457739190166, 32'sd1.1107866514090574e-119, 32'sd5.315922926879245e-116, 32'sd3.871075051815319e-115, 32'sd0.007092922539716831, 32'sd0.034091256658658954, 32'sd-0.02084401879106588, 32'sd0.1359341026998994, 32'sd0.07254027321785021, 32'sd-0.0917844690158054, 32'sd-0.10164456810163074, 32'sd-0.10047632637969804, 32'sd-0.0826690443342244, 32'sd-0.0939426912898513, 32'sd0.002168882175667843, 32'sd-0.04553536718478294, 32'sd-0.10492683056396891, 32'sd0.026481340873887396, 32'sd-0.08325783932258678, 32'sd-0.08505917713871862, 32'sd-0.14516678327920185, 32'sd-0.05600336838495429, 32'sd-0.009098587453266287, 32'sd-0.06430849561988587, 32'sd-0.0047645567444765625, 32'sd-0.05998924314824713, 32'sd-0.055504707038794926, 32'sd0.03092953662402751, 32'sd0.027924874416343785, 32'sd4.900743213539957e-124, 32'sd1.1296867009266272e-119, 32'sd-1.0381969020431222e-121, 32'sd5.663606372852779e-124, 32'sd0.07063947084962707, 32'sd-0.0101120685183947, 32'sd0.08579709600896676, 32'sd0.15758942632230563, 32'sd-0.10090060524203197, 32'sd-0.0741722021817881, 32'sd-0.1249817349500322, 32'sd0.020384586594091553, 32'sd-0.0919378247432089, 32'sd0.058133814897620234, 32'sd-0.14051005959228274, 32'sd-0.08705006303606157, 32'sd-0.04214949416205347, 32'sd0.07486750047532427, 32'sd-0.057516445154054414, 32'sd-0.11041569431678064, 32'sd0.03559976892451719, 32'sd-0.03977324456907036, 32'sd0.013767698396172662, 32'sd0.0039726680909678075, 32'sd0.025141271014966878, 32'sd0.030401725132676423, 32'sd0.08148445930663248, 32'sd5.784586811995034e-117, 32'sd1.480482366828581e-124, 32'sd-3.739510496143063e-119, 32'sd8.059168359563248e-125, 32'sd3.9679901297567233e-119, 32'sd-3.8505744631825716e-117, 32'sd0.02775569472680228, 32'sd-0.013802758714465183, 32'sd0.04217324899219098, 32'sd0.08491170228916547, 32'sd0.011599259961191318, 32'sd0.08374446279115076, 32'sd0.008740672754327484, 32'sd-0.019170038964611585, 32'sd-0.05289925529912641, 32'sd0.06308162630096767, 32'sd0.0412229782307643, 32'sd0.07704118139875618, 32'sd-0.06639428564531302, 32'sd0.0819046964341606, 32'sd-0.03834105938740788, 32'sd0.03199855385189388, 32'sd0.025254127094971802, 32'sd0.09424221007101452, 32'sd0.00648010682644269, 32'sd-0.005617988920404663, 32'sd-2.885996431365976e-125, 32'sd-3.3041652192121506e-115, 32'sd-2.059074326225528e-118, 32'sd1.0162531394426584e-124},
        '{32'sd3.1309981839676158e-114, 32'sd-1.7391328743758287e-125, 32'sd2.458428677924629e-124, 32'sd3.373093679496209e-126, 32'sd-6.89212231957709e-126, 32'sd-3.950676131580129e-119, 32'sd-1.526351847291776e-125, 32'sd1.0185242060129337e-127, 32'sd-3.2206470515148654e-114, 32'sd3.8006074495471885e-122, 32'sd-4.1708144878078645e-123, 32'sd-5.274292310724582e-127, 32'sd0.09465164778468367, 32'sd0.025712581907833036, 32'sd0.126134770507576, 32'sd0.13295993347144558, 32'sd2.5018520257232458e-114, 32'sd1.3965705674860773e-118, 32'sd-1.754642863865154e-117, 32'sd-4.4014156959500594e-123, 32'sd1.4902221565256056e-124, 32'sd3.090092317057109e-121, 32'sd2.6395867686109835e-125, 32'sd5.7434626977383924e-120, 32'sd4.947524770510739e-126, 32'sd-3.3115683534035056e-121, 32'sd7.925872899154436e-125, 32'sd-1.805215978308046e-123, 32'sd-4.341026724859704e-128, 32'sd-2.5579955977911527e-124, 32'sd-3.523012010868994e-128, 32'sd3.2794309515502193e-119, 32'sd-0.0305141669219792, 32'sd0.0047063414372331535, 32'sd-0.016154749935181657, 32'sd0.0812788874690666, 32'sd0.10232931067446867, 32'sd0.010694744192561924, 32'sd-0.0007061441156589184, 32'sd0.03947043478172505, 32'sd-0.0013051649710915207, 32'sd-0.061376035492205924, 32'sd-0.030671186706027264, 32'sd0.0790907073014481, 32'sd0.05252271973161158, 32'sd0.039119459277222546, 32'sd-0.02018252991725711, 32'sd0.00807866492159943, 32'sd0.03245418308078425, 32'sd-0.0239021529087794, 32'sd0.01665772881574959, 32'sd0.06030225883790559, 32'sd-7.629027601986107e-117, 32'sd4.551193867941101e-123, 32'sd3.334009255714322e-121, 32'sd-1.341732134235035e-122, 32'sd-2.9015291039051656e-120, 32'sd-2.859824645597968e-125, 32'sd0.10882698270452121, 32'sd0.03736082990165074, 32'sd0.0040604715027682476, 32'sd0.047174093481503705, 32'sd0.08690122288794054, 32'sd-0.054861381303446845, 32'sd-0.032344118129788206, 32'sd0.08743729195060165, 32'sd0.018458144030768744, 32'sd-0.03682436895646036, 32'sd-0.026437585592461517, 32'sd-0.0613936836943298, 32'sd-0.00128897144331603, 32'sd-0.0432376062315462, 32'sd0.053783426215151725, 32'sd0.03218095915497939, 32'sd0.003391108329157719, 32'sd0.09119389497798243, 32'sd0.027361795205059082, 32'sd-0.03984358710126238, 32'sd-0.05000356544184883, 32'sd0.02512647624508379, 32'sd-0.004693225076024335, 32'sd0.06581705097569322, 32'sd-3.0508244589837325e-119, 32'sd-2.2947663717429436e-118, 32'sd4.265608926759956e-123, 32'sd1.3139390062738078e-120, 32'sd0.008626746584619512, 32'sd-0.03294351469594444, 32'sd-0.07772896924441922, 32'sd-0.008171220384366185, 32'sd-0.010223434090273615, 32'sd-0.02461228916999472, 32'sd-0.04538286294598194, 32'sd-0.09206761488060299, 32'sd0.13815877891290954, 32'sd-0.06544128909975111, 32'sd-0.07683800626504855, 32'sd-0.06924523221664564, 32'sd-0.0440664593681276, 32'sd0.026734971644436962, 32'sd0.07516721737865079, 32'sd0.10518640525695663, 32'sd-0.035550363721935506, 32'sd0.026736150423824226, 32'sd0.06894691725019815, 32'sd-0.08208147052208492, 32'sd-0.06857071260377585, 32'sd-0.016866706638851252, 32'sd-0.0974618464478927, 32'sd-0.10074591077851758, 32'sd0.01735225258415672, 32'sd1.7394188766591802e-125, 32'sd1.1827430959908942e-117, 32'sd0.03916345151503948, 32'sd-0.010038425387195906, 32'sd0.05151657012532142, 32'sd-0.03704810968877774, 32'sd-0.11903317996820065, 32'sd-0.053866450004049514, 32'sd-0.13615996845738756, 32'sd-0.16700793722749396, 32'sd-0.11243219132594687, 32'sd0.017458155633532157, 32'sd0.06963431319965872, 32'sd-0.09757838322657678, 32'sd-0.06664210885661213, 32'sd-0.008421325147073664, 32'sd-0.01549757037023937, 32'sd0.09927786729361145, 32'sd0.17573163749276885, 32'sd0.03206148748483006, 32'sd0.15389188058171702, 32'sd0.06977511329176062, 32'sd-0.023595224857346952, 32'sd-0.0013940808242038623, 32'sd-0.0978772682105503, 32'sd-0.025438494122143634, 32'sd0.07803401831669118, 32'sd-0.09760180654272554, 32'sd0.01986674305234493, 32'sd4.312188884007981e-125, 32'sd0.06337735855239697, 32'sd0.026284108107306945, 32'sd0.04200768978792545, 32'sd-0.04240921102546991, 32'sd0.0301030243259322, 32'sd-0.01764848676466931, 32'sd-0.05830283510899757, 32'sd-0.03796851387357424, 32'sd-0.10560999215843174, 32'sd0.10859044855723748, 32'sd-0.02784350430587872, 32'sd0.036200961897812335, 32'sd-0.08457602025751948, 32'sd-0.16261981511395207, 32'sd-0.03729510614820775, 32'sd0.05708915038011633, 32'sd0.07446730046791339, 32'sd0.018600158807727467, 32'sd0.06355557829445985, 32'sd-0.06383985757581967, 32'sd-0.005176437038220669, 32'sd0.08990832340768605, 32'sd0.020424318902838613, 32'sd-0.16054043075490504, 32'sd0.0263199405305147, 32'sd-0.08507732312805806, 32'sd0.014496032572754303, 32'sd3.477770206470918e-122, 32'sd0.011495746753065137, 32'sd0.14368268576234347, 32'sd0.11693891032654076, 32'sd0.11550003688359349, 32'sd-0.0365058796947432, 32'sd-0.007762142908396158, 32'sd-0.016261922631171342, 32'sd0.04622791852683135, 32'sd0.052928810284077615, 32'sd0.24676955974884596, 32'sd0.17934790578505805, 32'sd0.10861255826124681, 32'sd-0.043124312715925074, 32'sd-0.05383415240955924, 32'sd0.05035445197620751, 32'sd-0.006638883509110983, 32'sd0.023651679429916084, 32'sd0.09330091347988474, 32'sd0.020347007729879962, 32'sd-0.04086056503608157, 32'sd0.05903318300511451, 32'sd0.08183514376632708, 32'sd-0.06241150581719143, 32'sd-0.0726747341990502, 32'sd0.04555391772020815, 32'sd-0.004312954272000709, 32'sd0.038630785238172316, 32'sd0.056080841828352934, 32'sd0.02351810452009532, 32'sd0.01017127518315892, 32'sd-0.0658726107195001, 32'sd0.03856465253085093, 32'sd0.014599220321677474, 32'sd0.08955258895771542, 32'sd0.1645851414750976, 32'sd0.14361553027056387, 32'sd-0.004175702047095202, 32'sd0.10057844464536718, 32'sd0.24717018197958396, 32'sd0.12011820554157274, 32'sd-0.12114937331532419, 32'sd-0.10543040266933101, 32'sd0.005973162557691311, 32'sd0.0539057830454942, 32'sd-0.021811084504791522, 32'sd0.047184844401616584, 32'sd0.16920580208906827, 32'sd0.07063960285883226, 32'sd-0.027114824062294443, 32'sd-0.07979985958377867, 32'sd0.07862956123646606, 32'sd0.13451494333664393, 32'sd0.06688881054548247, 32'sd0.06309193008280824, 32'sd0.003916082773916916, 32'sd0.04093237013804769, 32'sd0.004514366184856198, 32'sd0.059032269390440886, 32'sd0.011549735360057229, 32'sd0.02994456874215631, 32'sd-0.1039264153368006, 32'sd-0.08191155784117038, 32'sd0.06175544419246757, 32'sd0.06344803032597421, 32'sd0.04695573202600519, 32'sd-0.03276660467148033, 32'sd0.11285840429756164, 32'sd0.02746529699131986, 32'sd-0.012489840124908405, 32'sd-0.054563522827606445, 32'sd-0.04028766682856796, 32'sd-0.057693173961458614, 32'sd0.04395217707247568, 32'sd0.13347139941261024, 32'sd0.11254457491592422, 32'sd0.12826079600379972, 32'sd0.05403403020694042, 32'sd0.09881158459661771, 32'sd0.003662594945239605, 32'sd-0.008559436574775117, 32'sd0.07806811187293136, 32'sd-0.04045583248269922, 32'sd0.02057437779408666, 32'sd0.03733980850820103, 32'sd0.03650797860755126, 32'sd0.026878337476199173, 32'sd0.07911809723123958, 32'sd-0.009582452680755452, 32'sd-0.12562282184415302, 32'sd-0.14556078303698045, 32'sd-0.06529580371900154, 32'sd-0.1138706391767844, 32'sd-0.10632945294891373, 32'sd-0.08528254160637411, 32'sd-0.17151633324235596, 32'sd-0.1742774320769175, 32'sd-0.19622488186661832, 32'sd-0.16219758141366145, 32'sd-0.029931741638359138, 32'sd0.05963630392263305, 32'sd0.10860496497272248, 32'sd0.14770883154089282, 32'sd-0.0003328166963521274, 32'sd0.12238702836163931, 32'sd-0.013872086950012205, 32'sd6.981925915308051e-05, 32'sd0.026321373491142823, 32'sd-0.10378092910229779, 32'sd-0.09070156476011618, 32'sd-0.048406702220443, 32'sd-0.01773910810157062, 32'sd-0.012496591087411451, 32'sd0.019629590730295448, 32'sd0.08080400039192903, 32'sd0.11382930992041482, 32'sd0.016248771589029196, 32'sd0.02341304498078229, 32'sd-0.06562029535756264, 32'sd-0.21762476034321732, 32'sd-0.13802526666121986, 32'sd-0.22446410459192506, 32'sd-0.22388926208685442, 32'sd-0.23927143575610252, 32'sd-0.10216003591216335, 32'sd-0.1925225393355088, 32'sd-0.21397963435095307, 32'sd-0.030767466156813368, 32'sd0.04114127221819709, 32'sd0.031022934232833546, 32'sd0.05021132725649402, 32'sd-0.04083186023431, 32'sd0.12276953164120621, 32'sd0.11427078360735174, 32'sd0.09039565347486211, 32'sd0.006244830830795642, 32'sd-0.21074229664975525, 32'sd0.07090580134815053, 32'sd-0.010797853472336845, 32'sd-0.013552651498417558, 32'sd0.0007354857259816961, 32'sd0.09500201222189718, 32'sd0.06355034658964874, 32'sd0.02367151387060496, 32'sd-0.016906739020927715, 32'sd-0.14041592795820565, 32'sd-0.235225869967988, 32'sd-0.10775273140773813, 32'sd-0.19935537174255769, 32'sd-0.28820431732302065, 32'sd-0.25625676290787525, 32'sd-0.17563113392725138, 32'sd-0.12035026189583027, 32'sd0.03720877521727497, 32'sd-0.002380001132740576, 32'sd0.02715225809596079, 32'sd-0.12153167031698718, 32'sd-0.002630985290148806, 32'sd0.1268510324499888, 32'sd-0.07209982749942768, 32'sd-0.02382369354240016, 32'sd0.03970093676901648, 32'sd0.10273734269982883, 32'sd-0.041666183916668424, 32'sd-0.07254816662435455, 32'sd-0.1192458156645164, 32'sd0.006891208394691716, 32'sd0.0416146409027128, 32'sd0.08137035908952105, 32'sd-0.03289334029947425, 32'sd-0.0012833696226491012, 32'sd0.005254192198072679, 32'sd-0.03182304483021406, 32'sd0.008702758393912933, 32'sd-0.1531342131267318, 32'sd-0.1273562353769478, 32'sd-0.22255078108729331, 32'sd-0.2395406177807988, 32'sd-0.1008291659077752, 32'sd-0.003816046834803851, 32'sd0.0869576665513353, 32'sd0.06801988927892648, 32'sd0.004075066173608181, 32'sd-0.08863718039529757, 32'sd0.10074716215062754, 32'sd0.07760823381830334, 32'sd0.03835932551728082, 32'sd0.0051802537835547655, 32'sd0.04377018441276891, 32'sd-0.1105265079010279, 32'sd-0.021987052912463948, 32'sd-0.07321469061748277, 32'sd-0.014374909194018532, 32'sd-0.10334629888546068, 32'sd0.04425410896008913, 32'sd-0.01583078866120877, 32'sd0.0650465032922909, 32'sd-0.07735978256116872, 32'sd0.07529542807770784, 32'sd0.08734681849087428, 32'sd0.1060832430942492, 32'sd0.057580567887903056, 32'sd0.009717518963754657, 32'sd-0.05858231164940346, 32'sd-0.020285335482136714, 32'sd-0.061125939985758895, 32'sd0.03237996195107588, 32'sd0.07835992176245661, 32'sd0.021012336937027816, 32'sd-0.0013422772974555535, 32'sd-0.021020125818236864, 32'sd-0.11881549643433145, 32'sd-0.02378383006213258, 32'sd-0.01192443836445267, 32'sd0.04971010102391542, 32'sd-0.06352999420676214, 32'sd0.07802010989971501, 32'sd0.06331194202209997, 32'sd-0.01596796508353925, 32'sd0.04646462779860056, 32'sd0.026874105524159548, 32'sd0.04635128303512993, 32'sd0.05223634850193682, 32'sd0.05958233575856458, 32'sd0.08550066024948598, 32'sd0.0007159363735341215, 32'sd-0.03588395820113317, 32'sd-0.060753022282919865, 32'sd0.06387131694326205, 32'sd0.08327074063316818, 32'sd0.028610233819246562, 32'sd0.0387879058359528, 32'sd0.0727777852476075, 32'sd0.2016937731077168, 32'sd0.12616678817432586, 32'sd0.1475058715290435, 32'sd0.07950853668094224, 32'sd0.019264011528922074, 32'sd-0.09512511951590437, 32'sd-0.04116295042438108, 32'sd0.0489792112146053, 32'sd0.09275592471039423, 32'sd-0.013475927766430341, 32'sd-0.005934235709088773, 32'sd0.024571481598408204, 32'sd0.07004002047381057, 32'sd0.13451327250995967, 32'sd0.014305186125077087, 32'sd0.02410883533413178, 32'sd-0.013042763669007645, 32'sd0.04898882306492794, 32'sd-0.02318455556825231, 32'sd-0.08245459129410933, 32'sd-0.04524289631139207, 32'sd-0.050567712243229174, 32'sd0.13657307092491378, 32'sd0.03322711382418356, 32'sd0.07930129870222401, 32'sd0.09328306804809901, 32'sd0.01835750217269949, 32'sd-0.023856362017780165, 32'sd0.16546555910218602, 32'sd0.093577510289652, 32'sd0.13055046244182425, 32'sd0.17631715334203388, 32'sd0.153632550883866, 32'sd-0.008186326255459227, 32'sd0.036529396830549635, 32'sd0.11672534476549702, 32'sd0.04808006619034632, 32'sd0.002672454436564554, 32'sd-0.08022298091130937, 32'sd0.039988218736446146, 32'sd0.11329862221132476, 32'sd0.04484945250005789, 32'sd0.006188401277813245, 32'sd0.034792882748057044, 32'sd-0.015343778801718158, 32'sd0.02145064037043815, 32'sd0.0011419442022729345, 32'sd0.041613912233495705, 32'sd0.057257577566627096, 32'sd0.042974385315292296, 32'sd0.0642989923847533, 32'sd0.032442324782562384, 32'sd0.11944595825001382, 32'sd0.10041667922636752, 32'sd0.008872291575249417, 32'sd0.06155362284906856, 32'sd0.16053369107873855, 32'sd0.1307146416635053, 32'sd0.11136529029757723, 32'sd0.16383108153173206, 32'sd0.17124985643750745, 32'sd0.09688039354329187, 32'sd0.00417826814605762, 32'sd-0.002031313508058378, 32'sd0.048725604220919955, 32'sd0.028627793393421815, 32'sd-0.0218942172585912, 32'sd-0.04729476931265202, 32'sd0.04447065611678672, 32'sd0.014613740711819695, 32'sd-0.014354899477298372, 32'sd0.004546675122784712, 32'sd-0.024657089228477445, 32'sd-0.01682814821511403, 32'sd0.03975823211428027, 32'sd-6.91063243476695e-124, 32'sd0.07507379530112206, 32'sd-0.006158141894590072, 32'sd-0.051410250163409665, 32'sd0.09297962507922644, 32'sd0.10356271544825438, 32'sd-0.1176918287655388, 32'sd-0.07445919566600623, 32'sd-0.059312736348431684, 32'sd-0.08298825532689164, 32'sd-0.10589629247640807, 32'sd-0.15093735123579297, 32'sd-0.05157975095235784, 32'sd0.050274295519710376, 32'sd-0.052942590419020004, 32'sd0.020947318771408655, 32'sd-0.08960251541464366, 32'sd-0.019034782412485938, 32'sd0.04333358339061978, 32'sd-0.04686297851173358, 32'sd-0.1435903079499192, 32'sd-0.12921216695811522, 32'sd-0.18953632315995333, 32'sd-0.026517266211956915, 32'sd-0.03955999702273774, 32'sd-0.06550480977005205, 32'sd-0.03945562137408874, 32'sd0.05121933927553633, 32'sd0.01420176264206659, 32'sd0.06454755249434817, 32'sd0.03358268935347588, 32'sd0.05664405462530715, 32'sd-0.029911768893832454, 32'sd-0.0899377335715254, 32'sd-0.18527075251772418, 32'sd-0.06882800547112129, 32'sd-0.046456965740304924, 32'sd-0.06765940410463137, 32'sd-0.2120873138871307, 32'sd-0.13649391666275373, 32'sd-0.33321486488522584, 32'sd-0.11646663673502906, 32'sd-0.10242163036656103, 32'sd-0.06836871170060649, 32'sd-0.017180150533619883, 32'sd-0.05362306908998953, 32'sd-0.053818697381312515, 32'sd-0.1414575119490939, 32'sd-0.1311448682675722, 32'sd-0.08480270126948938, 32'sd-0.11095408490352038, 32'sd0.01948144830958752, 32'sd-0.048634004004952915, 32'sd-0.07365432877820734, 32'sd-0.06388151862656005, 32'sd-0.009296505435989637, 32'sd0.06424389672513497, 32'sd0.04728955189229714, 32'sd0.04739129178864349, 32'sd-0.0072217122086292, 32'sd-0.1438837762553388, 32'sd-0.05191105592735081, 32'sd-0.04214792112173146, 32'sd-0.030430164327326956, 32'sd0.00451380322437006, 32'sd-0.04325553804916791, 32'sd-0.16013258168473143, 32'sd-0.1223631563649336, 32'sd-0.21579126347074531, 32'sd-0.03856128830379788, 32'sd0.009790691323234952, 32'sd0.05208177684846795, 32'sd0.02817104520811746, 32'sd-0.05733693163297939, 32'sd-0.07633618271425434, 32'sd-0.13860748251744018, 32'sd0.03353389126013305, 32'sd-0.07479745882382571, 32'sd-0.03507666072826912, 32'sd0.06601490852070477, 32'sd-0.07708157891284426, 32'sd-0.0071431049015567355, 32'sd0.006098187075320337, 32'sd0.04717525254378604, 32'sd-1.495757217269872e-126, 32'sd-0.08794347148253409, 32'sd0.0661215165702937, 32'sd0.012157630107895575, 32'sd0.06787269255182939, 32'sd-0.10406965062836276, 32'sd-0.032268703163950335, 32'sd-0.016981040031795163, 32'sd0.05328312496212171, 32'sd-0.07348309948998273, 32'sd-0.051750045751666404, 32'sd-0.049232737126020346, 32'sd-0.0538492393779933, 32'sd-0.0052484982656756055, 32'sd0.1400277858347688, 32'sd0.036053739371893975, 32'sd0.01418296299279027, 32'sd-0.006928779558993964, 32'sd0.04090672793909618, 32'sd-0.035058919960273154, 32'sd0.0007074215267360005, 32'sd-0.09165898242587632, 32'sd-0.05499169165885769, 32'sd-0.07743755795390893, 32'sd0.07329091294004869, 32'sd-0.00610745938959631, 32'sd-0.041094211526058924, 32'sd0.04732714812964934, 32'sd0.030779823885523847, 32'sd0.028346587433260247, 32'sd0.0010599306492242288, 32'sd0.12274536729787328, 32'sd0.041415592127465206, 32'sd-0.047536462831981666, 32'sd0.02299147087827043, 32'sd0.029250620662034123, 32'sd0.06429324391258445, 32'sd-0.05707836007730894, 32'sd-0.09558964263523823, 32'sd-0.05757138284242764, 32'sd-0.012441144929994898, 32'sd0.042402525999397304, 32'sd0.021139911078132848, 32'sd0.15244155938905865, 32'sd-0.015122727213033356, 32'sd-0.00338794519532266, 32'sd0.02066953667112407, 32'sd0.020613668349487177, 32'sd0.04649971529354584, 32'sd-0.04537537048963619, 32'sd-0.03240025769187015, 32'sd-0.053176670814243876, 32'sd0.16901000562367274, 32'sd0.15098010188155753, 32'sd-0.00580556552514772, 32'sd0.06512611911300893, 32'sd0.09542981071623272, 32'sd0.07216650924139799, 32'sd0.04522969245589467, 32'sd0.07652774599694073, 32'sd0.07078207458121777, 32'sd0.0986670848488438, 32'sd0.08017361086500956, 32'sd0.09344046600587068, 32'sd-0.08424744035830259, 32'sd-0.15448608591459015, 32'sd-0.11096371183205331, 32'sd-0.021258078747034354, 32'sd-0.09978040208002172, 32'sd0.09960422241203411, 32'sd0.0062915611888501215, 32'sd0.11689210673012958, 32'sd-0.008670678514688229, 32'sd0.019845080794749996, 32'sd0.054465715528680035, 32'sd0.004871513296292175, 32'sd-0.001025903910454619, 32'sd-0.14179847365522152, 32'sd-0.04860797130856274, 32'sd-0.02587076453810123, 32'sd-0.012362031652044424, 32'sd0.05796543771822036, 32'sd0.10182167885233899, 32'sd0.09655309084828136, 32'sd-3.615199727641262e-114, 32'sd0.08631977198548144, 32'sd0.04871452307184178, 32'sd-0.051566885410226235, 32'sd0.04220913817008437, 32'sd0.02275345945068113, 32'sd0.038982056880162666, 32'sd0.09467136936719496, 32'sd0.05911729248753576, 32'sd-0.041225628001846495, 32'sd-0.0034722487646617482, 32'sd0.00903296666206385, 32'sd-0.06424698359759555, 32'sd0.040190866843218195, 32'sd-0.03412160355945048, 32'sd0.0576569436963742, 32'sd-0.017981372010808645, 32'sd-0.10437472233610419, 32'sd-0.08413601798936501, 32'sd0.03470125267188644, 32'sd-0.011884749199631318, 32'sd-0.10410540021707658, 32'sd-0.011766475965358335, 32'sd0.03605856475296923, 32'sd0.0859493616068306, 32'sd-0.03635382750419965, 32'sd0.08897517737262417, 32'sd5.895326873000953e-116, 32'sd4.539524817113874e-117, 32'sd5.270704608029367e-118, 32'sd0.03176806796879246, 32'sd-0.006149072846365999, 32'sd0.04948042118176834, 32'sd-0.005636530342367905, 32'sd-0.05802161136873974, 32'sd-0.043394232395268566, 32'sd0.10379093384431427, 32'sd-0.06913162106504155, 32'sd-0.0927664083768898, 32'sd-0.05907164925956777, 32'sd-0.09168583426039552, 32'sd0.004405056122528673, 32'sd0.007739940775987701, 32'sd-0.08499896959206148, 32'sd0.05711950466220996, 32'sd0.015253794660452676, 32'sd0.021171331206521767, 32'sd-0.07864145505322816, 32'sd0.04664076087679054, 32'sd-0.0620432615891857, 32'sd0.05795221824777544, 32'sd0.07717767744232279, 32'sd0.07765235007267741, 32'sd0.10876946279471797, 32'sd0.051948722359967794, 32'sd1.3265303676528802e-127, 32'sd1.090974993259765e-121, 32'sd-2.2381577831286252e-116, 32'sd0.02158465235821856, 32'sd0.06812488106679558, 32'sd0.014689280328424505, 32'sd-0.05635610305609612, 32'sd-0.08227271425808348, 32'sd-0.004146980433743958, 32'sd-0.0384687301108282, 32'sd-0.07520767420888812, 32'sd0.03372440486868766, 32'sd-0.00950978093992386, 32'sd-0.023545182729236714, 32'sd0.052201956041857, 32'sd0.05967326620449193, 32'sd0.0314574266602558, 32'sd0.09788977930354142, 32'sd-0.02224147549890499, 32'sd0.0062297776431311505, 32'sd-0.05619200735464954, 32'sd-0.010460118428586511, 32'sd-0.026744554122483402, 32'sd-0.07220232402026458, 32'sd0.11463621082219681, 32'sd-0.029608473604162973, 32'sd0.031302322832667526, 32'sd0.09644938447190197, 32'sd-1.0464793238361953e-120, 32'sd1.3231460144028977e-124, 32'sd1.2621374708847647e-118, 32'sd-2.5629869280151582e-126, 32'sd0.08524633480784682, 32'sd0.06801589673942554, 32'sd0.027327221471805278, 32'sd0.047319947907433095, 32'sd-0.04814310432813665, 32'sd-0.06744789435510108, 32'sd-0.04938686311603057, 32'sd0.01577594007076897, 32'sd-0.16718179765681745, 32'sd-0.0721405287417263, 32'sd0.04588598028075692, 32'sd-0.07148062212173985, 32'sd0.03685815941808982, 32'sd0.08712951618771518, 32'sd0.058238031021756724, 32'sd0.02859665003313204, 32'sd-0.10279355000355245, 32'sd-0.055531909806906164, 32'sd-0.04979284136894243, 32'sd-0.04239209445659338, 32'sd-0.024296031678258893, 32'sd0.06327053410550323, 32'sd0.05293433064479936, 32'sd7.946716699100812e-127, 32'sd-9.666847953226871e-121, 32'sd-2.0602832211845497e-117, 32'sd3.279899536418858e-121, 32'sd3.276678906642396e-121, 32'sd2.282381956779831e-114, 32'sd0.048489746988489506, 32'sd0.04152198762118918, 32'sd0.013970913868754497, 32'sd0.031601975878899784, 32'sd0.06469340963335192, 32'sd0.03368361362629314, 32'sd0.0357443119581417, 32'sd0.008342172196323586, 32'sd0.05350939516713792, 32'sd0.007960439669300053, 32'sd-0.002768800730954759, 32'sd-0.08820139113387597, 32'sd-0.041697036556454285, 32'sd0.025580831420128, 32'sd-0.026299647091588853, 32'sd0.04414361102523675, 32'sd0.004067105594016192, 32'sd0.022808310233839658, 32'sd-0.03217643749109305, 32'sd0.08860762945212904, 32'sd4.34151893942575e-124, 32'sd-3.8018030168109983e-122, 32'sd-7.548312163041471e-115, 32'sd4.822831607733121e-115},
        '{32'sd-1.0787474858362034e-124, 32'sd-4.991043330488925e-118, 32'sd6.348443312405035e-124, 32'sd-4.557653910961269e-123, 32'sd-1.927375630063717e-117, 32'sd1.4966272069795542e-114, 32'sd1.0568774979981024e-117, 32'sd5.6732559174257745e-115, 32'sd-1.739261016620708e-125, 32'sd1.1526141292461528e-117, 32'sd2.0220100002131977e-127, 32'sd3.589673098411619e-121, 32'sd0.0031658476543910815, 32'sd0.01832442124782364, 32'sd0.09869060559199257, 32'sd-0.035921895346516325, 32'sd8.034086905283681e-121, 32'sd-2.6608744466542183e-121, 32'sd9.414846940590762e-119, 32'sd-2.080353855051339e-116, 32'sd3.6033462743368722e-118, 32'sd1.4160454223302885e-121, 32'sd-6.388222526653972e-123, 32'sd-5.0233335703594564e-126, 32'sd4.092003973636472e-125, 32'sd4.0545555525198075e-125, 32'sd-5.984617324071074e-126, 32'sd6.345712077403072e-117, 32'sd1.6312067138278624e-115, 32'sd4.164732951608714e-124, 32'sd-3.271583208708437e-116, 32'sd1.8744696086635725e-124, 32'sd-0.024305489037678155, 32'sd0.0001925289085519588, 32'sd0.08858292227949416, 32'sd-0.03768585314210431, 32'sd-0.01182402890024749, 32'sd0.054681561485811374, 32'sd0.11000983834086311, 32'sd0.05910453473411926, 32'sd0.05603316447959827, 32'sd-0.02194004280424344, 32'sd0.07802889619629864, 32'sd0.0482827124534221, 32'sd0.10521887605494389, 32'sd0.011405971053931128, 32'sd0.03441779296638897, 32'sd-0.027835002183432545, 32'sd0.03005299695196402, 32'sd0.050844316913306, 32'sd0.05785137499342535, 32'sd0.06068899043525758, 32'sd-1.1364460119187119e-119, 32'sd-1.0461507542589566e-124, 32'sd-2.1973802231722206e-119, 32'sd1.2110671348813383e-114, 32'sd-7.537377383575672e-121, 32'sd8.632994987552018e-127, 32'sd0.047050058057744606, 32'sd-0.03274111500309803, 32'sd0.02085449345040612, 32'sd0.06624905435020624, 32'sd0.09369175170296609, 32'sd0.059835581223989034, 32'sd-0.04364837297470871, 32'sd0.05601219140321098, 32'sd0.04312010644218578, 32'sd-0.05396071895945102, 32'sd-0.06661797952467569, 32'sd-0.01925719448124484, 32'sd-0.003411880918318252, 32'sd-0.006555933401508847, 32'sd0.040527353329358584, 32'sd-0.015262320372850961, 32'sd0.04660100781965706, 32'sd0.0984887760552745, 32'sd0.023150970131005554, 32'sd0.11728583591988041, 32'sd0.0676842436263079, 32'sd0.08532276165471658, 32'sd0.017258520264082682, 32'sd0.1474387972314221, 32'sd2.9461414984069896e-128, 32'sd1.1298942990143105e-123, 32'sd-7.288576641757816e-127, 32'sd8.901355900066886e-122, 32'sd0.009568465403889618, 32'sd-0.02393254034105485, 32'sd0.06666111808382554, 32'sd-0.1101240100995895, 32'sd-0.13069503064177165, 32'sd0.00397944323468568, 32'sd-0.08814746648378459, 32'sd-0.026155291165821326, 32'sd-0.07233706963063063, 32'sd0.02469072474746592, 32'sd-0.019465776169500907, 32'sd-0.07728306128433968, 32'sd-0.15674708216894073, 32'sd-0.045684445610921456, 32'sd-0.030302949919560347, 32'sd-0.0893045338695785, 32'sd-0.0273404398439594, 32'sd-0.028709070396817506, 32'sd-0.02759669845302288, 32'sd0.12662820892721252, 32'sd0.11691395650631965, 32'sd-0.06215170967706915, 32'sd0.013433620233840626, 32'sd0.029163811114739834, 32'sd0.053622665314151496, 32'sd7.740341183204293e-123, 32'sd-1.2786614054663016e-123, 32'sd0.04321843856812376, 32'sd0.003217045584173349, 32'sd0.01345676133174408, 32'sd-0.08183776314237765, 32'sd-0.03854859370168633, 32'sd-0.005174566667053329, 32'sd-0.04717128690399915, 32'sd-0.08557771611337242, 32'sd-0.04608624324817919, 32'sd-0.0013533212011222241, 32'sd-0.01958925757280768, 32'sd0.05619519427933952, 32'sd-0.002717824610887862, 32'sd0.0038433150875521547, 32'sd-0.06825700775564038, 32'sd0.0011133525910106813, 32'sd-0.03148018730664377, 32'sd-0.031828556519523495, 32'sd-0.11261637394257173, 32'sd0.010990734217587677, 32'sd0.04586622279483001, 32'sd-0.02854525680472771, 32'sd0.013217282321404462, 32'sd-0.14919869463967161, 32'sd0.009298802955970265, 32'sd0.01090533055174991, 32'sd0.03667428018788405, 32'sd4.657797128778753e-117, 32'sd0.10862394974413257, 32'sd0.0699989411682054, 32'sd0.08188803974682164, 32'sd0.01626082787881617, 32'sd-0.009489679652765863, 32'sd-0.07948537265695481, 32'sd-0.06009053101714511, 32'sd-0.049352771629048324, 32'sd-0.09101386807215318, 32'sd0.016688687629131466, 32'sd-0.02142347850129579, 32'sd-0.06233392406947048, 32'sd-0.08078155673708734, 32'sd-0.038761384865000956, 32'sd-0.06212441213896895, 32'sd0.0034814823615085784, 32'sd-0.07445575731465108, 32'sd-0.06952342990541585, 32'sd0.035302185973086375, 32'sd0.05310810115976856, 32'sd0.1464534739898987, 32'sd0.06765053878737927, 32'sd0.08186233997656701, 32'sd-0.013918651811165056, 32'sd0.029812718979985917, 32'sd-0.018029190106028527, 32'sd0.05189114201230949, 32'sd-1.190298047874619e-120, 32'sd0.0383092005637832, 32'sd-0.008552993452893764, 32'sd-0.02198036930230796, 32'sd0.030438296506625665, 32'sd-0.1164938105885338, 32'sd-0.05650373351650501, 32'sd-0.07518625191589678, 32'sd-0.049691973188407075, 32'sd0.05585150412543606, 32'sd-0.028432978040856028, 32'sd0.031603262086431425, 32'sd-0.06480981282276158, 32'sd0.03540901428777049, 32'sd0.11275248403291782, 32'sd0.04202647538384695, 32'sd0.05575212007869748, 32'sd0.029177405979585916, 32'sd0.05154015816034656, 32'sd0.020036347052811022, 32'sd-0.09262019027759454, 32'sd0.03730233479920832, 32'sd0.057076452343344825, 32'sd-0.03269710890608855, 32'sd-0.017192279741576853, 32'sd0.03529151977850567, 32'sd0.06915561717204652, 32'sd0.006935253211727601, 32'sd0.0997925931326706, 32'sd0.007781631232286134, 32'sd0.056411788587511044, 32'sd0.013293637982634008, 32'sd0.013124787359428592, 32'sd-0.07527777602689734, 32'sd-0.1736383589426946, 32'sd-0.09818564976487013, 32'sd0.012438709885787337, 32'sd-0.015991678367355027, 32'sd-0.10014752497509795, 32'sd0.008594618880774878, 32'sd-0.10155828214540683, 32'sd0.09281778653624263, 32'sd0.16155011353643398, 32'sd0.054285702286857265, 32'sd0.14992560095485694, 32'sd-0.037528161640013415, 32'sd-0.016249043329034697, 32'sd0.15915880028420637, 32'sd-0.024185903679776, 32'sd0.05021607036550391, 32'sd0.036871938979067494, 32'sd-0.11058807295689811, 32'sd-0.07757474291668005, 32'sd-0.03093055034786644, 32'sd0.01797478707316008, 32'sd0.04342406817488099, 32'sd0.04855603069179818, 32'sd0.014375058650205346, 32'sd-0.06690289039848901, 32'sd0.06097031831112353, 32'sd-0.0562696490682417, 32'sd-0.07864283947601763, 32'sd-0.17036482364721298, 32'sd-0.0844318474594721, 32'sd-0.07139501429092061, 32'sd0.050884042208464306, 32'sd-0.04777748019419894, 32'sd0.0053167607243887, 32'sd-0.03332773343175673, 32'sd0.12522478408635154, 32'sd0.15966793737622792, 32'sd0.17533219255377738, 32'sd0.03671164830194666, 32'sd-0.030114837895821655, 32'sd-0.19165975010735506, 32'sd0.0173561850855113, 32'sd0.000380822503352739, 32'sd-0.002219353216454741, 32'sd-0.035275251183387875, 32'sd0.017905258887798377, 32'sd-0.05620523908536611, 32'sd-0.10117352890465352, 32'sd-0.04388507649259961, 32'sd-0.03048440650114919, 32'sd0.040596115795932, 32'sd-0.07213733184141244, 32'sd0.004322686033816265, 32'sd0.08904259805261701, 32'sd0.13689821028900584, 32'sd0.02995801626660511, 32'sd-0.09219044610839348, 32'sd0.05970611742872901, 32'sd-0.037043040280683816, 32'sd0.0764266483091458, 32'sd0.023332805249567292, 32'sd0.005493784965212603, 32'sd-0.019961375296670972, 32'sd0.1296213061225625, 32'sd0.18467786397960242, 32'sd0.17682822871499915, 32'sd0.02008168442461273, 32'sd-0.01288005634739056, 32'sd-0.032015895216352994, 32'sd-0.10601960637498002, 32'sd-0.028701923511065243, 32'sd-0.05049368113404171, 32'sd-0.028361977254205785, 32'sd-0.014742573669578415, 32'sd-0.01799604767516422, 32'sd0.032162743294649965, 32'sd0.02494914766893305, 32'sd-0.0047197861965569115, 32'sd-0.0019218085312155794, 32'sd0.07492512539414431, 32'sd0.012788808768551091, 32'sd-0.10730192855198863, 32'sd0.02755547793848646, 32'sd0.030871223513048437, 32'sd-0.0552631437422691, 32'sd-0.06887777696834074, 32'sd0.011204083026504856, 32'sd-0.03510213973110784, 32'sd-0.0051901950437162865, 32'sd-0.009918074778338897, 32'sd-0.0027919440243965553, 32'sd0.08477048478152201, 32'sd0.10993150724440681, 32'sd0.02504374314551277, 32'sd-0.03018301633867168, 32'sd-0.05505265375694544, 32'sd-0.11820697857443183, 32'sd-0.0014188453142622945, 32'sd-0.07688103183718564, 32'sd-0.044555101150018005, 32'sd-0.029717914098155482, 32'sd0.050650207259416075, 32'sd0.04078426928795271, 32'sd-0.0009122590398416011, 32'sd-0.0518771119688869, 32'sd-0.027429538368222924, 32'sd0.04028610561678516, 32'sd0.06164180041919881, 32'sd0.029027972186995335, 32'sd-0.03367987958322596, 32'sd-0.009246592923525457, 32'sd-0.10554532635178895, 32'sd-0.06904891041102558, 32'sd-0.07262143642240114, 32'sd-0.03384188447801552, 32'sd-0.056251562744667506, 32'sd0.040852628634333275, 32'sd0.008257128548065826, 32'sd-0.15599752372897174, 32'sd-0.1818376863989371, 32'sd0.04727070432745822, 32'sd0.0033594428702859503, 32'sd-0.05268065352006153, 32'sd-0.23748485185393736, 32'sd-0.15111514675015023, 32'sd0.018905938567561755, 32'sd0.005996215202645893, 32'sd-0.054305876546656286, 32'sd0.08754360263589128, 32'sd0.1290557001826627, 32'sd-0.029260232158822935, 32'sd-0.0264059513592507, 32'sd-0.03725030147925096, 32'sd-0.0021409861215133845, 32'sd0.035782574554781454, 32'sd-0.057238946838093926, 32'sd-0.02220715736127421, 32'sd-0.11522145534781318, 32'sd-0.13583887670486358, 32'sd-0.11743943112506113, 32'sd-0.10270352841886117, 32'sd-0.11620185579601021, 32'sd-0.03204129361433931, 32'sd0.035713843492127535, 32'sd-0.0022163126787454043, 32'sd-0.2183569025080819, 32'sd-0.2631499671400478, 32'sd-0.20380254968780656, 32'sd0.024366197478786523, 32'sd-0.05217711139034934, 32'sd-0.11948787536322175, 32'sd-0.1648600603436855, 32'sd-0.11220146327075498, 32'sd-0.1545595018227264, 32'sd-0.004818863372265407, 32'sd0.007055490835851548, 32'sd0.09674326450541201, 32'sd0.07024119702934549, 32'sd-0.02388778039549338, 32'sd-0.08596645655763245, 32'sd0.0467409020628373, 32'sd-0.05935102500072456, 32'sd0.04299184558314292, 32'sd0.03797740632606329, 32'sd0.016416671113607374, 32'sd-0.11164097071609871, 32'sd-0.024027199461380832, 32'sd-0.13566951028279098, 32'sd-0.11554501968385068, 32'sd-0.06868364534456896, 32'sd-0.08183182800715473, 32'sd-0.11106207056911829, 32'sd-0.20309539160855958, 32'sd-0.2054460971222516, 32'sd-0.03893574190223452, 32'sd-0.05373611575619822, 32'sd0.09486937271150146, 32'sd-0.07421458257023895, 32'sd0.00738552827923082, 32'sd-0.1404984532727576, 32'sd-0.1198009031913764, 32'sd-0.041522111365920024, 32'sd-0.06618838451886712, 32'sd-0.08410641538639425, 32'sd0.023367047673478712, 32'sd0.0010995880174573688, 32'sd-0.0480012328525164, 32'sd0.0328905141172191, 32'sd0.09119754789910636, 32'sd0.081046071330156, 32'sd0.06545660494565637, 32'sd0.007681853315776365, 32'sd-0.030713750009751014, 32'sd0.04465275819357208, 32'sd-0.07489975128743064, 32'sd-0.05751189494333088, 32'sd-0.05423835504855088, 32'sd-0.08771297989980299, 32'sd-0.0728904858964999, 32'sd-0.10609223546758396, 32'sd-0.13233836852965186, 32'sd-0.07045524904218135, 32'sd0.0037286603296954835, 32'sd0.038626065559296936, 32'sd0.22561901318607083, 32'sd0.0432226277935591, 32'sd-0.0046225363266742285, 32'sd-0.13323821808264666, 32'sd-0.12220506316732975, 32'sd-0.14570059835411922, 32'sd-0.20896701315997948, 32'sd-0.12246493188634015, 32'sd-0.11950209015796069, 32'sd0.0044974552892265195, 32'sd0.08408356494126812, 32'sd0.048383222247296506, 32'sd0.04172051480406331, 32'sd0.11661830133341067, 32'sd-0.03710697674526825, 32'sd0.0816289641183884, 32'sd0.01699837699129614, 32'sd0.0007737296463883914, 32'sd-0.025715459708836867, 32'sd-0.029127461379831826, 32'sd-0.03216685956866368, 32'sd-0.08631287329611986, 32'sd-0.07747966728918738, 32'sd0.02163856505523513, 32'sd0.15013512819656885, 32'sd0.12220550815454431, 32'sd0.2078517040589079, 32'sd0.3022526579226463, 32'sd0.047969964489602446, 32'sd-0.010577874819229437, 32'sd-0.06381730862821612, 32'sd-0.1250293049791445, 32'sd-0.06388932547302935, 32'sd-0.15705487917196584, 32'sd-0.1310277258923687, 32'sd-0.10840116924193179, 32'sd-0.1907038668813033, 32'sd-0.1641360233704751, 32'sd-0.11182008169474504, 32'sd-0.06308931178057885, 32'sd0.040756313214644915, 32'sd0.012661286304266195, 32'sd0.006129216991428612, 32'sd0.06274525494766854, 32'sd-0.07071960976474861, 32'sd-0.06310572970681572, 32'sd0.021608836866222607, 32'sd-0.06632677619541841, 32'sd0.10490813965453258, 32'sd-0.04240222120428776, 32'sd-0.04896073749528888, 32'sd0.30485559933642575, 32'sd0.3053449413338614, 32'sd0.11398198565955182, 32'sd0.10545890641814912, 32'sd0.12022982028118592, 32'sd0.13669186167215103, 32'sd-0.006614620622045564, 32'sd-0.06898508047999613, 32'sd-0.1510734628640592, 32'sd-0.09254611618392793, 32'sd-0.19699781400196845, 32'sd-0.17093585225108412, 32'sd-0.025342599065905882, 32'sd-0.04027110585633599, 32'sd-0.020595285717070824, 32'sd-0.03748420205293232, 32'sd0.04180635719960265, 32'sd0.03511819039246537, 32'sd0.023648135925105614, 32'sd2.2896599302081607e-118, 32'sd-0.05381509817125083, 32'sd-0.010912809193479998, 32'sd-0.012311319309157936, 32'sd0.015687596247481665, 32'sd-0.008414024605882822, 32'sd0.12367902754370658, 32'sd0.08599291321896843, 32'sd0.1489845397497956, 32'sd0.05357561227189948, 32'sd0.08679676749615138, 32'sd0.07034923709525932, 32'sd0.07588676817199337, 32'sd0.11495562433536528, 32'sd0.1489222731463128, 32'sd-0.04227831264966416, 32'sd-0.06305232181380914, 32'sd-0.005938289024147392, 32'sd-0.02272861326310103, 32'sd-0.03885975257483002, 32'sd-0.08039667470368436, 32'sd0.08974831870216067, 32'sd-0.04255961500160817, 32'sd-0.036526937163240424, 32'sd-0.09328384888583903, 32'sd0.01391589993932163, 32'sd0.11662279460534264, 32'sd0.045175583408654886, 32'sd0.012308341790556721, 32'sd0.09354592542662458, 32'sd0.017139688311004677, 32'sd-0.052253245108965854, 32'sd-0.007333719451534343, 32'sd0.09960791697977978, 32'sd0.057172986144768234, 32'sd0.12027544201767731, 32'sd0.03933055646252702, 32'sd0.016779325037011877, 32'sd0.09745010763731236, 32'sd-0.047451243982955124, 32'sd0.03207007672608384, 32'sd0.10998323330123516, 32'sd0.02152200557166223, 32'sd-0.09180578210403889, 32'sd-0.1184664321992117, 32'sd0.06058382706614012, 32'sd0.15049747965329538, 32'sd0.13552688594301546, 32'sd0.11839986559354952, 32'sd0.13545576190779873, 32'sd-0.03965303019377538, 32'sd0.0490986764030791, 32'sd-0.033667391940625714, 32'sd0.050077518626832386, 32'sd-0.03490600461346125, 32'sd0.05476594806455962, 32'sd0.07653066950910437, 32'sd0.04576015026946771, 32'sd0.054398701336715656, 32'sd-0.05577030468186418, 32'sd0.11203408020683052, 32'sd-0.012370792330280572, 32'sd0.12055494864512732, 32'sd0.11740960365490752, 32'sd0.13184581727264524, 32'sd0.07329301474289181, 32'sd-0.0022989671683046747, 32'sd0.08820850582412078, 32'sd0.04459371256132583, 32'sd0.053407674064447304, 32'sd-0.0047231447317968665, 32'sd0.02899192243071202, 32'sd0.034800394651662174, 32'sd0.10113148585560557, 32'sd0.12607222796411885, 32'sd0.14105642468565782, 32'sd0.09746423008911334, 32'sd0.09618448106364726, 32'sd0.08458133957384432, 32'sd0.10436190990635041, 32'sd-0.10313892118918007, 32'sd0.09888043438917948, 32'sd0.03613554336424778, 32'sd0.13342054742191045, 32'sd1.9035191983539218e-116, 32'sd-0.008723967865559824, 32'sd-0.01687774770350568, 32'sd-0.05196728418050693, 32'sd0.03525238225105316, 32'sd0.06506948280170383, 32'sd0.18756254029068134, 32'sd0.14296375701393824, 32'sd0.06426763502152619, 32'sd-0.046927408195839355, 32'sd0.003031593077715121, 32'sd-0.06306598169875959, 32'sd-0.06849353923175173, 32'sd-0.09105949725206576, 32'sd-0.05318015692417723, 32'sd0.1457063946120901, 32'sd0.09235769471892012, 32'sd0.0699003284282906, 32'sd0.17919272187022728, 32'sd0.15043851510443654, 32'sd0.19610460972090651, 32'sd0.1806057912838189, 32'sd0.10810517513634946, 32'sd0.17027555784432716, 32'sd0.0173857629114697, 32'sd0.032548570062309164, 32'sd0.007232942243347605, 32'sd0.06580973805400393, 32'sd-0.038866880104818424, 32'sd-0.06367190454629247, 32'sd0.11421805738308315, 32'sd0.1053713549662398, 32'sd0.027316442495805483, 32'sd0.1027749594035861, 32'sd0.06437622252213847, 32'sd-0.05183672285235467, 32'sd0.008068483484734112, 32'sd0.01415241951494682, 32'sd-0.05468680913693913, 32'sd-0.0614554404107764, 32'sd0.05634442647608074, 32'sd-0.010204255304994025, 32'sd0.07752555152052037, 32'sd0.0361390445394012, 32'sd-0.040832295371599665, 32'sd0.11873512493069396, 32'sd0.052165974562925585, 32'sd0.13939227840149968, 32'sd0.11009834713820839, 32'sd0.1184045301063154, 32'sd0.05882576382765512, 32'sd0.002612051627959457, 32'sd0.061251274596665885, 32'sd-0.026929897092459756, 32'sd-0.021816817613984258, 32'sd0.013146779958943961, 32'sd0.024868811816939097, 32'sd-0.04021062198549292, 32'sd-0.010102866301453878, 32'sd0.05281462508817359, 32'sd0.02077548224161981, 32'sd0.11079950902529669, 32'sd0.10283815568835145, 32'sd0.11032993543287116, 32'sd-0.05013448890200442, 32'sd0.031965460183526674, 32'sd-0.04315124652199872, 32'sd0.0008802000131331228, 32'sd0.11142852558338599, 32'sd0.1284726414432169, 32'sd-0.0976182199464871, 32'sd-0.037591708319824946, 32'sd-0.06009945679319322, 32'sd-0.0921018712594334, 32'sd-0.01428459917716226, 32'sd0.04121261839109942, 32'sd0.1383000051873851, 32'sd0.006832034117939735, 32'sd0.056727402508944764, 32'sd0.13092452834336732, 32'sd0.030709021523478878, 32'sd-0.0013260943797477128, 32'sd0.03603637188142327, 32'sd-0.005246322038449075, 32'sd1.5262361012898784e-125, 32'sd0.10510260905356307, 32'sd0.04716892587040597, 32'sd-0.0579050108713574, 32'sd0.03614516137618071, 32'sd-0.06150279541793455, 32'sd0.08177934269980704, 32'sd-0.0515440927735558, 32'sd-0.013261172954991489, 32'sd-0.09199545713049638, 32'sd0.011467400154285238, 32'sd-0.03036659487279869, 32'sd0.09961366449247593, 32'sd-0.03696403380748789, 32'sd-0.09280616310045615, 32'sd0.05646207152508117, 32'sd0.02782201071978921, 32'sd0.014783117853774118, 32'sd-0.021013113800412885, 32'sd-0.05741531471292723, 32'sd-0.02342471105387571, 32'sd0.043625546357504257, 32'sd0.06252333070498019, 32'sd0.09767780430032828, 32'sd-0.011175647054513028, 32'sd0.04060240058290309, 32'sd0.08394448173168778, 32'sd8.600703331919523e-117, 32'sd1.9203361017580123e-117, 32'sd-2.063522760644314e-127, 32'sd-0.06246984172968619, 32'sd0.033386610445381125, 32'sd0.10874794317534527, 32'sd0.04038264032192631, 32'sd-0.06038301841026148, 32'sd-0.04645392854069105, 32'sd0.0033615874888999714, 32'sd-0.07093477306903109, 32'sd-0.19253558499781934, 32'sd-0.16726060251269817, 32'sd-0.15101000192701824, 32'sd-0.06785107842993778, 32'sd-0.12488005187646767, 32'sd-0.21123834195510943, 32'sd-0.11605089610333082, 32'sd-0.09038771516943779, 32'sd-0.15836685332874526, 32'sd-0.16312795463460694, 32'sd-0.1227015029686081, 32'sd-0.0752236873659983, 32'sd0.05339959133260614, 32'sd0.020534928698763968, 32'sd-0.03562483587407188, 32'sd-0.0030960608697828233, 32'sd0.03012880345154949, 32'sd-1.9100090496990342e-121, 32'sd7.800940631040997e-126, 32'sd-2.488634603247927e-126, 32'sd0.06111351261244025, 32'sd0.06121562791301673, 32'sd0.024026870819272128, 32'sd-0.03131631114678014, 32'sd-0.044277001506512495, 32'sd-0.04578038505787645, 32'sd-0.009700525647350612, 32'sd-0.16887933643404596, 32'sd-0.22626159171914886, 32'sd0.0021736634547991165, 32'sd-0.06295436468304409, 32'sd-0.006921068108383442, 32'sd0.009059680759023941, 32'sd-0.03636427953544957, 32'sd-0.0247828614853689, 32'sd0.033523844706902076, 32'sd0.039033353718343905, 32'sd-0.05562505856661314, 32'sd-0.13953879799460356, 32'sd-0.014372589556714378, 32'sd0.020361047454938216, 32'sd-0.05023861278248324, 32'sd-0.0060998943530656624, 32'sd0.07604013387084263, 32'sd0.05568664589107617, 32'sd-3.415961484110646e-116, 32'sd3.583825966852851e-116, 32'sd-1.9289445710858783e-117, 32'sd2.7605037089878606e-123, 32'sd0.09855713271558514, 32'sd0.036496087498023196, 32'sd-0.015284474081612083, 32'sd0.011180541608980441, 32'sd0.0607299259590842, 32'sd-0.054483324668089264, 32'sd-0.0268828973027413, 32'sd-0.008059203841652979, 32'sd0.04150495322817852, 32'sd0.022244899827613875, 32'sd0.009072918132103069, 32'sd-0.029633758258641795, 32'sd-0.03090346121053856, 32'sd-0.11860882679776373, 32'sd-0.004120644167953084, 32'sd-0.008573855797671942, 32'sd0.01913507528699331, 32'sd-0.07197257168323636, 32'sd0.04286857406111308, 32'sd-0.05623576946729029, 32'sd-0.08748851368756304, 32'sd0.007830429403723676, 32'sd0.06257739595622665, 32'sd1.1534507798436736e-123, 32'sd1.3741595836365531e-125, 32'sd3.2204629242756716e-118, 32'sd3.605133116338163e-119, 32'sd3.5587781027635145e-122, 32'sd3.1667335470502956e-121, 32'sd0.06284096662010971, 32'sd0.06818766104659298, 32'sd0.02144721240978771, 32'sd0.06833169052191586, 32'sd-0.07981188062277578, 32'sd0.024224927297955046, 32'sd0.10407131626153542, 32'sd0.09969708391517186, 32'sd0.04754203964197386, 32'sd0.09894310376443781, 32'sd0.07242211229098831, 32'sd-0.018490721723781717, 32'sd0.07553720574448249, 32'sd0.011458859366209278, 32'sd-0.007437537977211441, 32'sd0.12767303867090637, 32'sd0.2171312586579731, 32'sd-0.023267564965632204, 32'sd-0.046064390080636626, 32'sd0.025932393176309635, 32'sd-3.9644827341654045e-115, 32'sd1.1294671523785113e-125, 32'sd-1.3794885516500135e-124, 32'sd-3.816002391703948e-118},
        '{32'sd-1.5178768073352874e-123, 32'sd-2.1378811951778075e-121, 32'sd-3.0977863968103187e-120, 32'sd2.6079740087146295e-126, 32'sd1.3392523506401807e-122, 32'sd-6.316033573235422e-115, 32'sd-3.466034587292866e-116, 32'sd4.8744768243584486e-123, 32'sd-1.340931525617781e-122, 32'sd8.138281223725472e-125, 32'sd6.879198020577529e-124, 32'sd-1.1099683823212323e-121, 32'sd-0.033068168165555856, 32'sd0.016548045821757392, 32'sd-0.044398796854716496, 32'sd0.06189536762535148, 32'sd1.2034282786320303e-123, 32'sd7.004914264049242e-127, 32'sd-4.990611650806373e-128, 32'sd3.757435817822057e-119, 32'sd3.6736661171663704e-123, 32'sd-3.669029146266369e-120, 32'sd-5.506705166380734e-127, 32'sd1.4864302561647057e-123, 32'sd-1.6073136392602997e-120, 32'sd-9.122040009486083e-121, 32'sd1.2767256571137657e-125, 32'sd-3.4424351368275164e-123, 32'sd1.6569408668634544e-127, 32'sd-6.002838505899082e-119, 32'sd1.958458086017528e-126, 32'sd6.602913704501861e-122, 32'sd0.0033608172762250844, 32'sd-0.04016713950531422, 32'sd-0.06653909354861647, 32'sd-0.01387806108209705, 32'sd-0.019753730351546702, 32'sd-0.044524963292311356, 32'sd0.03591841370588288, 32'sd-0.07595796796718751, 32'sd-0.011432011728552634, 32'sd-0.014839360686215693, 32'sd0.007981666428739355, 32'sd-0.012034143931849086, 32'sd0.06529542937361364, 32'sd0.08447895523694386, 32'sd0.07634208106825248, 32'sd0.06118512514817555, 32'sd-0.013874768591082137, 32'sd0.07239132371447962, 32'sd-0.002759522235280604, 32'sd-0.005664309338834809, 32'sd-1.2369667991109003e-127, 32'sd-1.8663192230251227e-121, 32'sd-1.292413125157501e-124, 32'sd-8.284382833238004e-122, 32'sd2.7517100914232163e-116, 32'sd-4.001375300756161e-125, 32'sd-0.009003768283849209, 32'sd0.009362581818375711, 32'sd0.0409725848127735, 32'sd0.10587227079829362, 32'sd0.04271567166935486, 32'sd-0.04592283538963697, 32'sd0.03761068538059449, 32'sd-0.06684936625595618, 32'sd0.0056803013855785236, 32'sd0.029468953210900255, 32'sd0.015262607599792605, 32'sd-0.11583717798755384, 32'sd-0.10357985084916312, 32'sd-0.06800443059964618, 32'sd-0.09562722521358262, 32'sd-0.005169447124690036, 32'sd0.010053205900248507, 32'sd-0.03903499686909529, 32'sd0.015925698942379066, 32'sd0.04104165327552266, 32'sd-0.012272800800141374, 32'sd0.015900617901776888, 32'sd0.024861696050570817, 32'sd-0.02134764027716197, 32'sd-6.582317065185851e-121, 32'sd-4.240741281804781e-121, 32'sd-2.370367405493154e-119, 32'sd2.5907786933105206e-124, 32'sd0.015811322948425383, 32'sd-0.04265780348243704, 32'sd0.0011229220768290385, 32'sd0.07031464516633293, 32'sd0.0320769912056303, 32'sd-0.035491915709784196, 32'sd-0.03211829245891734, 32'sd0.12986966574283001, 32'sd0.09198019417103538, 32'sd0.013283730903865294, 32'sd-0.05424644512044304, 32'sd0.0360921808277011, 32'sd0.0077214636857707705, 32'sd-0.0065849000339122, 32'sd-0.09024940314011087, 32'sd0.022028575870997085, 32'sd0.07809321042365516, 32'sd0.04017513107170683, 32'sd0.012745953846928844, 32'sd0.04039090043338343, 32'sd-0.04041919106921815, 32'sd0.06344832083771196, 32'sd0.035351792320390256, 32'sd0.06927870668246569, 32'sd0.02739933706977485, 32'sd-1.9753257517173827e-124, 32'sd5.289819346202123e-124, 32'sd0.04144144619204843, 32'sd0.025674541368940162, 32'sd-0.05546127780851798, 32'sd-0.075159888791555, 32'sd-0.011067147452968985, 32'sd0.0686208493651446, 32'sd0.008425082693797676, 32'sd0.025371730928427465, 32'sd0.13745213342156887, 32'sd0.0843639190782282, 32'sd-0.00963964533837217, 32'sd-0.023680027806724704, 32'sd-0.10107877909070415, 32'sd-0.10517871405191703, 32'sd0.018247396805986346, 32'sd0.042744091979738275, 32'sd0.0028998575915269256, 32'sd0.08904302935780489, 32'sd-0.033610019335597485, 32'sd-0.0040296032349360295, 32'sd-0.02969406837305285, 32'sd-0.08461614511849652, 32'sd0.0433969190103322, 32'sd0.038293545634023436, 32'sd0.02528588519940645, 32'sd0.06662308884623203, 32'sd-0.01668349015271252, 32'sd-3.6765208145499274e-116, 32'sd0.015013795819063274, 32'sd0.02972491349715835, 32'sd-0.12504717791691586, 32'sd0.04011272495216022, 32'sd0.0622120552884915, 32'sd-0.030405068936049766, 32'sd0.06766092054194783, 32'sd0.08539271855479934, 32'sd0.05657888788391929, 32'sd-0.05453653250013999, 32'sd-0.0322705720311817, 32'sd-0.02497268391073235, 32'sd0.06429533350618379, 32'sd0.0799905246310094, 32'sd-0.07620742213424013, 32'sd-0.12555669486543325, 32'sd-0.08536233366963913, 32'sd-0.004152583200014159, 32'sd-0.04118784855936774, 32'sd0.03468616809412582, 32'sd0.0943181630085987, 32'sd-0.06063120663470649, 32'sd0.05443093939526729, 32'sd-0.014118290292056785, 32'sd-0.02272163187804056, 32'sd0.02313662860465617, 32'sd-0.0009802723595211055, 32'sd-2.214581954925015e-126, 32'sd0.022252938607947755, 32'sd-0.054994183857201916, 32'sd-0.08910049288544522, 32'sd0.0010959465862799337, 32'sd0.032592013698623544, 32'sd-0.021309193954367166, 32'sd-0.002048529231992537, 32'sd0.057163568540654144, 32'sd-0.0353053844320543, 32'sd0.14192087905626188, 32'sd0.04695328175454719, 32'sd0.1108048582821039, 32'sd0.0412530426453726, 32'sd0.04023530823513001, 32'sd0.11615196012696, 32'sd0.0245501233035229, 32'sd-0.08334503312672217, 32'sd0.06002501646451634, 32'sd0.07731547460215843, 32'sd-0.001532739220367147, 32'sd0.11756679587285174, 32'sd0.04688550968296259, 32'sd0.003332673637836164, 32'sd0.04294861067303056, 32'sd0.00435070939319273, 32'sd-0.0036668686851500367, 32'sd-0.03908429079194767, 32'sd0.023796869514582496, 32'sd0.06330573283720928, 32'sd0.013698172495965989, 32'sd-0.19377671823038062, 32'sd-0.09622552258869986, 32'sd-0.0767342123516426, 32'sd0.028522904413346185, 32'sd0.016768750328994768, 32'sd0.057257555950898466, 32'sd0.07188248763275862, 32'sd0.13882648265325748, 32'sd0.1799726370708734, 32'sd0.06848468423951894, 32'sd0.25876964899849164, 32'sd0.1509501682242481, 32'sd0.12203453979337843, 32'sd0.1175847673367353, 32'sd0.036681239488121575, 32'sd-0.050412451374047144, 32'sd-0.050505630783405385, 32'sd0.08535420015899285, 32'sd-0.04724415828462067, 32'sd-0.06999581280413972, 32'sd-0.13029530041972642, 32'sd-0.08497065277400644, 32'sd-0.04242114519811852, 32'sd0.0063987837752258045, 32'sd-0.010954590876293104, 32'sd0.04178180760589359, 32'sd-0.016765365366405667, 32'sd-0.07252348567370222, 32'sd-0.043848257295137284, 32'sd-0.1241321397859594, 32'sd-0.006427316721400621, 32'sd0.061296790404730746, 32'sd0.03273497380443722, 32'sd-0.027466828305968347, 32'sd0.09174311574558343, 32'sd0.21001293014932176, 32'sd0.10413230089380507, 32'sd0.17512626780395427, 32'sd0.19231689300785978, 32'sd0.16654863178920637, 32'sd0.07110654855227581, 32'sd0.062134161120014936, 32'sd-0.013765494203892812, 32'sd-0.0612668497444785, 32'sd-0.037778080530369094, 32'sd0.010440732455110402, 32'sd-0.1365917142365761, 32'sd-0.1560144560407629, 32'sd-0.1925864715318001, 32'sd-0.034920890365822924, 32'sd-0.08699763940068661, 32'sd-0.06048316749733237, 32'sd-0.0932268177372063, 32'sd0.013114038229522056, 32'sd-0.07443395805582653, 32'sd0.10933869318765048, 32'sd0.016767096773928843, 32'sd0.03827841998171231, 32'sd-0.0019860883670516057, 32'sd0.05735480022282714, 32'sd0.042123527635248625, 32'sd0.008834525086951829, 32'sd0.2048270804129457, 32'sd0.0075137006991788415, 32'sd-0.07352148626067063, 32'sd0.061392685740901, 32'sd0.04746240922887512, 32'sd0.01640674481375667, 32'sd-0.056898688421728176, 32'sd-0.04745229442852513, 32'sd-0.03883280256423609, 32'sd0.12284738208346424, 32'sd0.034336892708241445, 32'sd-0.03294346167095208, 32'sd-0.0005974703782005642, 32'sd-0.044835827938876964, 32'sd-0.10345700519687086, 32'sd0.02402998458423792, 32'sd-0.01713496455009498, 32'sd-0.09254241587507334, 32'sd0.07717093747310981, 32'sd0.01485211304305904, 32'sd-0.10410445266006361, 32'sd0.11679422365560195, 32'sd-0.07443901104665639, 32'sd0.018764661496054574, 32'sd0.04138586088654861, 32'sd0.11930117365454042, 32'sd0.006766487689553117, 32'sd0.0404897352489115, 32'sd0.05839423314055584, 32'sd0.0910174950174882, 32'sd0.016631452551062086, 32'sd-0.14576038719970244, 32'sd0.006739149468469857, 32'sd-0.07251315474348323, 32'sd-0.0394452589192282, 32'sd-0.03431914347991539, 32'sd0.10314011573462309, 32'sd0.11180228464115394, 32'sd-0.02374815280415378, 32'sd-0.07065544109869519, 32'sd0.017046928395396246, 32'sd0.07921549986535359, 32'sd-0.025315188599479507, 32'sd-0.07614675920380701, 32'sd-0.04496254384147138, 32'sd-0.025068685794700132, 32'sd0.0017206047910971417, 32'sd0.02116313791106585, 32'sd-0.0043489656390743306, 32'sd-0.020922749350870497, 32'sd-0.027573729763760754, 32'sd-0.0038021192918361404, 32'sd0.07730465987129075, 32'sd0.06193943182205904, 32'sd-0.04300871779035596, 32'sd0.06490044530504484, 32'sd0.06457466479168943, 32'sd0.018636176687631466, 32'sd-0.006890683301833648, 32'sd-0.17817730813337396, 32'sd-0.17816279781865837, 32'sd-0.21801825632242047, 32'sd-0.10100166881732937, 32'sd-0.01743403748739003, 32'sd-0.05872063869828262, 32'sd0.015769960745527615, 32'sd-0.0010673182040721607, 32'sd0.028739074406483572, 32'sd0.0899525061147623, 32'sd0.11906169491651232, 32'sd0.12723231737273166, 32'sd0.02876891470370917, 32'sd-0.09965003961419573, 32'sd0.03270900351317303, 32'sd0.0729840081041993, 32'sd0.01413487067685097, 32'sd0.08433768853994596, 32'sd-0.03175297780008741, 32'sd-0.049009735350274426, 32'sd0.04644713260512992, 32'sd-0.04260250699096458, 32'sd0.10675134410042704, 32'sd0.03550087079719999, 32'sd-0.05246290594113831, 32'sd-0.029726353227114814, 32'sd-0.05898566533004888, 32'sd-0.15541495985624754, 32'sd-0.180738525164037, 32'sd-0.08542707262351196, 32'sd-0.06800407219996737, 32'sd-0.0517223693855581, 32'sd0.03886926835800422, 32'sd-0.06903469014021069, 32'sd-0.014044863114175596, 32'sd-0.07433480958394668, 32'sd0.07644483860703898, 32'sd0.1279155104334011, 32'sd0.03431746148710896, 32'sd0.059565407514164, 32'sd-0.09627154813300419, 32'sd-0.04694116817396208, 32'sd0.03275128832444818, 32'sd-0.06408719956044989, 32'sd-0.00029162733290722634, 32'sd0.02255931811314969, 32'sd0.0591653711969866, 32'sd0.08202330446539594, 32'sd0.0711292634035389, 32'sd-0.055923152092755925, 32'sd0.05852699740226247, 32'sd0.04227126991890732, 32'sd-0.001463746600738053, 32'sd-0.06211589018625066, 32'sd-0.04187438825463089, 32'sd-0.14685753546006422, 32'sd-0.02535968394408119, 32'sd-0.09003648579534598, 32'sd-0.049321966066572444, 32'sd-0.15497525393942976, 32'sd-0.10690512133268074, 32'sd-0.1084682228345305, 32'sd-0.07929398444401828, 32'sd-0.024029093312947957, 32'sd0.11769737914665929, 32'sd-0.014907139905902665, 32'sd-0.017645042029415595, 32'sd-0.0765755610039675, 32'sd0.11545054162669009, 32'sd0.12585153443055905, 32'sd0.018887221422652672, 32'sd0.0626445819546467, 32'sd-0.006059648280550392, 32'sd0.04146272741101601, 32'sd0.07715823080818673, 32'sd0.06078855154259254, 32'sd-0.09176159188008032, 32'sd-0.1281590040284896, 32'sd-0.1094934748013952, 32'sd-0.06368718863473928, 32'sd0.026570402684071414, 32'sd-0.07063395500381092, 32'sd-0.01166458843476464, 32'sd-0.12746513556059152, 32'sd-0.07702112705575712, 32'sd-0.07684737209292386, 32'sd-0.1112799634726733, 32'sd-0.08506672372061809, 32'sd-0.21841634447519886, 32'sd-0.0936451435711234, 32'sd0.007099946597554834, 32'sd0.010888512471784876, 32'sd0.11818984694868394, 32'sd-0.039167994589036054, 32'sd-0.051293111764574684, 32'sd-0.013241516874000341, 32'sd0.06353154845208835, 32'sd-0.022167083232621274, 32'sd0.06921147079920609, 32'sd0.0014112148995980595, 32'sd-0.008568027137747482, 32'sd-0.007063817866827227, 32'sd0.051796767885550696, 32'sd-0.000395271959619603, 32'sd0.020563097480716074, 32'sd-0.007056763994553339, 32'sd-0.14194548350255623, 32'sd-0.11407763226555315, 32'sd-0.05301740182981891, 32'sd-0.06920129535409955, 32'sd0.045934607170155205, 32'sd0.04169769289482544, 32'sd0.02159354303871288, 32'sd0.010159473136340072, 32'sd-0.11313496891083713, 32'sd-0.05178474560018819, 32'sd-0.15689505564036366, 32'sd-0.10550635553756979, 32'sd0.08842933927504519, 32'sd-0.04899232261956373, 32'sd0.09369987391931768, 32'sd0.10743034207152963, 32'sd0.05427722091668981, 32'sd0.021984447650673512, 32'sd0.08002937890038732, 32'sd-0.10047331169957531, 32'sd0.08199963641996384, 32'sd0.011704714248678066, 32'sd0.01987289230510501, 32'sd0.08050286820954336, 32'sd-0.030587513978000927, 32'sd-0.06599990609467427, 32'sd0.02177935183848349, 32'sd0.03401789059603502, 32'sd0.003671617717784333, 32'sd0.0067665519199444635, 32'sd-0.06177764347560621, 32'sd-0.040860335229924535, 32'sd0.1423784925531855, 32'sd0.10021844280272382, 32'sd0.16925567865558613, 32'sd0.0899483466131496, 32'sd0.02619258425895483, 32'sd-0.13859247407895992, 32'sd-0.20319231878787522, 32'sd-0.06377775368144925, 32'sd-0.10382763658367171, 32'sd-0.0025207987659368633, 32'sd0.040389120547734435, 32'sd-0.017152226285457532, 32'sd-0.03153285249183669, 32'sd0.08461675451552249, 32'sd-0.05256877161589363, 32'sd0.007469322208341596, 32'sd0.002558426807339055, 32'sd-0.09282979238490907, 32'sd1.0492070093094069e-120, 32'sd-0.017503422710435604, 32'sd-0.06048794609581514, 32'sd0.007203323209732229, 32'sd0.0013823285874543288, 32'sd0.1098097045153161, 32'sd0.0210052439617703, 32'sd-0.010940604052716643, 32'sd-0.08432258688339934, 32'sd-0.007295532452794123, 32'sd0.011662124773386387, 32'sd-0.03114621753571337, 32'sd0.047410650729129145, 32'sd0.0747472428326604, 32'sd-0.08781616153329314, 32'sd-0.12762619068202535, 32'sd-0.0605887259448599, 32'sd-0.14828618212457673, 32'sd-0.09161604276632204, 32'sd0.057233409497389344, 32'sd0.06069802279881223, 32'sd-0.08929434643141103, 32'sd0.03716287099981945, 32'sd0.12081223139746865, 32'sd0.04450519569437616, 32'sd0.020246145495641753, 32'sd-0.06964049910505848, 32'sd0.07590616496216789, 32'sd0.010339437893017129, 32'sd-0.061991904199981754, 32'sd0.05001656866695072, 32'sd0.006663363820942026, 32'sd-0.10694858095069401, 32'sd0.020564782566781913, 32'sd0.0005457447200687516, 32'sd0.10110570640196677, 32'sd-0.03643129092974766, 32'sd-0.036153664887425815, 32'sd0.0013616034439555432, 32'sd-0.042317013044314795, 32'sd-0.06820667962913059, 32'sd-0.04304373465463462, 32'sd-0.20898431264137546, 32'sd-0.043930095386750065, 32'sd-0.01312665220102445, 32'sd-0.03065972374691959, 32'sd-0.04470850643757982, 32'sd0.08082630498423177, 32'sd0.06944839348219768, 32'sd-0.02620338098043525, 32'sd0.05535472484496991, 32'sd0.08617567368932423, 32'sd0.013086415324268538, 32'sd-0.019818011227379882, 32'sd-0.08537722686344074, 32'sd0.028360753193698587, 32'sd0.027821395058350237, 32'sd0.00851782125176765, 32'sd0.011099864046002073, 32'sd0.029179528159377355, 32'sd0.040836912303151764, 32'sd0.027436562638391414, 32'sd-0.027985573869819605, 32'sd-0.030626114416534813, 32'sd-0.09510499593666367, 32'sd-0.04577493584365506, 32'sd-0.04947854668037545, 32'sd-0.0492446153330383, 32'sd-0.11559938378898714, 32'sd-0.23387813489228854, 32'sd-0.22783637950808586, 32'sd-0.06557878759515898, 32'sd-0.005435693718976333, 32'sd0.05248571420601956, 32'sd0.06007600051932605, 32'sd0.002270224900186086, 32'sd0.11675017905412567, 32'sd-0.1073370066674691, 32'sd0.022143776172520727, 32'sd0.10026974029200796, 32'sd0.11957249832491057, 32'sd-0.10099681241145446, 32'sd-0.08189459753423425, 32'sd-0.0073251963611676236, 32'sd6.805479086925313e-115, 32'sd0.060009949629162465, 32'sd0.057787059804712035, 32'sd0.034317188412553455, 32'sd0.050070390594895604, 32'sd-0.024716276242013172, 32'sd-0.060875620554446556, 32'sd0.006968648064721775, 32'sd0.012761608678813239, 32'sd-0.03366612173694948, 32'sd-0.1761946621607936, 32'sd-0.21948215791435916, 32'sd-0.17639983813883556, 32'sd-0.14764527293053115, 32'sd5.5171197991108416e-05, 32'sd0.13405550637983243, 32'sd0.17363198208514183, 32'sd0.1249294730645542, 32'sd0.0908715965010053, 32'sd-0.011808275500899454, 32'sd0.0007219831153937534, 32'sd-0.027711063525586162, 32'sd-0.03786362414542953, 32'sd-0.006840090275404566, 32'sd-0.06420787438327094, 32'sd-0.007976954936038136, 32'sd-0.035529426758754964, 32'sd0.03710325632228137, 32'sd-0.00962270439707765, 32'sd-0.08761116333239347, 32'sd-0.04661777587024103, 32'sd0.11514886596742856, 32'sd0.03704367838510407, 32'sd-0.04292256001750736, 32'sd0.03088460798300616, 32'sd0.06220963638516899, 32'sd-0.10618334036015437, 32'sd-0.08746254018138953, 32'sd-0.07549165728610219, 32'sd-0.08228324897820673, 32'sd-0.10377939915097642, 32'sd-0.0418682796312621, 32'sd0.17566249522135685, 32'sd0.23879718193790078, 32'sd0.06524745334571273, 32'sd-0.059897545687294655, 32'sd-0.04674852210623209, 32'sd-0.06382827460659436, 32'sd-0.08329151757355534, 32'sd-0.1046028211198404, 32'sd-0.024884543755697493, 32'sd-0.1376502895907287, 32'sd-0.13847886638446547, 32'sd0.10245842037817539, 32'sd0.06383406951948334, 32'sd0.02510868668162369, 32'sd-0.018116691596190802, 32'sd-0.009475025156419795, 32'sd-0.08423948479148459, 32'sd0.03772381138220355, 32'sd0.10298142365710995, 32'sd0.048818934697830385, 32'sd-0.011082075653344129, 32'sd-0.06403479999066557, 32'sd-0.04719197671918362, 32'sd-0.019836475219384885, 32'sd-0.04631024892411761, 32'sd0.0495612971237488, 32'sd0.009560842713688874, 32'sd-0.043463090732259305, 32'sd0.11338899589139649, 32'sd0.08782547159640217, 32'sd0.05075015289065436, 32'sd0.05792515765273309, 32'sd0.08067827563335753, 32'sd0.05655343011676912, 32'sd0.000697835206898366, 32'sd-0.01813655306493757, 32'sd-0.009062462822008453, 32'sd0.0023379421236271866, 32'sd-0.04270123225868418, 32'sd0.03395048094364153, 32'sd0.08477682863277156, 32'sd0.008390262954717823, 32'sd2.030667044239116e-124, 32'sd0.04742515752924869, 32'sd-0.034871869650042644, 32'sd0.017994068101662052, 32'sd-0.07760571571030496, 32'sd-0.05416184064959452, 32'sd0.013371006229139887, 32'sd-0.08569968477031865, 32'sd-0.03970729342488254, 32'sd0.005167287863649379, 32'sd0.07679319248258162, 32'sd0.05177168664413764, 32'sd0.0026578492429788223, 32'sd0.04155747530465646, 32'sd0.13481965942557916, 32'sd0.16569834557294166, 32'sd0.03878578439844835, 32'sd0.06336898762630373, 32'sd-0.022698262976412364, 32'sd-0.0018396825036791089, 32'sd-0.08737357160363457, 32'sd-0.10388331658548648, 32'sd-0.0005750234531193076, 32'sd0.08538452571611846, 32'sd0.03557620267848065, 32'sd0.0705623829170492, 32'sd0.0843693986685697, 32'sd-3.452230334224206e-114, 32'sd5.781489109410655e-122, 32'sd-1.0640503482640003e-118, 32'sd-0.025811310117327364, 32'sd0.0582732460655082, 32'sd-0.04403394937187341, 32'sd0.06214993221496683, 32'sd-0.035683172670666466, 32'sd0.10985167326562867, 32'sd0.1410701937450518, 32'sd0.09391001868633643, 32'sd0.11951282902693375, 32'sd0.08311440186927384, 32'sd0.16066270142831168, 32'sd0.08336110799919796, 32'sd0.20302051074049798, 32'sd0.09632748846757705, 32'sd0.04643041797291894, 32'sd0.07390549805242723, 32'sd0.09654613227416577, 32'sd0.022897211644103972, 32'sd-0.009701256470911945, 32'sd0.044082267960640485, 32'sd0.10670743578594014, 32'sd-0.004323185651360133, 32'sd0.014515212296620353, 32'sd0.026069919852294357, 32'sd-0.017652929820253547, 32'sd-8.527798765157891e-126, 32'sd-1.2742798874917524e-123, 32'sd3.25334424190091e-116, 32'sd-0.006034315977053626, 32'sd0.02267467209632286, 32'sd-0.057871295449418686, 32'sd-0.0154525703786314, 32'sd0.021784932277930668, 32'sd0.1153623972784301, 32'sd0.1994824962409545, 32'sd0.1858868649798471, 32'sd0.1436602529186373, 32'sd0.028199249295832274, 32'sd0.1835968043132205, 32'sd-0.0900758141747048, 32'sd-0.09671094833354554, 32'sd0.0954758301724713, 32'sd0.002565150595170547, 32'sd-0.04569658042297193, 32'sd-0.026279562668801926, 32'sd0.07404044344152663, 32'sd0.055299310529687916, 32'sd0.02248220615852549, 32'sd0.0035862775695476544, 32'sd0.0067050170668125865, 32'sd0.09589325134544119, 32'sd-0.007663188940185745, 32'sd-0.005821414004428119, 32'sd-5.169774146545798e-124, 32'sd2.6125314836779587e-126, 32'sd6.947537895009206e-128, 32'sd5.3317009500862825e-126, 32'sd0.04763075658506265, 32'sd-0.09524822105950484, 32'sd0.024721094965937558, 32'sd-0.08854979315820254, 32'sd0.002621886321783535, 32'sd-0.11013832745434489, 32'sd-0.051546943867326486, 32'sd0.045278783893423546, 32'sd-0.05288197202413123, 32'sd-0.035565452433428936, 32'sd0.052421751387969256, 32'sd-0.009263579601306015, 32'sd0.14374559098397766, 32'sd0.07465243362907724, 32'sd-0.03750194583983784, 32'sd-0.08940942946248025, 32'sd0.04038845030122284, 32'sd0.08014071853549151, 32'sd0.01774315753520816, 32'sd-0.028962176827690096, 32'sd0.025523272039772612, 32'sd0.02882136048094237, 32'sd0.04283739530776438, 32'sd1.5139729806840634e-123, 32'sd-7.450429091496902e-120, 32'sd5.4060254358549e-118, 32'sd-6.83019914336332e-117, 32'sd-1.988407628997084e-122, 32'sd1.372580975828325e-118, 32'sd0.03163937267098909, 32'sd0.028852624765942733, 32'sd0.028707214440939398, 32'sd0.057424405970016204, 32'sd-0.02485756220510007, 32'sd-0.008522458246820476, 32'sd0.0508157587647369, 32'sd0.07371217919501846, 32'sd-0.03410659705264504, 32'sd-0.043626500330913545, 32'sd-0.01921401321195381, 32'sd0.074720213848956, 32'sd0.07106030277976093, 32'sd0.05710226812170862, 32'sd-0.013465827367799114, 32'sd-0.023335368844693713, 32'sd-0.09813556849183036, 32'sd-0.021607193990114133, 32'sd0.08603725891412425, 32'sd-0.06750969629853294, 32'sd2.0120253561174824e-116, 32'sd1.0529490495818088e-126, 32'sd1.8183971693955886e-123, 32'sd-1.425585004746485e-116},
        '{32'sd7.142720769103899e-127, 32'sd-9.034516059134743e-118, 32'sd4.8174828855154485e-127, 32'sd1.3097583277543491e-124, 32'sd-1.793670282541665e-127, 32'sd4.2193638276843066e-117, 32'sd-1.255629269625971e-114, 32'sd1.7486020728338108e-123, 32'sd1.462823884943185e-116, 32'sd7.046204648082457e-128, 32'sd3.653762634620115e-124, 32'sd2.2638770247400272e-125, 32'sd0.10484768973874938, 32'sd0.0001063821446069797, 32'sd-0.006816595482440789, 32'sd0.04501732324148441, 32'sd-1.165591039398861e-118, 32'sd-1.2984588859700957e-121, 32'sd1.959256395313932e-123, 32'sd-1.0716333529830035e-122, 32'sd-9.523554343963474e-126, 32'sd-2.0855534647703465e-118, 32'sd1.0281527270209524e-118, 32'sd-2.615927223118298e-125, 32'sd-5.5734647573462645e-121, 32'sd7.0045122568578266e-121, 32'sd-7.501802969606799e-117, 32'sd-3.8681622737255844e-125, 32'sd-1.4226496022423731e-118, 32'sd9.02334142278854e-118, 32'sd-3.959417219165844e-119, 32'sd1.9940078734285574e-119, 32'sd0.01918831012786197, 32'sd-0.040871029874419096, 32'sd-0.026358431271259822, 32'sd0.118497814288545, 32'sd0.0909693951261921, 32'sd0.024197303495181937, 32'sd0.061260938940780774, 32'sd-0.07541060202086153, 32'sd0.01757851484877479, 32'sd-0.024568261673293897, 32'sd-0.0819188511254019, 32'sd-0.010373818942796304, 32'sd0.0003758092390373839, 32'sd-0.014027789940988524, 32'sd0.12326579874991994, 32'sd0.07890750097294771, 32'sd0.005353742486549925, 32'sd0.11386103641706642, 32'sd0.0853599803380002, 32'sd0.08468114976101554, 32'sd-3.361654920446711e-120, 32'sd-6.835460579199347e-126, 32'sd-3.3375532563865543e-127, 32'sd-3.964232641672803e-119, 32'sd6.899601415834925e-117, 32'sd-9.80158633895866e-125, 32'sd0.044905166569646694, 32'sd0.014394754864396796, 32'sd0.055639831166671254, 32'sd0.02750559046065679, 32'sd-0.06334638257140592, 32'sd0.09684727370659936, 32'sd0.08420099660200833, 32'sd0.10983005570090458, 32'sd-0.06813483254951588, 32'sd-0.05107611791550138, 32'sd-0.04910812099924986, 32'sd-0.03362813808582836, 32'sd-0.02738415147967998, 32'sd0.1160053876789997, 32'sd0.06457989577877282, 32'sd0.09086164068413016, 32'sd-0.03610587110994457, 32'sd-0.010810832739020757, 32'sd0.04414967268622315, 32'sd0.08235114234084105, 32'sd-0.012343987010740212, 32'sd0.02951780698732566, 32'sd0.06833486072111285, 32'sd0.0969758264600428, 32'sd1.3352944568929978e-122, 32'sd-1.922136912706873e-117, 32'sd1.2128048309336601e-128, 32'sd-3.263413680335442e-122, 32'sd0.005039722212765642, 32'sd0.020977905058357248, 32'sd-0.0936870097714972, 32'sd-0.0040619553564083125, 32'sd0.018703931224487432, 32'sd-0.01790758702494109, 32'sd0.16688360761387228, 32'sd-0.07995483579212298, 32'sd-0.026262507624364672, 32'sd0.11537890603213555, 32'sd-0.028214404811818458, 32'sd0.04726635559491225, 32'sd0.0502933282843078, 32'sd-0.01603141871919944, 32'sd0.11896413629364598, 32'sd0.028080804978586466, 32'sd-0.05056070904785234, 32'sd-0.03859875560755701, 32'sd-0.12080967394037034, 32'sd-0.01777239534006019, 32'sd-0.0414549409888806, 32'sd0.038766830997769994, 32'sd0.01574850445512949, 32'sd0.026791580328933706, 32'sd0.014943606329903623, 32'sd2.2486575749364365e-126, 32'sd-3.3711702884526586e-120, 32'sd0.019036989484140423, 32'sd0.014699315718782411, 32'sd0.10719145088961458, 32'sd-0.08420775939766317, 32'sd-0.05001292473715054, 32'sd-0.002848983490491828, 32'sd0.04712848027533418, 32'sd0.10877378350778977, 32'sd0.10843703727635964, 32'sd-0.0020853983432791673, 32'sd-0.025048743260247322, 32'sd0.007494636774925802, 32'sd0.03978470747494422, 32'sd-0.020271413736263837, 32'sd0.10405815185796789, 32'sd-0.018294378113175917, 32'sd0.016013096806692266, 32'sd-0.01863552299912548, 32'sd-0.05266510043290119, 32'sd-0.09059973932689515, 32'sd-0.0058118694731219365, 32'sd-0.07867043918785704, 32'sd-0.10239531394253142, 32'sd-0.03077289926195984, 32'sd0.027275579856563155, 32'sd0.04566073943475252, 32'sd-0.007174489924456035, 32'sd1.0118604364054224e-118, 32'sd0.08136443612754916, 32'sd0.038083847159673646, 32'sd0.03238793198341037, 32'sd0.0175106744275287, 32'sd-0.014280858303284776, 32'sd-0.11974613555947969, 32'sd-0.04737896857374242, 32'sd-0.09971765137138307, 32'sd0.04901699237102904, 32'sd-0.030483119151755878, 32'sd0.1577708204285994, 32'sd-0.037954330255571773, 32'sd0.020276026633201768, 32'sd0.18849414983110094, 32'sd0.0773805905832495, 32'sd0.004710484737474883, 32'sd0.013959707407657623, 32'sd-0.14385035927592926, 32'sd0.0008668179955710626, 32'sd0.011328917130332133, 32'sd-0.1464119153961642, 32'sd-0.0862079032977408, 32'sd-0.09356429445984293, 32'sd-0.06338377165421803, 32'sd-0.11864769296114647, 32'sd-0.05394256342359858, 32'sd0.08221092715909857, 32'sd-3.295094360960226e-121, 32'sd0.04036189483061159, 32'sd-0.021748062370810815, 32'sd0.024361401614096855, 32'sd0.06314381458769985, 32'sd0.07439041182249878, 32'sd0.015748296956375578, 32'sd0.004659827329881088, 32'sd0.029864855840440373, 32'sd-0.025942566172546807, 32'sd0.06100182125542892, 32'sd0.12178572552171262, 32'sd0.005625818063266604, 32'sd0.08090604489484264, 32'sd0.11194194966584503, 32'sd0.1883444845639539, 32'sd-0.017462942219109715, 32'sd-0.16744958989952857, 32'sd-0.07903290977678445, 32'sd-0.13458597452710883, 32'sd0.02612991538166231, 32'sd-0.08849567261808272, 32'sd-0.14375632813864148, 32'sd-0.1455533365499508, 32'sd-0.09480035389650913, 32'sd-0.11824672314677936, 32'sd0.10170481994613222, 32'sd0.052866716490417416, 32'sd0.022887315861631837, 32'sd0.014625897735775798, 32'sd-0.07231705902253995, 32'sd-0.06515993279038873, 32'sd0.010175417645170317, 32'sd0.04920160056246091, 32'sd0.08112935599263854, 32'sd-0.06615562907723978, 32'sd-0.04781161214917647, 32'sd-0.1236895703512699, 32'sd0.05021958583558361, 32'sd0.07818238819616263, 32'sd-0.024799899721319258, 32'sd0.12804185668497742, 32'sd0.12085048719502849, 32'sd0.03252578553806786, 32'sd-0.12231828578556139, 32'sd-0.20051432228851335, 32'sd-0.08667353733092636, 32'sd-0.1359578663454177, 32'sd0.007310211609445984, 32'sd-0.07702583287390612, 32'sd0.01206821676460619, 32'sd-0.12105490263112578, 32'sd-0.10746289490437663, 32'sd-0.12567896110070442, 32'sd0.01865675370799366, 32'sd-0.01891425776820706, 32'sd0.025496728812543064, 32'sd0.02510346798134415, 32'sd0.08592807586085521, 32'sd0.059110773845305435, 32'sd0.025396283829006897, 32'sd-0.06295716181727652, 32'sd-0.06652549727934423, 32'sd-0.09557320026792851, 32'sd-0.14369647342617747, 32'sd-0.12163378287392951, 32'sd-0.02162246764599574, 32'sd0.09876301922407492, 32'sd0.1148273738818079, 32'sd0.08135129240856177, 32'sd0.013380869160268052, 32'sd-0.1895986307846814, 32'sd-0.043234380245606316, 32'sd-0.09070551461737851, 32'sd-0.11507047506532614, 32'sd0.027763050232976982, 32'sd-0.06934447017598674, 32'sd-0.0450507009588506, 32'sd-0.06553686223194825, 32'sd-0.1647213766243602, 32'sd0.00740916252939017, 32'sd-0.00042196904880030333, 32'sd0.09579585321545381, 32'sd0.05716084003017655, 32'sd0.09391373882454962, 32'sd0.048965771132733094, 32'sd0.06011396731599131, 32'sd0.039654068693914975, 32'sd-0.09305371248823965, 32'sd0.0018641754003374282, 32'sd0.0236325473720848, 32'sd-0.08343343112604085, 32'sd-0.053093715937337305, 32'sd0.10832198339281046, 32'sd-0.010887886326467911, 32'sd0.120803337934789, 32'sd0.0924766560658427, 32'sd0.07918699091156249, 32'sd-0.05010883728667946, 32'sd-0.2267670636609748, 32'sd-0.07944357900295851, 32'sd0.015412554856742396, 32'sd-0.014232667537230464, 32'sd-0.07515859035339949, 32'sd0.042369494586025305, 32'sd0.069238331903504, 32'sd-0.006697011937990356, 32'sd-0.15963243266901156, 32'sd-0.12533211372144373, 32'sd0.0279232747782384, 32'sd0.018476856185594064, 32'sd0.009476559814882735, 32'sd-0.031525567199521896, 32'sd0.006442021451821601, 32'sd-0.023120608313817362, 32'sd0.042570234289779046, 32'sd-0.011095677212147756, 32'sd-0.09716675939071401, 32'sd-0.0734306394086836, 32'sd0.017961285781078886, 32'sd0.11732541311138246, 32'sd0.051486597117203575, 32'sd0.012835462805559457, 32'sd-0.013989100438987195, 32'sd0.013140570828631877, 32'sd-0.14797709829046152, 32'sd-0.2844134548641679, 32'sd-0.17222552954703224, 32'sd-0.01361146540265829, 32'sd0.019259889773313353, 32'sd0.04574433470483276, 32'sd0.042763037954341415, 32'sd-0.0225700272169643, 32'sd0.07758110854072163, 32'sd0.008439338178571636, 32'sd0.015063379207339432, 32'sd-0.16803097948976048, 32'sd-0.10075417982819568, 32'sd-0.00971570769240579, 32'sd0.03999742908682229, 32'sd-0.015051079895799924, 32'sd0.10644652778243467, 32'sd-0.05374288233972094, 32'sd-0.049617427245277596, 32'sd-0.06795408555934872, 32'sd-0.0717093588649806, 32'sd-0.03810916036725332, 32'sd-0.07533517716439714, 32'sd0.053072459563041234, 32'sd0.035440313268250215, 32'sd0.06909044815332752, 32'sd0.00222457365486224, 32'sd0.01923080180182656, 32'sd-0.17445664685337736, 32'sd-0.30901116377480053, 32'sd-0.07006249137387632, 32'sd0.03996893637766225, 32'sd0.017923953758671275, 32'sd-0.0023870386797729304, 32'sd-0.027883331341513974, 32'sd0.011899098470319485, 32'sd0.11896042184009471, 32'sd-0.06880027364379916, 32'sd-0.02057468054612277, 32'sd-0.05867049554946437, 32'sd-0.016732274180179738, 32'sd0.0245649979157688, 32'sd-0.03341444455662523, 32'sd0.015290161445047941, 32'sd0.013538347547436639, 32'sd-0.023793902110388853, 32'sd0.027766668742011464, 32'sd-0.023186074514949223, 32'sd0.09154346534393328, 32'sd0.02091973741528291, 32'sd0.0983679919752758, 32'sd-0.00843797612330587, 32'sd0.03215578153937482, 32'sd0.03837788825963169, 32'sd-0.039122797933991246, 32'sd-0.10858670488443548, 32'sd-0.15001455645990402, 32'sd-0.10129377301152691, 32'sd0.13719195078655747, 32'sd0.07917591784807639, 32'sd0.13166986959890914, 32'sd0.07597204712898702, 32'sd0.06214026460283938, 32'sd0.1031992018811406, 32'sd0.1702631589286794, 32'sd0.012091437572119848, 32'sd0.10243874497987686, 32'sd0.038994391036245704, 32'sd-0.07067410142805979, 32'sd0.06487769211827119, 32'sd-0.01981530403850393, 32'sd0.02193779796144953, 32'sd-0.031167485299309086, 32'sd-0.06784618053291219, 32'sd-0.03413341942576511, 32'sd-0.027284775389025403, 32'sd-0.02629398333283874, 32'sd0.09816867493661938, 32'sd0.19817056291428878, 32'sd0.11161349197780966, 32'sd-0.04823356997538035, 32'sd0.09525378216675622, 32'sd-0.08721137976260945, 32'sd-0.043038058836540674, 32'sd-0.08595346640521725, 32'sd0.030091424442024797, 32'sd0.02865358726784749, 32'sd0.07070708072265766, 32'sd0.018511917592307272, 32'sd-0.004402530311761354, 32'sd0.09367701529290809, 32'sd-0.007417466018855678, 32'sd0.08227791382105841, 32'sd0.10565026868653797, 32'sd0.08211822553652187, 32'sd0.03355077519985174, 32'sd-0.039252700628296965, 32'sd-0.027104885507373312, 32'sd0.0029757920441561966, 32'sd-0.062169315553933846, 32'sd-0.014343939683934333, 32'sd-0.0023827368742991655, 32'sd-0.01371358213270427, 32'sd0.003723879668594413, 32'sd0.12812414922522816, 32'sd-0.0033354842576899094, 32'sd0.06698171952696134, 32'sd0.0835289262940252, 32'sd0.11261227879316202, 32'sd-0.012601982902031577, 32'sd-0.013370650932793231, 32'sd-0.06899279581665374, 32'sd-0.07664839489875976, 32'sd-0.08420153486727358, 32'sd0.17344805915506875, 32'sd0.13971503884621153, 32'sd-0.06348531766404646, 32'sd0.09327217588704893, 32'sd0.019137782760893184, 32'sd-0.003346817144474101, 32'sd-0.009674859998066714, 32'sd0.050248423895717834, 32'sd0.0685630019558951, 32'sd0.0708851021132107, 32'sd-0.09783302744683854, 32'sd-0.02009374821604939, 32'sd-0.03138321840045629, 32'sd0.011603749949194829, 32'sd0.06205284863346572, 32'sd0.021946143993739415, 32'sd-0.036445728551901306, 32'sd-0.12508043843900293, 32'sd0.06607706186526051, 32'sd0.06752123541719508, 32'sd0.17865641084808728, 32'sd0.05861008422298772, 32'sd-0.0046899536907626625, 32'sd0.12036822888064098, 32'sd0.11360147083808485, 32'sd-0.03181642207980896, 32'sd-0.10779867770294986, 32'sd-0.09143263081440706, 32'sd-0.021267431366438362, 32'sd0.04867405947716003, 32'sd-0.02008667446727286, 32'sd0.04498649012014812, 32'sd-0.008732179494460233, 32'sd-0.00553454429972061, 32'sd-0.007883691032979165, 32'sd0.10366401795442262, 32'sd0.10341608942945972, 32'sd0.07888201952230464, 32'sd0.021225086451932013, 32'sd-0.13683476301437775, 32'sd0.03145571198975522, 32'sd0.03915737757555669, 32'sd-0.08005948021219364, 32'sd-0.03602316222053462, 32'sd-0.03265092461219678, 32'sd-0.07427467347952643, 32'sd-0.048239505115936866, 32'sd0.008646862385878043, 32'sd0.09951680475116041, 32'sd0.09845676037190938, 32'sd0.08642103558275874, 32'sd0.09809806435283323, 32'sd0.10190104370308074, 32'sd0.08164242041233966, 32'sd0.013365968783034757, 32'sd-0.026451261357138565, 32'sd-0.013470323193324219, 32'sd-0.23088376971962665, 32'sd-0.1287196231067613, 32'sd-0.04160073817165885, 32'sd-0.008908887664022534, 32'sd0.0111103038775924, 32'sd-0.07760152319610239, 32'sd-0.009947207620618645, 32'sd0.028101663126022646, 32'sd0.12259171917966968, 32'sd-0.03210782101070117, 32'sd-0.024165475286866103, 32'sd0.033055303868958275, 32'sd-5.257872186779376e-124, 32'sd0.07453394880656773, 32'sd0.002529249495207726, 32'sd-0.05559580557538544, 32'sd0.03074199198395309, 32'sd-0.005831944650261652, 32'sd-0.01448914138860232, 32'sd0.06934389202935816, 32'sd0.09456594860019318, 32'sd0.0876468831658941, 32'sd0.08875510094688957, 32'sd0.11786683371464825, 32'sd0.06451347386925738, 32'sd0.08731250225139632, 32'sd0.09012296151572756, 32'sd-0.1365952930806067, 32'sd-0.168704647481924, 32'sd-0.1460503592544092, 32'sd-0.12823243958252498, 32'sd0.05375838988110613, 32'sd0.09349879173187599, 32'sd-0.01498603919585384, 32'sd0.10268888648543162, 32'sd0.12437085677423625, 32'sd0.08673008733688482, 32'sd-0.053853695095160255, 32'sd-0.10604424235076484, 32'sd-0.05359213442742904, 32'sd0.023324522456262327, 32'sd-0.03584693652077839, 32'sd0.0222582243314535, 32'sd-0.03372711130822393, 32'sd-0.043367664991592954, 32'sd0.06731903136227942, 32'sd-0.0756636122707801, 32'sd-0.08654952607731616, 32'sd0.05609411835868111, 32'sd0.08967527749069068, 32'sd0.11074466099124951, 32'sd0.29755868021788257, 32'sd0.24435064634800546, 32'sd0.05614044340712805, 32'sd-0.08929048668909075, 32'sd0.012804356299734764, 32'sd-0.06836102434047961, 32'sd-0.15771888743168033, 32'sd-0.0009625162893430593, 32'sd0.08688521585504505, 32'sd0.03735555077317724, 32'sd-0.038212448005644835, 32'sd0.11145647622625673, 32'sd0.03904691698137721, 32'sd0.026297811994543323, 32'sd-0.0821525009828255, 32'sd0.011763978466483032, 32'sd0.036490744757606934, 32'sd0.03685787449679181, 32'sd-0.004725638920290662, 32'sd0.006466303673955281, 32'sd0.016901714452846016, 32'sd-0.053085831145155624, 32'sd-0.059475958840455354, 32'sd-0.10122912271559704, 32'sd-0.08375383649147806, 32'sd-0.15339956737055999, 32'sd-0.03943030864503976, 32'sd0.050572279062033335, 32'sd0.14759850469629865, 32'sd0.22232918284448677, 32'sd0.06589917629130028, 32'sd-0.05565421712484616, 32'sd0.02413161931134767, 32'sd-0.03295721576579448, 32'sd0.033798034598759324, 32'sd0.07714760476467983, 32'sd0.06163893815035955, 32'sd0.041945855761520795, 32'sd0.07691659614518928, 32'sd0.02648416065716021, 32'sd-0.05877819635829285, 32'sd0.015287250949918573, 32'sd-0.1139842090757904, 32'sd0.0419219788422801, 32'sd-0.08612233464449491, 32'sd-1.8037204561567666e-121, 32'sd0.00639229925758056, 32'sd0.035629094676023584, 32'sd0.04278584089380053, 32'sd-0.0012976154749661083, 32'sd0.00035840337407264686, 32'sd-0.09483604736027394, 32'sd-0.03255866040005949, 32'sd-0.0978372154690242, 32'sd-0.10145313172983221, 32'sd-0.057474973425416645, 32'sd0.006420378407516631, 32'sd7.266827121799206e-05, 32'sd0.08296306819910428, 32'sd0.06135491105684515, 32'sd0.10879000965554818, 32'sd0.03581583111760946, 32'sd0.04692168458092105, 32'sd0.011077191032653222, 32'sd0.06306651867295734, 32'sd-0.001753793824699187, 32'sd0.10193096244337346, 32'sd0.06642281330028836, 32'sd-0.025163124640063806, 32'sd0.0038340102055972876, 32'sd-0.007342223850372849, 32'sd0.060118979936979754, 32'sd0.03746225937116707, 32'sd0.014414695459062127, 32'sd-0.010022858637908905, 32'sd-0.0761618292224182, 32'sd0.05306628356417089, 32'sd0.014552501561846929, 32'sd-0.022454784284796584, 32'sd0.06536961943343306, 32'sd-0.041077775047562985, 32'sd-0.06736234120208003, 32'sd-0.11629719775108589, 32'sd-0.11529761325143476, 32'sd-0.09404046941264138, 32'sd-0.04469952612681617, 32'sd-0.07119386282406416, 32'sd0.18720200369774792, 32'sd0.2056177228579451, 32'sd0.060136291910632744, 32'sd0.06758426271246659, 32'sd0.05963795155131225, 32'sd-0.06666297246230383, 32'sd0.043921072865142026, 32'sd0.02095738987957862, 32'sd0.028058160485974586, 32'sd-0.052914276968664874, 32'sd-0.10859627781049405, 32'sd-0.05618966858693628, 32'sd0.020679265664372407, 32'sd0.021810837150380947, 32'sd0.020192621318781336, 32'sd-0.04756898157139078, 32'sd-0.05962333598242167, 32'sd-0.04963779196166572, 32'sd-0.037381124043216224, 32'sd0.041280734357645156, 32'sd0.02930306750050293, 32'sd-0.002207682908447961, 32'sd-0.03552892010520537, 32'sd0.0015481252482007594, 32'sd-0.18008548966777788, 32'sd-0.13153621062512544, 32'sd-0.048207381714986446, 32'sd0.04680382139288572, 32'sd0.09209022547170233, 32'sd0.06571993703018264, 32'sd0.13823452674725858, 32'sd0.0741257408453379, 32'sd-0.018831187774450895, 32'sd-0.01100777500219014, 32'sd-0.003071155329437953, 32'sd0.08138241368186035, 32'sd-0.03952377658583016, 32'sd-0.14295965940895797, 32'sd-0.09865703380180812, 32'sd-0.09502603827970295, 32'sd0.0872870817492546, 32'sd0.01990542652873807, 32'sd-6.014482715899934e-121, 32'sd-0.034079174868575965, 32'sd0.03432695367634356, 32'sd0.01402552467623462, 32'sd-0.0010656276086485046, 32'sd0.010287070477438797, 32'sd-0.011802846950883553, 32'sd0.03980046027128196, 32'sd-0.054905120983564565, 32'sd-0.01398550385746066, 32'sd0.03280198493600675, 32'sd-0.038970906352505254, 32'sd-0.08617704141657216, 32'sd-0.004980604379663255, 32'sd0.1540778229295219, 32'sd-0.053422225222148914, 32'sd-0.07825824421233256, 32'sd0.01582473737514108, 32'sd-0.006330540491616735, 32'sd0.029999179428027774, 32'sd0.08290477707967944, 32'sd0.00566755494841643, 32'sd-0.023136502489599368, 32'sd-0.07246202131968767, 32'sd-0.10601067900091475, 32'sd-0.03235213699011135, 32'sd0.04265865472417952, 32'sd-1.537946017171973e-115, 32'sd-4.142401327625928e-125, 32'sd-1.1338649028604982e-122, 32'sd-0.005108050727553186, 32'sd0.0362094886302314, 32'sd-0.02484320139269317, 32'sd-0.024239485245310628, 32'sd0.0856418150527059, 32'sd0.06305278102921054, 32'sd0.022749094787188364, 32'sd0.016837988670896257, 32'sd-0.016347113934819683, 32'sd-0.014397410560173978, 32'sd-0.025562248139926417, 32'sd0.19867320312857184, 32'sd0.035101659484783394, 32'sd0.037461032125967665, 32'sd0.17433850136169898, 32'sd0.0005146911052772428, 32'sd0.03731624755827692, 32'sd-0.052875808114446296, 32'sd-0.09579957638450358, 32'sd0.025834225390374152, 32'sd-0.05283175250277638, 32'sd0.09495396405957594, 32'sd-0.01990868640633883, 32'sd0.0326526397004792, 32'sd0.01091976796700003, 32'sd-1.5698872563278472e-124, 32'sd4.116824553001184e-118, 32'sd-4.783753528467836e-117, 32'sd-0.05384826156055707, 32'sd-0.05471882891264965, 32'sd0.004125872863714595, 32'sd0.026166989100454067, 32'sd-0.06437645869487363, 32'sd0.014154226187188632, 32'sd0.12395602286663195, 32'sd0.04315171752654044, 32'sd-0.017364277880882812, 32'sd0.005205018129818348, 32'sd0.015685910533258737, 32'sd0.10874106096554349, 32'sd0.032085258102253524, 32'sd-0.01118320957382866, 32'sd-0.014670820565293431, 32'sd-0.01714189171611187, 32'sd-0.0029946635473544585, 32'sd0.0844192985009877, 32'sd-0.026433282781167414, 32'sd-0.008315538552441921, 32'sd-0.019105798979841, 32'sd0.12627116350142853, 32'sd-0.004530510250088315, 32'sd0.036101714663591675, 32'sd0.05316962228170098, 32'sd3.2252225438016447e-122, 32'sd2.233529721062806e-126, 32'sd-8.058890108311604e-116, 32'sd3.1773633187271954e-120, 32'sd0.03841168478547495, 32'sd0.015531264537351302, 32'sd-0.00869408692792084, 32'sd-0.07929022938574547, 32'sd0.011284225140770387, 32'sd0.04486745971153979, 32'sd-0.09258804038831381, 32'sd-0.1578034885386953, 32'sd-0.06629502179840073, 32'sd-0.04453522340864958, 32'sd-0.11758724844469744, 32'sd0.010840878601423548, 32'sd-0.06432450958646707, 32'sd0.054007965604630705, 32'sd-0.0854813062745853, 32'sd-0.080937747356467, 32'sd0.062007951383060644, 32'sd0.0916783224772492, 32'sd-0.018387718056850886, 32'sd-0.12636791596208125, 32'sd-0.09503085759499534, 32'sd-0.010761219278100911, 32'sd0.07659511843146949, 32'sd-1.190211439399758e-121, 32'sd-7.0557425860354425e-115, 32'sd-1.5146154631650418e-116, 32'sd4.221272818266704e-117, 32'sd-3.1140568138544265e-125, 32'sd-1.1804709464296743e-125, 32'sd0.10287301262402475, 32'sd0.003528515617291592, 32'sd0.05896875334524129, 32'sd0.08640451067656736, 32'sd0.09101540172389046, 32'sd-0.006225913750501907, 32'sd0.06533226282025684, 32'sd0.016586214172633385, 32'sd0.08434497137341844, 32'sd-0.028254479794523196, 32'sd-0.04222279291012858, 32'sd-0.046744110010517495, 32'sd0.008128016612135143, 32'sd0.01849723682866588, 32'sd0.007311113903884326, 32'sd-0.010006080917242479, 32'sd0.013472252507345583, 32'sd-0.04074397791784064, 32'sd0.010927379914938792, 32'sd0.06971996436716701, 32'sd8.867105741297906e-127, 32'sd-7.911455977888364e-117, 32'sd-2.631195153861816e-118, 32'sd5.854711111876575e-117},
        '{32'sd3.318254968438445e-118, 32'sd8.82717520939195e-127, 32'sd9.322886404675698e-121, 32'sd-1.0401163588290068e-122, 32'sd4.83365538328934e-118, 32'sd1.416088692339165e-124, 32'sd2.609591385326196e-116, 32'sd-1.3605143192866176e-123, 32'sd-7.046942549476053e-128, 32'sd-9.82351708063763e-122, 32'sd-9.116057367956231e-122, 32'sd3.214332607198129e-121, 32'sd0.007883776760953755, 32'sd-0.005397131982459687, 32'sd-0.00944152657733016, 32'sd0.06819528072541811, 32'sd4.265090497004275e-125, 32'sd1.3706989630934626e-118, 32'sd-9.951593461452645e-116, 32'sd2.9996377569407413e-115, 32'sd-2.2845545778058217e-125, 32'sd3.3374146103560374e-121, 32'sd-2.6564808885259792e-120, 32'sd2.5342849475275592e-114, 32'sd-1.49041499817361e-119, 32'sd-2.294896041693073e-121, 32'sd1.3796358681330966e-122, 32'sd-9.075580594236585e-128, 32'sd-1.4290497207428855e-118, 32'sd-9.895559494668018e-116, 32'sd-1.0561303745350228e-119, 32'sd3.447440815447975e-125, 32'sd0.07231235218706278, 32'sd0.028886347187084625, 32'sd0.04130685879304055, 32'sd0.09708853683902255, 32'sd-0.020892662566583987, 32'sd-0.06599472797092171, 32'sd-0.03577259457243071, 32'sd-0.008732122238800329, 32'sd0.03678182272426225, 32'sd-0.0377372206382568, 32'sd-0.020743796427712582, 32'sd0.010757796187145273, 32'sd-0.023680419379104707, 32'sd0.07038774633908017, 32'sd0.020350414567751902, 32'sd0.044785632223949226, 32'sd-0.030679872849434776, 32'sd0.10850890781401615, 32'sd0.04825282908793742, 32'sd0.03859024150862815, 32'sd2.141612980808202e-124, 32'sd-5.0696028999111575e-121, 32'sd1.2032428240903524e-122, 32'sd1.42029633196625e-120, 32'sd-1.4480909240532225e-125, 32'sd-4.752888078319529e-127, 32'sd0.11224894271917998, 32'sd0.05927650982843544, 32'sd0.0937910264126159, 32'sd-0.015749151793198666, 32'sd-0.012444200990172512, 32'sd0.036201259852374906, 32'sd0.10076191686907521, 32'sd0.06543843479695478, 32'sd-0.007972613423139376, 32'sd-0.03380344907340846, 32'sd-0.12039526600919594, 32'sd-0.009228755361885171, 32'sd-0.13561783557322882, 32'sd-0.03654543746133284, 32'sd0.031994678923455346, 32'sd0.1857661285407106, 32'sd0.18490450602141706, 32'sd0.018153314444983516, 32'sd0.06942420263133395, 32'sd-0.07664293918890402, 32'sd0.06439863606351102, 32'sd0.05996788358705808, 32'sd0.0825580738268462, 32'sd0.07072436469259871, 32'sd2.3688937120736556e-120, 32'sd9.499175829912662e-120, 32'sd-3.774105980633912e-124, 32'sd-1.3089120048523728e-118, 32'sd0.07815587438694435, 32'sd0.025141458662345132, 32'sd-0.016236481973728324, 32'sd0.04399593493549939, 32'sd0.13884171977302223, 32'sd-0.012265346936623223, 32'sd0.060724871607111, 32'sd0.018442893385887598, 32'sd-0.05493988355584408, 32'sd-0.03685142037551101, 32'sd-0.07778030888573911, 32'sd0.08844172581752699, 32'sd0.0242117495168132, 32'sd0.0024440401355836903, 32'sd0.08502779936540825, 32'sd-0.055500452898134926, 32'sd0.07830136665369858, 32'sd0.036047124256954347, 32'sd-0.04693870509728253, 32'sd0.07019917064622846, 32'sd-0.010045681586643651, 32'sd0.025525869544157812, 32'sd-0.07656203398028345, 32'sd0.09265454757651462, 32'sd-0.032824144881180135, 32'sd-6.376507021356064e-121, 32'sd3.5973844258744e-119, 32'sd0.07312508815824471, 32'sd0.02119012868678711, 32'sd0.02902796531029685, 32'sd0.06508471859306453, 32'sd0.03975383365620463, 32'sd0.07241049092397979, 32'sd0.04837810610171184, 32'sd-0.019500815769650324, 32'sd-0.08055130137309385, 32'sd0.0034323612999749924, 32'sd0.004728773565305636, 32'sd0.006368943588802684, 32'sd-0.10758873429765047, 32'sd0.08243372170844158, 32'sd0.05754895777092246, 32'sd0.007077350489092819, 32'sd0.06132018157541565, 32'sd0.08870018986773633, 32'sd0.06498456080627067, 32'sd0.09356461430557533, 32'sd0.06111357569741023, 32'sd-0.11149958553350069, 32'sd0.0730603928028324, 32'sd0.10902092187361871, 32'sd-0.03261730949010012, 32'sd0.024664849640416278, 32'sd0.0006283922094260481, 32'sd-6.930769224030133e-120, 32'sd0.0353615786750488, 32'sd0.02599636703954424, 32'sd-0.13240059911585586, 32'sd-0.005052848858583998, 32'sd-0.026229842064064562, 32'sd0.012775257939138798, 32'sd-0.09701903398212205, 32'sd0.011965776738672766, 32'sd-0.0716590434757067, 32'sd0.09102212587055332, 32'sd0.08225232996235085, 32'sd0.1476017416057771, 32'sd0.05438747636593275, 32'sd0.06929801502816782, 32'sd0.1436229379782572, 32'sd0.20284103471927464, 32'sd0.1447462239738422, 32'sd0.19640583177556326, 32'sd0.07840271397854752, 32'sd0.09602373399588589, 32'sd0.18471511594631493, 32'sd0.09415669798359898, 32'sd0.1253575999861179, 32'sd0.1692231594721626, 32'sd-0.05508042264661108, 32'sd-0.04378094968543149, 32'sd0.059789290778152086, 32'sd-5.101402926999426e-121, 32'sd0.01898644183752582, 32'sd-0.026459149426475405, 32'sd-0.0711671080038853, 32'sd0.019434406915604652, 32'sd-0.06527315235451736, 32'sd-0.036750423024368505, 32'sd0.09416956955172857, 32'sd0.09959087051502771, 32'sd-0.02869101264181357, 32'sd0.057566972469960294, 32'sd0.21546413776126028, 32'sd0.07523051682707776, 32'sd0.05432240464465816, 32'sd0.058049731035051746, 32'sd0.21764747748925178, 32'sd0.18140440930814342, 32'sd0.14558286085691705, 32'sd0.14439578641641448, 32'sd0.1590732211054468, 32'sd0.04362723919847855, 32'sd0.0032342292767117043, 32'sd0.0020492017210154982, 32'sd0.0013025634225897465, 32'sd0.14653106968427707, 32'sd-0.017392474030654272, 32'sd-0.040084332271598584, 32'sd0.013113408895352337, 32'sd0.027146571829866982, 32'sd0.11899810114395162, 32'sd-0.05301918080578163, 32'sd-0.06700326585840978, 32'sd-0.02631949955908836, 32'sd0.06866965319650213, 32'sd0.06209033562733275, 32'sd-0.028674501444212918, 32'sd0.04398932100817255, 32'sd0.024644866373284325, 32'sd0.031361327034844386, 32'sd0.07956305915636504, 32'sd0.07181272611414112, 32'sd0.014812391145437826, 32'sd0.13263905158135986, 32'sd0.016867828479977573, 32'sd0.09829070328724684, 32'sd-0.02309782980423958, 32'sd-0.019368515232225308, 32'sd-0.041924495846215416, 32'sd-0.13347706414462826, 32'sd-0.08092887901484411, 32'sd-0.016758425286004387, 32'sd-0.2000606536187101, 32'sd-0.1122447572742875, 32'sd0.03976540627895329, 32'sd0.019429111061320038, 32'sd0.05955583492360307, 32'sd0.07733261715086637, 32'sd0.03080931434814151, 32'sd-0.0010060108524427502, 32'sd-0.02435064564296902, 32'sd-0.021192135795843874, 32'sd-0.0548522071722747, 32'sd0.017817603452017394, 32'sd-0.022916386252774545, 32'sd0.026007289774629138, 32'sd0.002814580767115171, 32'sd0.04395262473187804, 32'sd0.08473842789770031, 32'sd0.0719689423837751, 32'sd-0.023052202727471945, 32'sd0.05718954038879842, 32'sd-0.16220982164322184, 32'sd-0.204295288110136, 32'sd-0.1378427977401692, 32'sd-0.03921050280700169, 32'sd-0.13103320149600467, 32'sd-0.21490382460773502, 32'sd-0.10724261623832756, 32'sd-0.021647903619315765, 32'sd-0.20060228464758056, 32'sd-0.18116646129330904, 32'sd-0.07926398114009382, 32'sd0.020092419272228604, 32'sd-0.01269028069308507, 32'sd0.025761279559176526, 32'sd-0.029716141403275522, 32'sd-0.007398569132532904, 32'sd-0.005231250106528008, 32'sd-0.019243700293403262, 32'sd-0.0272509072035026, 32'sd0.11495811219276357, 32'sd-0.0044186849807603705, 32'sd0.027405649091436043, 32'sd-0.01578886234500683, 32'sd0.08791205846363333, 32'sd-0.05424397669016307, 32'sd-0.05928008457853182, 32'sd-0.009008113701142939, 32'sd-0.07512955970419782, 32'sd-0.21263844918519528, 32'sd-0.2508275781101314, 32'sd-0.07615981020659073, 32'sd-0.08791198009103326, 32'sd-0.22797949789675823, 32'sd-0.17723274783430745, 32'sd-0.08560196546759397, 32'sd-0.11386256690944375, 32'sd-0.2975760894883103, 32'sd-0.059301791348481805, 32'sd-0.06467141091916973, 32'sd-0.03148714120219117, 32'sd0.034661763819943264, 32'sd0.014550759533838015, 32'sd-0.10209707022435223, 32'sd-0.055391171194523504, 32'sd-0.08190394651960914, 32'sd-0.036617722863743235, 32'sd0.07333316567086288, 32'sd0.13628153141062607, 32'sd-0.00046236250431205275, 32'sd0.010068851947312895, 32'sd0.0001079833066181419, 32'sd-0.07478562008972282, 32'sd-0.11637700270852702, 32'sd-0.13322972288493895, 32'sd-0.14690956855615905, 32'sd-0.2597034151389877, 32'sd-0.2128525734225143, 32'sd-0.2339950882260673, 32'sd-0.2654124161776506, 32'sd-0.15089765301570238, 32'sd-0.17103637078379832, 32'sd-0.11805041616594916, 32'sd-0.12809939046979074, 32'sd-0.2162770593221895, 32'sd-0.046888084745046264, 32'sd-0.1422664155210873, 32'sd-0.06839596382802297, 32'sd-0.060086443278693, 32'sd-0.002303321768785482, 32'sd0.01656784746993354, 32'sd-0.017118149227209063, 32'sd0.034684296713215275, 32'sd-0.005951508731929205, 32'sd0.0915235674794158, 32'sd0.017103563258792587, 32'sd0.06330619357645256, 32'sd-0.058310743931021064, 32'sd-0.06389501646860125, 32'sd-0.12732816007666756, 32'sd-0.018970404399342746, 32'sd-0.1750161850248888, 32'sd-0.009603837008405858, 32'sd-0.16006968825444567, 32'sd-0.09828624926715127, 32'sd0.03378654247563993, 32'sd-0.10950826935043086, 32'sd-0.037655506913851305, 32'sd-0.02652605488488272, 32'sd-0.16670767051204866, 32'sd-0.16164360015637236, 32'sd0.0027830316974592055, 32'sd0.00850611030548071, 32'sd-0.05005817553812979, 32'sd0.0435646993813749, 32'sd-0.04250601679333253, 32'sd-0.029630212640012518, 32'sd-0.016802135670963662, 32'sd0.02537166362052236, 32'sd0.04526625966042789, 32'sd-0.05855761566716622, 32'sd0.13218823523882503, 32'sd-0.012435674564941372, 32'sd0.006071823086798162, 32'sd-0.044980767567516095, 32'sd-0.1128975371648463, 32'sd-0.05818143187249011, 32'sd-0.06807189869391614, 32'sd-0.0570818811910493, 32'sd-0.09031843801704433, 32'sd-0.08000903995701529, 32'sd-0.18659896892935707, 32'sd-0.020915678405426817, 32'sd0.09698225487215466, 32'sd0.044246048752529625, 32'sd0.07366801862652152, 32'sd-0.04107725163895117, 32'sd0.051715016141607194, 32'sd0.04239579384485486, 32'sd-0.04703218362405428, 32'sd-0.03379799126072329, 32'sd0.06862607090078847, 32'sd0.10938684301721958, 32'sd-0.06423803495756296, 32'sd-0.11275607635488853, 32'sd-0.021544613164743473, 32'sd0.01988551211470991, 32'sd-0.09966174540707992, 32'sd-0.005925052481943631, 32'sd0.01717974488326222, 32'sd-0.01725311636392113, 32'sd-0.09708037096555445, 32'sd-0.002524877212122861, 32'sd0.07564876736525586, 32'sd0.03062644710298019, 32'sd-0.056684232816394016, 32'sd0.019872895659054063, 32'sd0.02502866917708056, 32'sd-0.07795878928506203, 32'sd-0.06484228311934588, 32'sd0.05790425005980355, 32'sd0.007440078903720486, 32'sd0.0729634762894112, 32'sd0.07104316030279705, 32'sd0.07366084188572299, 32'sd0.1919067895410462, 32'sd0.22245375859561994, 32'sd-0.08951010107764565, 32'sd-0.07448468369252584, 32'sd0.007452928090812094, 32'sd0.0643966721338577, 32'sd0.004501728679925525, 32'sd0.010319695868946021, 32'sd-0.009556967485488, 32'sd0.12698652544942202, 32'sd0.06428067064889506, 32'sd0.011666735057124787, 32'sd0.051471621478713925, 32'sd0.049227576184500035, 32'sd0.059568253576460235, 32'sd0.028255638125049262, 32'sd-0.024591648397362276, 32'sd-0.008937658530610763, 32'sd-0.0508073198699876, 32'sd0.0936646116268219, 32'sd0.07828525819772995, 32'sd-0.07668542527060868, 32'sd-0.0501001584821146, 32'sd0.0018426650555764612, 32'sd-0.06322352944345362, 32'sd0.02212811268025159, 32'sd0.011157287489499304, 32'sd0.07506905014280268, 32'sd0.12184187513066, 32'sd0.10426240118035261, 32'sd0.004379685211109688, 32'sd-0.08096575617822106, 32'sd-0.034971351071419784, 32'sd0.0416723698283069, 32'sd-0.048606199556373575, 32'sd-0.01574955126224755, 32'sd0.027505724559478827, 32'sd0.051403118509977454, 32'sd0.010793880332680418, 32'sd0.02295154272218216, 32'sd0.004587076180749024, 32'sd-0.0500627668513828, 32'sd-0.010785507295519803, 32'sd0.1351791761134358, 32'sd0.09097977962429445, 32'sd0.11553123802231176, 32'sd0.005035859559046844, 32'sd-0.1050101845995565, 32'sd-0.1319371466433339, 32'sd-0.093217904943236, 32'sd-0.03210940096032416, 32'sd-0.021322419543715197, 32'sd-0.10847316163208762, 32'sd0.01378637338486258, 32'sd0.055226534700293976, 32'sd0.030767035736290037, 32'sd0.08749231888165804, 32'sd0.08369059217281052, 32'sd0.029295465135999777, 32'sd-0.1467807841604948, 32'sd0.05637838364527664, 32'sd0.014787447185241763, 32'sd0.08622272805483855, 32'sd0.03815057238238227, 32'sd-0.054373095570692066, 32'sd0.06909153292574993, 32'sd0.08065992891668047, 32'sd-0.039559306636967724, 32'sd0.07711016127499958, 32'sd0.08572601237003684, 32'sd-0.0066388103004411635, 32'sd-0.05529287323743527, 32'sd0.0019271189429589067, 32'sd-0.04337235017367565, 32'sd-0.046781104745404437, 32'sd-0.03145227164545906, 32'sd-0.06158439475343387, 32'sd0.026812115837065175, 32'sd0.06138319131982607, 32'sd-0.00660630793709235, 32'sd0.08281058363606912, 32'sd0.09227741309059471, 32'sd0.09630618580505412, 32'sd0.10644168830678721, 32'sd0.03449004370934259, 32'sd0.039791189650285434, 32'sd-0.020440442198548247, 32'sd-0.039170554538929474, 32'sd0.08947823361320033, 32'sd-0.0623197951847219, 32'sd0.03681531242855773, 32'sd-0.044312579986693766, 32'sd0.03490457548508543, 32'sd2.7510100178907068e-120, 32'sd-0.023114968011379636, 32'sd0.007959463358157321, 32'sd0.07616717778964478, 32'sd0.05994710677696692, 32'sd-0.027345286279016216, 32'sd-0.05282487525468393, 32'sd-0.15182308405113207, 32'sd-0.062150808117059926, 32'sd0.01640349365798565, 32'sd0.018298815055911216, 32'sd0.013197592155501117, 32'sd0.1412490029389167, 32'sd-0.013632494551036264, 32'sd-0.04735562704803375, 32'sd0.06769869846597032, 32'sd0.1193196138400467, 32'sd-0.02431520339104259, 32'sd-0.022603608962731125, 32'sd0.0025991061170114057, 32'sd0.009820408171801166, 32'sd0.04026531529349549, 32'sd0.050160080391984566, 32'sd-0.06725031622124678, 32'sd-0.07296392768521155, 32'sd0.014839153484922664, 32'sd-0.10100999721961086, 32'sd0.05896723648979244, 32'sd0.057796231176485635, 32'sd0.07838263372838979, 32'sd0.008281951683120934, 32'sd-0.0008572688483739049, 32'sd0.017692644092123313, 32'sd0.09449106882262666, 32'sd0.08415381072590525, 32'sd-0.15795777389035182, 32'sd-0.07260419466448231, 32'sd-0.10492259495388437, 32'sd0.12019857015341602, 32'sd0.15243255255939228, 32'sd0.0991244499545661, 32'sd0.020639169044533636, 32'sd0.03553600432264657, 32'sd0.08952753364388841, 32'sd0.04457669957209542, 32'sd-0.003001846893305199, 32'sd-0.00804505411578226, 32'sd0.018339451650522698, 32'sd-0.0371617875849866, 32'sd-0.053127944142158955, 32'sd0.06751040883648916, 32'sd0.005962759345469841, 32'sd-0.0026156475512254993, 32'sd0.048426596028807514, 32'sd-0.0183879625558356, 32'sd0.07031389243608342, 32'sd0.060166798537484606, 32'sd0.04532221948754231, 32'sd0.0017889216444574394, 32'sd-0.040921474729030814, 32'sd0.005621532229701049, 32'sd0.051458571800920706, 32'sd0.0022264028396631716, 32'sd-0.09861269441810398, 32'sd-0.03431584518868442, 32'sd-0.01625411311338227, 32'sd0.19841359758065408, 32'sd0.16423472417738816, 32'sd0.1377344647427901, 32'sd0.061692092907543614, 32'sd-0.02387205345037552, 32'sd-0.0446641052833443, 32'sd0.03625655095816575, 32'sd0.025601470757189545, 32'sd0.13486968549979633, 32'sd0.012284643963902246, 32'sd-0.060039201792652507, 32'sd-0.09576418380237113, 32'sd0.04932989334966943, 32'sd0.041960195536488165, 32'sd0.025065517474030397, 32'sd0.1276732091729353, 32'sd0.0979636670035236, 32'sd-0.052569200232064406, 32'sd-6.650135099525283e-124, 32'sd-0.07325873081894793, 32'sd0.06402417321732516, 32'sd-0.01475925311034813, 32'sd0.17498411838199757, 32'sd0.07255054563959891, 32'sd0.10051921262252839, 32'sd-0.018055872321799022, 32'sd-0.08463289453827763, 32'sd0.0948410703268516, 32'sd0.05692574163496438, 32'sd-0.0007720259126273324, 32'sd0.12430456722267394, 32'sd0.02262585316896823, 32'sd-0.013877673153514354, 32'sd-0.023042029566546038, 32'sd-0.04853533973926604, 32'sd0.03351262951609054, 32'sd0.06171878488767496, 32'sd-0.0134680716864991, 32'sd-0.035339559807519204, 32'sd0.02514622381371689, 32'sd0.058373989968433425, 32'sd0.09495121389281502, 32'sd0.053340234699644225, 32'sd0.0333511220077251, 32'sd-0.06893434142626925, 32'sd0.0358763193325012, 32'sd0.10324192774586781, 32'sd0.04740028731847988, 32'sd-0.06806896243756257, 32'sd0.06720351249007214, 32'sd0.10158191265331341, 32'sd0.04586459508717661, 32'sd0.13958602402013465, 32'sd-0.05325067543417965, 32'sd0.03520959969690638, 32'sd0.10067535261661024, 32'sd0.07330342660304616, 32'sd0.10283380149789555, 32'sd0.11437633022119349, 32'sd0.07437012144438121, 32'sd-0.0003894827036740074, 32'sd0.11619270427686242, 32'sd0.106740650244178, 32'sd0.013757702536635307, 32'sd0.06536670167212295, 32'sd0.02421862038482055, 32'sd-0.030628207898695352, 32'sd0.002099919055033602, 32'sd-0.010729142749987408, 32'sd0.07495446392995775, 32'sd0.07707605559170341, 32'sd-0.050915795649855475, 32'sd-0.04318852028635581, 32'sd0.07036070004639959, 32'sd-0.005063465514431026, 32'sd-0.0053608617786207475, 32'sd-0.04329583688420472, 32'sd0.046789051674316434, 32'sd0.06922478330764711, 32'sd0.07100912380539558, 32'sd-0.05388256497032793, 32'sd-0.010615000099866998, 32'sd0.02805707751611392, 32'sd0.08252451730267622, 32'sd-0.029339445959526672, 32'sd-0.02756732751831938, 32'sd0.08959240387276347, 32'sd-0.008806054425371091, 32'sd0.059695632187855154, 32'sd-0.02600090363035836, 32'sd-0.07232918280151658, 32'sd-0.11901827543205314, 32'sd0.024455639326918893, 32'sd-0.06744491915648253, 32'sd-0.03994406273958205, 32'sd0.02864158305353898, 32'sd0.08255682762600473, 32'sd0.09972881459809083, 32'sd0.011446345457289165, 32'sd0.04078437698370628, 32'sd-0.024273171014266483, 32'sd0.036657091344495775, 32'sd-1.0557659012912163e-116, 32'sd0.03695641459639222, 32'sd-0.08782927970160546, 32'sd-0.023162367588537496, 32'sd-0.01523798696080982, 32'sd0.08868678544334789, 32'sd-0.0941688972673811, 32'sd0.020410503525302742, 32'sd0.05257852165586959, 32'sd-0.07829367067654372, 32'sd-0.015486768171108152, 32'sd-0.1445184318807758, 32'sd0.0082062043558648, 32'sd-0.051572323891321686, 32'sd-0.03685325241052563, 32'sd-0.0011338291453371185, 32'sd-0.07166025125286035, 32'sd-0.08472715616724219, 32'sd-0.06426300999267388, 32'sd-0.016929789382021915, 32'sd0.0062830573713360816, 32'sd0.07890878376658789, 32'sd0.049617869514029835, 32'sd0.08263953653642782, 32'sd0.07443000992237297, 32'sd0.09083942257167088, 32'sd-0.02739403216979299, 32'sd-3.011450095890944e-116, 32'sd3.7944908767488107e-115, 32'sd3.7520086222511606e-122, 32'sd-0.02706801751522095, 32'sd-0.02341559710180081, 32'sd-0.02304712762110799, 32'sd0.025645960694679795, 32'sd-0.0974241248129616, 32'sd-0.032518102923988774, 32'sd-0.03696535350144351, 32'sd0.012636826702043195, 32'sd0.019356935778233882, 32'sd-0.060776039012240754, 32'sd-0.11422533846327218, 32'sd0.004572441387226568, 32'sd-0.011679076968684152, 32'sd-0.025746905638135267, 32'sd-0.03659755412006177, 32'sd0.01574116760195719, 32'sd0.101838865539631, 32'sd0.0350656819138132, 32'sd0.07562896753196449, 32'sd0.07159961634448296, 32'sd-0.014407760050015345, 32'sd-0.016749639471786173, 32'sd0.04137309469211985, 32'sd-0.027284735657483062, 32'sd0.026573753358963052, 32'sd-6.469165132070457e-119, 32'sd-8.454108030894457e-121, 32'sd3.0412102708943254e-120, 32'sd0.09259796716146847, 32'sd0.03765164581806103, 32'sd-0.0909093231548804, 32'sd0.02360438538512174, 32'sd-0.0835375529902364, 32'sd-0.033261732127790745, 32'sd-0.12486365034508387, 32'sd-0.13566206195656075, 32'sd-0.059295970137264294, 32'sd-0.012179108195913717, 32'sd0.05913133247987704, 32'sd-0.10555922413920882, 32'sd0.03295171031508097, 32'sd-0.0779844564440132, 32'sd0.046503940237528185, 32'sd0.010693484696676064, 32'sd0.044523782615247726, 32'sd0.05626510753368674, 32'sd0.04924170329412443, 32'sd-0.0035483853646373895, 32'sd0.03503156197436902, 32'sd0.10649250507269721, 32'sd0.08998247951954126, 32'sd0.049960832328277076, 32'sd0.025421452095928894, 32'sd2.883628535458931e-118, 32'sd7.909513154692478e-130, 32'sd-7.76499969475863e-123, 32'sd5.743456572293224e-123, 32'sd0.03708249657895279, 32'sd0.001500910367366074, 32'sd-0.013611523994148193, 32'sd-0.05125244617849805, 32'sd0.0425599116833369, 32'sd0.09504707390901333, 32'sd-0.014310570478986517, 32'sd0.06050876556451328, 32'sd0.008731526170396542, 32'sd0.001410721822202662, 32'sd-0.020983544699865787, 32'sd0.0034935146467250356, 32'sd-0.020092795059861873, 32'sd-0.07140484975728377, 32'sd-0.0049723341044674635, 32'sd0.04681725664849451, 32'sd0.08239436294021442, 32'sd0.1151442577799984, 32'sd0.011766514521962687, 32'sd0.024951681202535957, 32'sd0.030469637680321657, 32'sd0.1353208039273776, 32'sd0.05013237796264427, 32'sd-1.0578843013829188e-121, 32'sd1.6868721135877338e-116, 32'sd1.5863542627026295e-125, 32'sd9.325545965819841e-116, 32'sd-2.5715635970803902e-123, 32'sd-4.944533607586074e-122, 32'sd0.03190232885547138, 32'sd0.09511065841734993, 32'sd-0.0004109838626908269, 32'sd0.05413681366804121, 32'sd0.006006850099529618, 32'sd-0.006496375095504329, 32'sd0.06761335513678499, 32'sd0.06022857617512931, 32'sd0.005412588748508844, 32'sd0.036632122763774276, 32'sd0.11191818623201893, 32'sd0.060124015598232966, 32'sd0.03875893223333909, 32'sd-0.046831979293497576, 32'sd0.01603420007719653, 32'sd-0.001897893163659443, 32'sd0.0008057488919951624, 32'sd0.037055226762351096, 32'sd0.032098470187280834, 32'sd-0.018737016654286214, 32'sd3.4620838991994704e-116, 32'sd-6.866504966383186e-119, 32'sd-8.356416478540229e-117, 32'sd-1.3418908556955087e-118},
        '{32'sd5.627775897246409e-125, 32'sd-2.5473282392690375e-126, 32'sd-9.735162442326883e-115, 32'sd1.0303320551075065e-114, 32'sd6.636371334706435e-115, 32'sd-1.506187390084516e-116, 32'sd3.283461474829954e-120, 32'sd6.4285160112005975e-121, 32'sd2.3924268480622047e-126, 32'sd1.5485380773836298e-118, 32'sd-5.5818019813239425e-117, 32'sd-4.60851898211666e-123, 32'sd0.027223202401703273, 32'sd-0.08907684019115043, 32'sd-0.001556828298150854, 32'sd0.03304615299678536, 32'sd-6.264713169524408e-125, 32'sd-3.348161874100968e-116, 32'sd3.636760450832536e-116, 32'sd1.6814001894013494e-116, 32'sd9.087704725065917e-124, 32'sd-2.842460475808514e-121, 32'sd-3.991740724561488e-123, 32'sd-1.1819922430668995e-123, 32'sd5.496605348395271e-125, 32'sd7.528394156652281e-115, 32'sd4.963697874084345e-124, 32'sd-9.853178286837115e-123, 32'sd-6.450213625941719e-126, 32'sd-1.751834955539317e-123, 32'sd1.3608079911157299e-115, 32'sd-1.593479878013724e-123, 32'sd-0.005763749484374804, 32'sd-0.023634676400318366, 32'sd-0.012850577840207156, 32'sd0.002461471688946099, 32'sd-0.09013409730440897, 32'sd-0.021040736994160113, 32'sd0.02157251819565932, 32'sd-0.10780156068050668, 32'sd-0.07890984541979866, 32'sd-0.03194230915193508, 32'sd0.017783611355813078, 32'sd-0.12477302324654038, 32'sd0.08559998125226878, 32'sd0.023432243748224425, 32'sd0.0846698067611572, 32'sd0.10176037396853108, 32'sd-0.04363234705008163, 32'sd0.07671202064994595, 32'sd0.02348245553180037, 32'sd0.008213030928103035, 32'sd-7.465114250693467e-115, 32'sd-7.2261130842921095e-127, 32'sd-1.5464000976471743e-117, 32'sd1.077145908630869e-124, 32'sd3.6790186215727113e-119, 32'sd-1.4876424512121216e-115, 32'sd-0.028118541589025724, 32'sd-0.04583084419389728, 32'sd0.024460239489117356, 32'sd0.029734090429274513, 32'sd-0.039240629208783975, 32'sd0.016732149040519406, 32'sd-0.06389899361627213, 32'sd-0.03675879108647796, 32'sd-0.12576225813348368, 32'sd0.03572940746587167, 32'sd-0.150879714624035, 32'sd-0.0701943745774512, 32'sd0.02808844686475724, 32'sd0.06577048086949011, 32'sd-0.026791820558951462, 32'sd0.1769427386767912, 32'sd0.06237247759581416, 32'sd0.08977108388075411, 32'sd-0.010852859081130763, 32'sd0.09362031536168848, 32'sd0.11280867088502837, 32'sd-0.011499231486255328, 32'sd0.019289019286642006, 32'sd-0.04404085014981252, 32'sd3.0856664755330056e-121, 32'sd6.927698225579465e-123, 32'sd-1.5744797868348947e-123, 32'sd-7.69057284688103e-127, 32'sd-0.020783154669638343, 32'sd-0.018490547135721215, 32'sd0.0828554230307076, 32'sd-0.09239059883614582, 32'sd-0.05175328822063446, 32'sd0.003877614128639723, 32'sd0.0657721899757848, 32'sd-0.12010144896844878, 32'sd-0.09723450668739157, 32'sd0.0093127782366951, 32'sd-0.11403422053508067, 32'sd-0.011786502875602043, 32'sd0.07855739204299717, 32'sd-0.11079464959870726, 32'sd0.013883887204042584, 32'sd0.048504218281674116, 32'sd0.0060937012912219155, 32'sd0.06899956422833545, 32'sd-0.051902587214186745, 32'sd0.06780205068471055, 32'sd-0.0014391718653736897, 32'sd0.07897784637918082, 32'sd0.016119423740973336, 32'sd-0.019956217078261708, 32'sd-0.040447235843817854, 32'sd1.5119951975631762e-120, 32'sd1.8171400440320475e-123, 32'sd0.04057430818195146, 32'sd-0.09884296343543329, 32'sd-0.04267128654245134, 32'sd-0.029864579734872852, 32'sd0.06328726804130565, 32'sd-0.008082863551095866, 32'sd-0.014760956925877597, 32'sd-0.1770084536718103, 32'sd-0.16718501575637423, 32'sd-0.17446705324550812, 32'sd-0.03332712298950541, 32'sd-0.046332824637527276, 32'sd-0.01122086948161714, 32'sd0.07484100280953351, 32'sd0.05676780974675677, 32'sd0.09976736249514762, 32'sd0.11219276123772964, 32'sd0.09388039110666549, 32'sd-0.02193676445136498, 32'sd0.020427225362230884, 32'sd0.09556426370363337, 32'sd-0.03841156841400788, 32'sd-0.0006106698903737165, 32'sd-0.04602081557136393, 32'sd-0.028901447256147406, 32'sd0.020809144139471998, 32'sd-0.029939105132368384, 32'sd3.6737248556406426e-123, 32'sd-0.06008560707925292, 32'sd0.0833736122857579, 32'sd0.0045807432746922064, 32'sd-0.084313133739253, 32'sd-0.07773942247905982, 32'sd-0.10408085191900517, 32'sd-0.20163347416827276, 32'sd-0.12770353468558301, 32'sd-0.08637525128649554, 32'sd-0.11280458618596752, 32'sd0.0595547977707677, 32'sd0.013941189966257258, 32'sd-0.12031219479324623, 32'sd-0.09141944782848292, 32'sd-0.04609406120968969, 32'sd-0.025522101133337464, 32'sd0.0070471452568503816, 32'sd0.05129868714239808, 32'sd0.12488014742466272, 32'sd-0.003040059262163063, 32'sd-0.106896217277345, 32'sd-0.09903349274863535, 32'sd-0.09167216062610205, 32'sd-0.05944601992201127, 32'sd-0.031137531469751217, 32'sd-0.03137419539709855, 32'sd0.015667117839757546, 32'sd-7.162755792105449e-115, 32'sd-0.05861382476582555, 32'sd0.03344839526569534, 32'sd0.014229905647811607, 32'sd-0.0930114247086318, 32'sd-0.12477591294381608, 32'sd-0.09004519763712526, 32'sd-0.10091310607395243, 32'sd-0.1801718750111721, 32'sd-0.1298476784503692, 32'sd-0.018280547392905334, 32'sd-0.056769589786756815, 32'sd-0.09386097217841613, 32'sd0.028807842062704946, 32'sd0.14518633359871186, 32'sd0.1519221039472956, 32'sd0.018162304303644374, 32'sd0.03544692312272678, 32'sd0.09339760714195061, 32'sd0.11039294864648146, 32'sd0.12351754971354147, 32'sd0.028050464996590002, 32'sd-0.1258122445785087, 32'sd-0.10755548502846199, 32'sd-0.11718081832558454, 32'sd0.058766911622146874, 32'sd-0.03335019589890461, 32'sd0.0505162054062296, 32'sd-0.021942778535134846, 32'sd-0.07083447548847885, 32'sd-0.003564252570538471, 32'sd0.007483249502340379, 32'sd-0.015881306912777508, 32'sd-0.1657433200951073, 32'sd-0.22066142697814622, 32'sd-0.1804820692529336, 32'sd-0.22213215473337083, 32'sd-0.1718157215708206, 32'sd0.056426598814496166, 32'sd-0.046015458812188575, 32'sd-0.002930880265127431, 32'sd0.07331787400714261, 32'sd0.14676078615636656, 32'sd0.14178653796347554, 32'sd-0.01240040403813126, 32'sd-0.06976698051534141, 32'sd0.03925889105294501, 32'sd-0.027318251486781256, 32'sd0.13608340452485496, 32'sd0.14981660191557863, 32'sd-0.038028448010611254, 32'sd-0.1320640164939147, 32'sd0.019433749506466317, 32'sd0.014051825573150791, 32'sd-0.031543983945989805, 32'sd-0.0689616348719105, 32'sd-0.027609923900512087, 32'sd0.036889809922020136, 32'sd0.10095341298206204, 32'sd0.003414120432145754, 32'sd-0.1250835605190255, 32'sd-0.24973268772307206, 32'sd-0.15739737251399383, 32'sd-0.17456810589350943, 32'sd-0.1396815835979406, 32'sd-0.1137263778424046, 32'sd0.02183118856363413, 32'sd0.13274908999250062, 32'sd0.053052663554605924, 32'sd0.17640828536347988, 32'sd0.04471715913678101, 32'sd0.028397335085225774, 32'sd0.04018188529051507, 32'sd-0.04545493522087295, 32'sd-0.0012167317069543676, 32'sd-0.016663135289950715, 32'sd-0.0774807204328341, 32'sd0.09020293210905996, 32'sd-0.10696303227447755, 32'sd-0.10586551253722197, 32'sd0.04491722446704646, 32'sd-0.06987016864953789, 32'sd-0.014477172521799558, 32'sd-0.07191386273758155, 32'sd-0.05894008777455661, 32'sd-0.10077186881072334, 32'sd0.02991701086030191, 32'sd0.06442829422783462, 32'sd-0.1592087061150123, 32'sd-0.1644191065368439, 32'sd-0.2115190109111699, 32'sd-0.22829250418166655, 32'sd-0.11499688105705479, 32'sd0.04958659780406257, 32'sd0.16727272156935175, 32'sd0.0038143979836733704, 32'sd0.03415092782754814, 32'sd0.14559703365389892, 32'sd0.10094182777033867, 32'sd0.03158694324074148, 32'sd0.00896833919054645, 32'sd-0.209518034229316, 32'sd-0.07875802833742382, 32'sd-0.10836959058532514, 32'sd-0.04547452302918498, 32'sd-0.111969774636336, 32'sd0.0037585882565959712, 32'sd0.04025849523973152, 32'sd0.04703347629210655, 32'sd7.137210921388549e-05, 32'sd-0.0668056012863774, 32'sd-0.10007352292907921, 32'sd0.02280312473256829, 32'sd-0.0833473576860096, 32'sd0.061376453909448424, 32'sd0.0024751934770543284, 32'sd-0.1626157757502097, 32'sd-0.1747346303744461, 32'sd-0.1407185848351909, 32'sd0.0018612837226632754, 32'sd-0.04387903460763643, 32'sd0.03869555010254933, 32'sd0.043487756907477575, 32'sd-0.02072491950863615, 32'sd-0.06652831187647627, 32'sd0.016716285109094373, 32'sd0.15594388892192906, 32'sd-0.07018337056414767, 32'sd-0.09246095635636407, 32'sd-0.11159298085048536, 32'sd-0.12921260644365257, 32'sd-0.2129577637831899, 32'sd-0.012128958304289377, 32'sd-0.06288689841060092, 32'sd-0.0981872966632489, 32'sd0.04701089204321216, 32'sd0.055225569949724516, 32'sd-0.018435076342081337, 32'sd-0.06585350255532456, 32'sd-0.05356973708160637, 32'sd-0.056269378217737205, 32'sd-0.11528984777550251, 32'sd-0.0565108275982899, 32'sd-0.032153750866910934, 32'sd-0.1610712343292837, 32'sd-0.10381340325037884, 32'sd-0.2138033395992837, 32'sd0.06754001793532205, 32'sd0.07844002545930673, 32'sd0.16213282222727401, 32'sd0.018520344301569788, 32'sd-0.09023119964226405, 32'sd0.024262245291288276, 32'sd0.13092892803096337, 32'sd-0.0005204317872167086, 32'sd-0.13050100185150854, 32'sd-0.29748047080230844, 32'sd-0.24195634618870424, 32'sd0.0011566440227483122, 32'sd-0.16474312619770556, 32'sd-0.02785165648184517, 32'sd-0.027446835058578145, 32'sd-0.02253287245972766, 32'sd-0.020417654830960762, 32'sd0.06913655725511203, 32'sd0.11326137802238753, 32'sd0.025159608390362503, 32'sd-0.06648957819642264, 32'sd0.005208780330034928, 32'sd-0.028705036554884714, 32'sd-0.13323130706210895, 32'sd0.019567190911316507, 32'sd-0.07176197441089348, 32'sd-0.20604461701261345, 32'sd-0.18330723257877832, 32'sd-0.005748783053077257, 32'sd0.11733057754247955, 32'sd0.02013724382710333, 32'sd-0.06264164178225905, 32'sd0.08366187216429066, 32'sd0.06183666537817829, 32'sd-0.011375692409814626, 32'sd-0.06804153748405405, 32'sd-0.29382459016569246, 32'sd-0.11950052884574101, 32'sd-0.128605682180841, 32'sd-0.06368255909901889, 32'sd0.01179545858299892, 32'sd0.09144914035205835, 32'sd0.12082296899804955, 32'sd0.035778112784190456, 32'sd0.15752201961052545, 32'sd0.11017294054275736, 32'sd-0.0007559405036220171, 32'sd0.0390301920408766, 32'sd-0.07142306360522023, 32'sd-0.01164139932702576, 32'sd-0.07149244038529991, 32'sd-0.08432461517715747, 32'sd0.014114316614393014, 32'sd-0.05528182462015085, 32'sd-0.1283963616210748, 32'sd0.05141675648959221, 32'sd0.027562364736329434, 32'sd0.10134647049813185, 32'sd-0.026792078895309386, 32'sd0.0050017125597551755, 32'sd0.0680907062077444, 32'sd0.04970119994311614, 32'sd-0.049605708315767424, 32'sd-0.11938650202643858, 32'sd-0.04133222178514429, 32'sd0.07285844351110576, 32'sd0.003382793067135386, 32'sd0.010157546347242679, 32'sd0.16569422331929867, 32'sd0.10794961063980496, 32'sd0.013785421012777748, 32'sd0.1976752119152667, 32'sd0.10916079355712623, 32'sd-0.03958753050970535, 32'sd-0.1223430251237259, 32'sd-0.013737765615331965, 32'sd-0.06785903332069636, 32'sd-0.03314891304997747, 32'sd-0.03486288773919331, 32'sd0.020228191481021056, 32'sd-0.04872314283326647, 32'sd-0.07327113740277354, 32'sd0.02056921725419266, 32'sd0.033921644937628025, 32'sd-0.0032869265975716123, 32'sd0.001488146281466577, 32'sd0.005497624258283998, 32'sd-0.04458412587819832, 32'sd-0.07173832984421961, 32'sd-0.12509413414790496, 32'sd-0.0963068989951948, 32'sd0.013383945186075432, 32'sd-0.03423055021493784, 32'sd0.18317409858225583, 32'sd0.04292251408398292, 32'sd0.02160778403944496, 32'sd0.102005391882202, 32'sd0.08631226529976348, 32'sd0.07724819118365989, 32'sd0.09048456528526999, 32'sd-0.027300024109365363, 32'sd-0.05547773391612979, 32'sd-0.015909513583103677, 32'sd0.017271549978652302, 32'sd0.022705046139663093, 32'sd-0.04370672961151314, 32'sd0.005233816999338945, 32'sd0.06359500362367856, 32'sd-0.08447471516426368, 32'sd-0.14374706715242555, 32'sd-0.01620614842663926, 32'sd-0.017541978446954744, 32'sd0.12761106194038718, 32'sd0.15618691526764714, 32'sd-0.049746453134922285, 32'sd0.06576325948969526, 32'sd-0.0858177092016193, 32'sd-0.06576680233271447, 32'sd-0.016727712044776983, 32'sd0.00476376838253486, 32'sd0.018167640352375183, 32'sd0.09659070715665626, 32'sd0.0024050046779686314, 32'sd-0.0324639066798929, 32'sd0.04486319571363053, 32'sd0.047270016978911214, 32'sd-0.09093325972198306, 32'sd0.014655660433627168, 32'sd-0.03081146507859059, 32'sd-0.08292368113720182, 32'sd0.03771124004713496, 32'sd-0.04132415058321274, 32'sd0.029869231271429604, 32'sd0.004325143129205073, 32'sd0.0279800534681822, 32'sd0.0136527290901451, 32'sd-0.07351263607052426, 32'sd-0.13975223151882293, 32'sd-0.046743240526300016, 32'sd-0.05861352695096517, 32'sd0.1450621542930979, 32'sd0.14251572761598477, 32'sd-0.021943834971263603, 32'sd-0.02408851380561291, 32'sd0.06116656171282716, 32'sd-0.07160229453085842, 32'sd-0.018789730459095155, 32'sd-0.03459432747997974, 32'sd0.04329490293648599, 32'sd-0.016219007867667997, 32'sd-0.037844007649949704, 32'sd-0.013731157092543439, 32'sd-0.0033393345049631817, 32'sd0.09359222329611915, 32'sd0.005344207202774697, 32'sd-0.10596675791778576, 32'sd0.05264423357320004, 32'sd-0.04571384807487076, 32'sd0.08642682984550192, 32'sd0.05289108246861524, 32'sd0.023444373451173946, 32'sd1.0141939276648058e-115, 32'sd-0.06581273506468076, 32'sd-0.006670232003388025, 32'sd0.028928713968320842, 32'sd0.01545469872096832, 32'sd-0.002224596637415445, 32'sd0.07216490280456633, 32'sd0.020582221357902296, 32'sd0.01133075908896164, 32'sd-0.007033553059096129, 32'sd-0.10190684813687607, 32'sd-0.11234167667861311, 32'sd0.04171038782067048, 32'sd-0.023745000414495013, 32'sd0.04152485854557286, 32'sd-0.11501200570957888, 32'sd-0.06676771835161835, 32'sd0.06322344741556568, 32'sd-0.050982204004016395, 32'sd-0.08344683566134109, 32'sd0.08360005787909493, 32'sd0.05713794153749163, 32'sd0.06241631330497463, 32'sd-0.037483415683513176, 32'sd0.007271273136855601, 32'sd-0.14168231915315818, 32'sd-0.018344234439212594, 32'sd0.05603063584930102, 32'sd-0.025487125520168793, 32'sd-0.06322020520646592, 32'sd0.021589818277173944, 32'sd0.0463409708768358, 32'sd-0.11477496005213951, 32'sd-0.04518544011552167, 32'sd-0.10050907506407722, 32'sd0.11223438432610904, 32'sd0.14797193318112753, 32'sd0.11268127972011813, 32'sd-0.004878601869838399, 32'sd-0.09992417220153303, 32'sd0.06324808619528603, 32'sd0.04888381543637905, 32'sd-0.035863097342186956, 32'sd-0.10122223870925201, 32'sd-0.037077799899923644, 32'sd0.1378108913911326, 32'sd-0.0915515824811351, 32'sd-0.014045730120577807, 32'sd0.02748089797706546, 32'sd0.06778910030328072, 32'sd0.050121373083680865, 32'sd0.06921333297879902, 32'sd-0.004816959895843779, 32'sd0.03040052425003151, 32'sd-0.035284850741260886, 32'sd0.009191734798274724, 32'sd-0.038097597634565654, 32'sd-0.0018789142643679344, 32'sd-0.05135325216873625, 32'sd-0.0801811925898668, 32'sd-0.06140781143578006, 32'sd0.01928833521023894, 32'sd-0.05352057235996562, 32'sd0.14725670421789686, 32'sd0.21321549421997402, 32'sd0.1288122641921939, 32'sd0.1388201792017039, 32'sd0.01295628594071469, 32'sd-0.059286711793397055, 32'sd-0.0015844056125625713, 32'sd-0.01584578216069348, 32'sd-0.0756059171041741, 32'sd-0.1010821994411126, 32'sd-0.026139233780749907, 32'sd0.013748387454228362, 32'sd-0.06531742557971043, 32'sd-0.06832518841107346, 32'sd0.17772721623680682, 32'sd0.2444704097123498, 32'sd0.20347584435097194, 32'sd-0.005832050262029244, 32'sd-0.12318578930190847, 32'sd-0.02343114558687784, 32'sd0.040289941370328784, 32'sd-1.3193040677589894e-118, 32'sd-0.05292593859345442, 32'sd-0.03969749107594328, 32'sd-0.04121483252737322, 32'sd-0.08624518419588059, 32'sd0.09458210187460146, 32'sd-0.003862921245413953, 32'sd0.00847596574868973, 32'sd0.05488954324834683, 32'sd0.21642669687349528, 32'sd0.23128206147821054, 32'sd0.04593049127324458, 32'sd-0.06483209258685611, 32'sd0.041300265542927886, 32'sd-0.058096599634123086, 32'sd-0.033199053353096517, 32'sd-0.06172333528230154, 32'sd0.05401867979322128, 32'sd-0.05575345669313226, 32'sd-0.04263576571415864, 32'sd0.12657963799109895, 32'sd0.14906667007160196, 32'sd0.14021114730573286, 32'sd0.10099888974514307, 32'sd-0.04406668686576013, 32'sd0.0064408436227037826, 32'sd0.07719839012587852, 32'sd-0.03378141029016274, 32'sd-0.0016390415239128122, 32'sd0.01582362004378848, 32'sd0.05623726744445043, 32'sd-0.028388265071683072, 32'sd0.010416112496853664, 32'sd-0.05644596199989265, 32'sd-0.06917755530642065, 32'sd0.03494783755465101, 32'sd0.003106718312731442, 32'sd0.11825056689896175, 32'sd0.1414386323510271, 32'sd0.04608356123892311, 32'sd0.043633750404927646, 32'sd0.15828145247035696, 32'sd0.0012137520071267957, 32'sd0.0027088616997223017, 32'sd-0.01661625865135564, 32'sd-0.008317169954525465, 32'sd-0.028835786739837787, 32'sd-0.024222302703242337, 32'sd0.12820954151434993, 32'sd0.052531848413076794, 32'sd-0.0062095465969874575, 32'sd0.1104147638698287, 32'sd0.09705388628620705, 32'sd-0.10118393684813042, 32'sd0.0245430913461192, 32'sd-0.05637561746441089, 32'sd-0.030558063058466964, 32'sd-0.02995105462673955, 32'sd-0.06680378862883987, 32'sd0.11071669170158938, 32'sd0.0932363769387335, 32'sd0.016142839374826218, 32'sd0.021433494775232344, 32'sd0.02130202812566836, 32'sd-0.03320111112865068, 32'sd-0.06450950748923105, 32'sd-0.04196460910038142, 32'sd-0.11444129243519653, 32'sd0.12140827626868812, 32'sd0.1487900527937925, 32'sd0.13820418513902627, 32'sd0.18833478267616377, 32'sd-0.00916353055150129, 32'sd-0.09620151024052702, 32'sd-0.02732970568137918, 32'sd0.012119595788302887, 32'sd-0.05986676030676254, 32'sd0.09234184010525413, 32'sd-0.06492184928972164, 32'sd0.06616668343198538, 32'sd0.057731931211861855, 32'sd-0.016816895915236434, 32'sd0.1021855331249353, 32'sd0.0069779454317323835, 32'sd1.0456204504638936e-120, 32'sd-0.003435370433709804, 32'sd0.06610606357837248, 32'sd0.022347373984775525, 32'sd0.0316998193023969, 32'sd0.19684848917000242, 32'sd0.018254198394699724, 32'sd-0.05232475876781967, 32'sd-0.053849320667135256, 32'sd-0.17609330542582421, 32'sd-0.09376855655155757, 32'sd-0.11067340164249677, 32'sd0.011267829903812254, 32'sd0.07427662570593264, 32'sd0.03680039153585611, 32'sd0.13677655021154658, 32'sd0.08014173808325427, 32'sd0.10148995518163459, 32'sd0.09539505694856655, 32'sd-0.014267409569999761, 32'sd-0.031319329716820984, 32'sd-0.13607309107109034, 32'sd-0.019549304360009345, 32'sd-0.032059526673770655, 32'sd0.043021902226417115, 32'sd0.00391000576610183, 32'sd0.028743209992572693, 32'sd2.338733765826409e-120, 32'sd2.4794707532549398e-126, 32'sd-1.4333851540779728e-117, 32'sd-0.02878901130751367, 32'sd-0.11845690334286237, 32'sd0.01118080043974236, 32'sd0.08060938867783986, 32'sd-0.07839931157567936, 32'sd-0.015596228666576655, 32'sd-0.05750223098355966, 32'sd-0.08182754568836127, 32'sd0.054428185024841265, 32'sd-0.04777811494521329, 32'sd-0.039396955197171825, 32'sd-0.139035276192792, 32'sd-0.08587578170969092, 32'sd-0.01452898962796075, 32'sd0.09533852931548477, 32'sd-0.01813129793740469, 32'sd-0.11521822760470993, 32'sd-0.10867363028716857, 32'sd-0.13972046748557268, 32'sd-0.1580015292026124, 32'sd0.009164319737939328, 32'sd0.08171738554105676, 32'sd-0.04202747206082648, 32'sd0.009843402486757368, 32'sd-0.03666418031959869, 32'sd-1.211104937260233e-114, 32'sd-1.5825936139360215e-115, 32'sd-3.511548412777491e-119, 32'sd0.06400525322037429, 32'sd-0.06470981697668765, 32'sd-0.10496193152031821, 32'sd0.06699764508363992, 32'sd-0.06946596474536317, 32'sd-0.15351237396118741, 32'sd0.030766205851220436, 32'sd0.05423418307374405, 32'sd-0.027283059843301396, 32'sd0.05436810610723034, 32'sd-0.006658531013133548, 32'sd-0.014771483893533255, 32'sd-0.0958591598675609, 32'sd0.01672583315017712, 32'sd0.06143415175150842, 32'sd0.06704105735569628, 32'sd-0.1187499169467913, 32'sd0.040257600776759266, 32'sd0.05323979386458725, 32'sd-0.06559427468027575, 32'sd-0.056869211211489655, 32'sd0.05588215188692007, 32'sd-0.013977716851183587, 32'sd-0.04953835129057416, 32'sd-0.052268782984548304, 32'sd-4.7639468623634904e-120, 32'sd6.510777764903799e-115, 32'sd5.285592043147753e-118, 32'sd-3.702780690860637e-123, 32'sd-0.02569308908378357, 32'sd-0.05089333741262306, 32'sd-0.1244958487767677, 32'sd-0.031127890140402778, 32'sd0.006614657991731609, 32'sd-0.0563725277679526, 32'sd-0.11568025412496231, 32'sd0.012577321057076018, 32'sd0.041684306621781055, 32'sd-0.09060956972538538, 32'sd-0.19516419348913752, 32'sd-0.1797514559826115, 32'sd-0.15474791441250726, 32'sd-0.06292299935515826, 32'sd-0.14112392485857672, 32'sd0.025306200288899988, 32'sd-0.05145360425067814, 32'sd0.04325604034369711, 32'sd0.05964948775335004, 32'sd-0.1052743454211863, 32'sd0.05668715085274279, 32'sd-0.034675022802918086, 32'sd-0.020209557060211828, 32'sd7.560659805171209e-115, 32'sd-1.3097791906514583e-118, 32'sd-2.5450130105481833e-124, 32'sd-1.598297826050344e-126, 32'sd2.5638914373217896e-124, 32'sd5.242104361035733e-116, 32'sd-0.0010445019202580373, 32'sd0.021096247465389687, 32'sd0.037976841298251934, 32'sd-0.004220509791578899, 32'sd-0.07074967674227316, 32'sd0.017479849285736825, 32'sd-0.08419734450854674, 32'sd-0.11634312267655597, 32'sd-0.05485848503826219, 32'sd-0.06212155560217934, 32'sd0.05444628574612398, 32'sd0.06141922282928376, 32'sd-0.017911648118865055, 32'sd0.06211895014820934, 32'sd-0.06575412242948196, 32'sd-0.04160031312624241, 32'sd-0.06986940812736137, 32'sd-0.04220434119521487, 32'sd0.006966556777457378, 32'sd0.04470338049286142, 32'sd2.574822566774599e-124, 32'sd-3.248298676688146e-122, 32'sd3.0125149601348057e-123, 32'sd3.374560171045072e-115},
        '{32'sd-3.424868523179919e-117, 32'sd-3.3833116007844834e-120, 32'sd-6.469423611128426e-123, 32'sd-1.0507749588962546e-125, 32'sd3.466699848569813e-119, 32'sd1.1620744518161175e-114, 32'sd1.1531760544870538e-125, 32'sd-1.3191433539831598e-123, 32'sd-6.214490891299311e-126, 32'sd1.0757318940374375e-124, 32'sd-3.737100487391129e-122, 32'sd-7.921157770342681e-115, 32'sd0.07834146171739868, 32'sd0.029452175419769917, 32'sd0.052956783490310994, 32'sd0.09170220755847812, 32'sd4.790796164905676e-130, 32'sd-6.438608334405643e-124, 32'sd-9.686046634515383e-122, 32'sd1.4005683504601299e-117, 32'sd1.02514140664105e-118, 32'sd-8.679399103598564e-122, 32'sd-5.615118485702354e-126, 32'sd-3.8218492510183057e-119, 32'sd-7.6036893258053e-118, 32'sd-4.744137692600798e-115, 32'sd-6.479527707080239e-121, 32'sd-2.4710078370416546e-121, 32'sd-9.339030000871872e-126, 32'sd-2.5679953637529102e-123, 32'sd8.977227310689547e-123, 32'sd1.8061628696016846e-127, 32'sd0.098450325514622, 32'sd0.06772175376593374, 32'sd0.06490161415521455, 32'sd0.07072565899450571, 32'sd0.11503621318401587, 32'sd0.05453380028271632, 32'sd0.1986725380063926, 32'sd0.13352386367958405, 32'sd0.10833906209656732, 32'sd0.02778109355051676, 32'sd-0.02651611895751412, 32'sd0.017909862731089826, 32'sd0.06514890912185925, 32'sd0.07431596706940616, 32'sd0.11335040621795972, 32'sd0.005132970817307831, 32'sd0.08724530234280937, 32'sd0.07919753322851163, 32'sd0.12922530003473454, 32'sd0.09268590517725052, 32'sd-1.8155383710462946e-123, 32'sd1.4750117205507934e-123, 32'sd-2.4674179284161885e-121, 32'sd-4.102663039326335e-126, 32'sd1.165981670561735e-122, 32'sd1.238604418047026e-122, 32'sd0.06522085089366723, 32'sd0.07237222970687272, 32'sd-0.04581967256082397, 32'sd0.08167802221311249, 32'sd-0.01932471632594092, 32'sd0.0031753975836447705, 32'sd-0.039188474153521204, 32'sd-0.040029018553426665, 32'sd0.028487450353344757, 32'sd0.05805817332606131, 32'sd0.10763719553857953, 32'sd-0.05873310376120825, 32'sd0.0651666711116942, 32'sd0.11971358381377134, 32'sd0.1286956669637287, 32'sd0.05749078633856373, 32'sd0.13094153861837107, 32'sd-0.002529655539308355, 32'sd0.03423104803545189, 32'sd0.08278760092744193, 32'sd0.049104824091271496, 32'sd0.09002801619023834, 32'sd0.10112828756327848, 32'sd0.08668805013025783, 32'sd-1.4767410546879101e-125, 32'sd-3.9240809113707082e-115, 32'sd9.56019034236689e-125, 32'sd3.5943863899094556e-125, 32'sd0.09683237356010889, 32'sd0.0730776697670832, 32'sd0.01334019330516688, 32'sd0.10096759411005495, 32'sd0.045410338243863015, 32'sd0.07948209339643385, 32'sd0.0075301125642045184, 32'sd0.09792188895301754, 32'sd0.03045440430479686, 32'sd-0.04233691456170781, 32'sd-0.009831743367136212, 32'sd-0.02660950426268752, 32'sd-0.02255839872641502, 32'sd0.0973151139970923, 32'sd0.0027242121352913035, 32'sd-0.010538956284983457, 32'sd0.013119348733977928, 32'sd-0.0506652975828294, 32'sd0.09991484530249704, 32'sd0.08551003891278042, 32'sd-0.028539294317056433, 32'sd0.013360686557070798, 32'sd0.003264192764145227, 32'sd0.02194408794769567, 32'sd-0.03599769865045855, 32'sd1.1793476006326022e-122, 32'sd-7.171414940509419e-121, 32'sd0.07789998501571936, 32'sd-0.027286056160484292, 32'sd0.03857899834721367, 32'sd-0.030969640927603737, 32'sd0.01767430171070569, 32'sd0.08849864845561944, 32'sd0.07505465973958358, 32'sd0.09930168906394318, 32'sd0.04210198692170381, 32'sd0.09114422761326005, 32'sd0.05225004449029601, 32'sd0.024740266259645323, 32'sd0.010101029364531345, 32'sd0.04128702374240883, 32'sd0.011283858823813778, 32'sd0.09804202546536306, 32'sd-0.0769863117912253, 32'sd0.056911179275090505, 32'sd-0.06433277279164207, 32'sd0.026766131712604422, 32'sd0.06435343436930496, 32'sd-0.02570123151970788, 32'sd-0.08905788263914337, 32'sd-0.03622646762933337, 32'sd0.0655558665295381, 32'sd-0.0152866450873612, 32'sd-0.014584248274508002, 32'sd1.4557222177073595e-122, 32'sd0.03435947965167901, 32'sd0.023388352621879504, 32'sd0.07197070107166129, 32'sd0.0526401060269076, 32'sd0.12631827748741853, 32'sd-0.030332526937635083, 32'sd0.057245744135405945, 32'sd0.041309553600931026, 32'sd0.0234339918954208, 32'sd0.07970334670507924, 32'sd0.08797394910574471, 32'sd-0.050666988681904744, 32'sd0.037067780758896475, 32'sd-0.0373433248363809, 32'sd-0.0924116434276852, 32'sd-0.087078184424455, 32'sd-0.08879698752340867, 32'sd0.10613730951658229, 32'sd0.008760095395138742, 32'sd0.06292341439197155, 32'sd0.08239107872026423, 32'sd0.08577678942420719, 32'sd-0.07692555623515171, 32'sd-0.06091814692642432, 32'sd0.0625056323091043, 32'sd0.012703748789921865, 32'sd0.0693249451613563, 32'sd3.3238263991694027e-116, 32'sd0.0056423459582095915, 32'sd-0.002081209146679315, 32'sd0.07475689339355718, 32'sd0.004733203308345787, 32'sd0.14161004622292206, 32'sd0.08610019430115817, 32'sd0.10452244912491154, 32'sd0.03413116517096126, 32'sd-0.053850426081052186, 32'sd-0.0018941650911079558, 32'sd0.04725895704967715, 32'sd0.08140094861828515, 32'sd-0.011898099629546044, 32'sd0.01138701891333043, 32'sd-0.064725882900087, 32'sd-0.12324356548428521, 32'sd-0.018294525257988112, 32'sd0.08381855143875502, 32'sd-0.00035967712889034087, 32'sd0.06950565275995034, 32'sd0.007041950136173089, 32'sd0.05371515082105565, 32'sd-0.031737322677625135, 32'sd0.11913401245051695, 32'sd0.11274226662539817, 32'sd0.06554629824163738, 32'sd0.02324630805604517, 32'sd0.07864061925072445, 32'sd0.07003611567744603, 32'sd0.014921413645552432, 32'sd-0.018975211871425757, 32'sd0.07250290667482442, 32'sd0.08936435339073766, 32'sd0.08680339264136756, 32'sd0.05630238214164134, 32'sd0.053221732152037515, 32'sd0.003040450051585909, 32'sd0.1134180347507873, 32'sd0.07601976421653536, 32'sd0.11156520945374736, 32'sd0.03789988175647933, 32'sd0.09701878755562432, 32'sd-0.02920244289081127, 32'sd0.014916571922221714, 32'sd0.07400567271716939, 32'sd-0.0019217204038142642, 32'sd0.06166619267075309, 32'sd0.22985685717814955, 32'sd0.13432968549885518, 32'sd0.10262554437365111, 32'sd-0.0063976697462379654, 32'sd-0.0025377879342241088, 32'sd-0.007721810779773635, 32'sd-0.004397600038859964, 32'sd-0.021288316560544904, 32'sd0.08856514123404671, 32'sd-0.014857748915046813, 32'sd0.010013022136896144, 32'sd0.05603431628458596, 32'sd-0.09500617391385333, 32'sd0.01291029506714588, 32'sd-0.07123802958047319, 32'sd0.046474592158705655, 32'sd-0.004506890369239329, 32'sd0.08933296419073002, 32'sd0.01639819040201409, 32'sd0.0014418093322811792, 32'sd0.13066036651199003, 32'sd0.09005080972555637, 32'sd0.0017708440484611814, 32'sd0.09675835008376524, 32'sd-0.04313646034315063, 32'sd-0.0873052971273043, 32'sd-0.069004594102765, 32'sd-0.0654961952051309, 32'sd0.047255888644280215, 32'sd0.01984170266668061, 32'sd0.09124898729576397, 32'sd-0.07775688359270895, 32'sd0.09031671632329157, 32'sd-0.07727935940353332, 32'sd0.04966321055698077, 32'sd0.06965828940210407, 32'sd0.0022594768058184587, 32'sd-0.020424493381485342, 32'sd0.08553080623059638, 32'sd-0.03966832711384506, 32'sd0.02455757179370394, 32'sd0.05562377807923611, 32'sd0.018377454379700033, 32'sd0.06186604046876372, 32'sd-0.006010356043775253, 32'sd0.11535061953005676, 32'sd0.13107757546400253, 32'sd0.0005656594509739721, 32'sd0.06248470223187377, 32'sd0.08615928559424303, 32'sd0.10233189819271951, 32'sd0.06829290833354262, 32'sd-0.06389177613930508, 32'sd-0.14765613912529127, 32'sd-0.02984732306567297, 32'sd-0.11018244496056236, 32'sd-0.04534885635559603, 32'sd-0.05706052677723152, 32'sd-0.013303446499170883, 32'sd0.012196988044458528, 32'sd0.04314260655006358, 32'sd-0.039773133891917924, 32'sd-0.0480318825493927, 32'sd-0.00313491645359077, 32'sd-0.023106210840086017, 32'sd0.013539286665075105, 32'sd0.003664263769544769, 32'sd-0.07245584032776753, 32'sd-0.11885528452078915, 32'sd-0.1403519656813572, 32'sd0.06128514366984794, 32'sd0.013002298985047848, 32'sd-0.0009182524688577119, 32'sd0.0696703953177964, 32'sd0.12294842855838777, 32'sd0.005409279463673661, 32'sd-0.06001246077102858, 32'sd0.06518874455683657, 32'sd-0.0036105188031593763, 32'sd-0.03800072172736204, 32'sd-0.14201471100410898, 32'sd-0.06439675876945344, 32'sd-0.008190171649187027, 32'sd-0.17090493392205516, 32'sd-0.15876795480844746, 32'sd-0.02020267235253965, 32'sd-0.09310525338732055, 32'sd-0.16157107342775517, 32'sd-0.11704324777420128, 32'sd-0.050678671913114294, 32'sd-0.049840872500151526, 32'sd-0.03381074722530779, 32'sd0.029419280005144606, 32'sd-0.0329010448802294, 32'sd-0.036918502718772304, 32'sd-0.04243956768279945, 32'sd0.05266972357078159, 32'sd-0.006149835882314463, 32'sd-0.0975394680653387, 32'sd-0.009773982424453657, 32'sd0.018697422417098587, 32'sd-0.018633735317872203, 32'sd-0.08464054463943575, 32'sd-0.19482895073336468, 32'sd-0.13691863394420462, 32'sd-0.08340412779628775, 32'sd-0.017817017383636266, 32'sd-0.1479078958337616, 32'sd-0.1915278601596366, 32'sd-0.06792572599003932, 32'sd-0.0011115919550495953, 32'sd-0.1330486675069847, 32'sd-0.20543376101216423, 32'sd-0.16177786906471842, 32'sd-0.12478171986303697, 32'sd0.0451648374827079, 32'sd0.10544960946722134, 32'sd0.007829008984726117, 32'sd0.13903288992650353, 32'sd-0.05275597065198114, 32'sd0.07506313539200832, 32'sd0.04646253496682417, 32'sd0.0667004921114437, 32'sd0.04076276430451143, 32'sd-0.02634247719354323, 32'sd-0.0934927257346033, 32'sd0.00011007119357275174, 32'sd0.004218872216042667, 32'sd0.017015262049479098, 32'sd0.07790140159462938, 32'sd-0.13090543353152187, 32'sd-0.12374129190923264, 32'sd-0.020146416561182667, 32'sd-0.0761173529445364, 32'sd-0.020404395453697308, 32'sd-0.2093047163898071, 32'sd-0.0362827783541148, 32'sd0.003076638894792323, 32'sd0.035128495448398835, 32'sd-0.05093593349376626, 32'sd0.03233545772869132, 32'sd-0.06498317493022802, 32'sd-0.2126006411550669, 32'sd0.05644435782616159, 32'sd-0.014547334631288038, 32'sd0.08143350724579632, 32'sd0.1369761590156121, 32'sd-0.06444233383078798, 32'sd-0.011313581200341392, 32'sd0.012104234490949297, 32'sd0.04089502238187358, 32'sd0.006003862677819899, 32'sd-0.0829645372586673, 32'sd0.006915273797322443, 32'sd-0.020315239875430036, 32'sd0.08804038959052074, 32'sd0.12549741595951155, 32'sd-0.07986462016191193, 32'sd-0.12690456376517667, 32'sd-0.11528607638281023, 32'sd-0.13942455550249833, 32'sd-0.004347343691037821, 32'sd0.011584282356555191, 32'sd-0.1585559599895115, 32'sd-0.1699901924110933, 32'sd-0.07651078421286925, 32'sd-0.07537239435611323, 32'sd0.04114491762815459, 32'sd-0.06697031888057697, 32'sd-0.0470745842409278, 32'sd-0.16267341802902255, 32'sd-0.0805980183182128, 32'sd-0.010765079464274746, 32'sd0.011119531405117804, 32'sd-0.01726651673459239, 32'sd0.06069886734183988, 32'sd0.0800870367869694, 32'sd0.06231697360367359, 32'sd0.0030338232978645795, 32'sd0.03674714628773772, 32'sd0.010647577612627612, 32'sd-0.009803542613704936, 32'sd0.08765526012607905, 32'sd0.15315801427321293, 32'sd0.015465538917139943, 32'sd-0.03734061964690875, 32'sd-0.1400652253935274, 32'sd-0.14989320403242973, 32'sd-0.12756957558569398, 32'sd-0.028246107023252864, 32'sd0.09313096726905189, 32'sd-0.022077773751380102, 32'sd-0.1527865922399851, 32'sd-0.1984100586931966, 32'sd-0.07722204054971037, 32'sd-0.14390453389079824, 32'sd0.01747719779586003, 32'sd-0.04200942548306798, 32'sd0.003812571881619427, 32'sd0.09108317623832855, 32'sd-0.016843466772323516, 32'sd-0.008140278140685898, 32'sd-0.01228594815445835, 32'sd-0.02570622491223993, 32'sd0.02539313362423349, 32'sd-0.029576205757402243, 32'sd0.16286672816976291, 32'sd0.045279583778635384, 32'sd-0.09910703699921282, 32'sd0.042918717869391255, 32'sd0.010429280592351863, 32'sd0.03161865072284231, 32'sd-0.11814124344907444, 32'sd-0.0831067288184278, 32'sd-0.05927122332865006, 32'sd-0.1666483679709285, 32'sd-0.01143977116323252, 32'sd-0.008499280753851342, 32'sd-0.07485174726614897, 32'sd-0.09047366396926844, 32'sd-0.1387962907636765, 32'sd-0.19062942839248456, 32'sd-0.15114009255654223, 32'sd-0.19773377326084945, 32'sd-0.0491775146986461, 32'sd0.0907139260709738, 32'sd-0.04367107021032991, 32'sd0.022933767334653243, 32'sd0.038920902490646093, 32'sd0.005832820980881177, 32'sd-0.11791850211036994, 32'sd0.04717038576200876, 32'sd0.052415235697641706, 32'sd0.05736424352123656, 32'sd0.003067138974964327, 32'sd-0.08737978123248678, 32'sd-0.1663257802954066, 32'sd-0.1609535817530516, 32'sd-0.15914011903855202, 32'sd-0.17491713873953266, 32'sd-0.1886481140832679, 32'sd-0.1379491735035153, 32'sd-0.13412502872284993, 32'sd-0.10610009127585543, 32'sd-0.0316229400955621, 32'sd0.011714585330899231, 32'sd0.00010369901193203531, 32'sd-0.05733199240766414, 32'sd-0.08346676881934377, 32'sd-0.06571112615712256, 32'sd-0.1550631208177122, 32'sd-0.11282372053529852, 32'sd-0.1030189580571113, 32'sd0.024275626575775533, 32'sd0.10668343277408168, 32'sd0.07569792570655355, 32'sd0.04097994108105526, 32'sd-0.06587801299204463, 32'sd0.09275846790943439, 32'sd0.07983131935369832, 32'sd7.17772498421811e-118, 32'sd0.07397179014268293, 32'sd0.0485157749770698, 32'sd-0.011980922709679702, 32'sd-0.0653699917200031, 32'sd-0.020728437264660938, 32'sd-0.02690046448003902, 32'sd-0.06183182944749438, 32'sd-0.13358908918121423, 32'sd-0.11320778130437911, 32'sd-0.1785103641759816, 32'sd-0.2546476785702249, 32'sd-0.19152418260099474, 32'sd-0.11301429721215521, 32'sd-0.029586094892830754, 32'sd-0.0399760391692129, 32'sd-0.06678844637347697, 32'sd-0.05941039464690537, 32'sd-0.14538232396255965, 32'sd-0.13015697358535241, 32'sd0.04247039993899171, 32'sd0.09785161186828022, 32'sd0.10612201331037371, 32'sd0.05249694261892395, 32'sd0.013704345291455982, 32'sd-0.04316751019099925, 32'sd0.019597873938574435, 32'sd-0.018066334758632802, 32'sd0.027467584766294222, 32'sd0.022950822655291594, 32'sd0.12479650749777273, 32'sd0.08684827720017535, 32'sd-0.018355579885194324, 32'sd-0.09734187177410285, 32'sd-0.07513341678884088, 32'sd-0.11704221594281264, 32'sd-0.11849268407673466, 32'sd-0.19741722111505075, 32'sd-0.12577587969319243, 32'sd-0.14998017556288298, 32'sd-0.17583947821740578, 32'sd-0.11250963885880458, 32'sd-0.07691178885219167, 32'sd-0.19713984058513578, 32'sd-0.01252110123957168, 32'sd-0.052402925823238404, 32'sd-0.09366499700875373, 32'sd-0.009180142641829536, 32'sd0.03537270879295725, 32'sd0.13190166661134986, 32'sd0.10190363857759165, 32'sd0.10717682834235352, 32'sd0.07727356417685334, 32'sd0.02438432634281388, 32'sd-0.1329113056583785, 32'sd0.08165122181903302, 32'sd0.06915557000452893, 32'sd-0.06569186391464071, 32'sd0.10641942923454982, 32'sd0.11482181106229916, 32'sd0.01805641289573148, 32'sd-0.0005556548228769162, 32'sd0.07179875448879323, 32'sd0.00445979432555705, 32'sd-0.10905333167815387, 32'sd-0.16923988808049437, 32'sd-0.2523797277796675, 32'sd-0.12405681970533594, 32'sd-0.14004030699400763, 32'sd-0.03107062499564138, 32'sd-0.14254443049733082, 32'sd-0.12925363434311604, 32'sd-0.000537128615172884, 32'sd-0.05064974437442929, 32'sd0.05184309192701064, 32'sd0.04260006248265331, 32'sd0.049366054899738464, 32'sd0.0019528550263468844, 32'sd0.11160315293104588, 32'sd-0.01947063776406683, 32'sd0.005827810746405663, 32'sd0.05552028954061337, 32'sd-0.04558106662749198, 32'sd0.026565308660262382, 32'sd-1.7168379805425924e-122, 32'sd-0.04542050099369917, 32'sd-0.022417133745793082, 32'sd0.06890039112682206, 32'sd0.08237296947074949, 32'sd0.09064215768054103, 32'sd0.08932857749217253, 32'sd0.004808242984217999, 32'sd0.050017176198399384, 32'sd-0.021874609607996382, 32'sd0.002750047704207531, 32'sd0.05835464950797051, 32'sd0.02638737645917047, 32'sd0.07252852068719212, 32'sd0.0032359559059373893, 32'sd-0.030524209235437597, 32'sd0.1102235662658374, 32'sd0.033864138129071256, 32'sd-0.012236282151902672, 32'sd0.15969990467476278, 32'sd-0.010052785690480508, 32'sd-0.00875725053941626, 32'sd0.026897076492266973, 32'sd-0.02098664528368967, 32'sd0.04991919890850391, 32'sd-0.03684544949456933, 32'sd-0.026633466107338553, 32'sd0.06110437080719595, 32'sd0.09269680939738105, 32'sd-0.006640178854779079, 32'sd0.015445610346967736, 32'sd0.03495593526188403, 32'sd0.15994360616357323, 32'sd0.14060061125183734, 32'sd0.04638107700907043, 32'sd0.1276990709879546, 32'sd0.15563442029371227, 32'sd0.14698501316054566, 32'sd0.061070618572322585, 32'sd0.10763225933747822, 32'sd0.13791044809115335, 32'sd0.12963823368268435, 32'sd0.23214088654256304, 32'sd0.09617067010942319, 32'sd-0.09725647297219396, 32'sd-0.016311494659372604, 32'sd0.07838059699423498, 32'sd-0.05062899859234692, 32'sd-0.013645192489000644, 32'sd0.005594074666853, 32'sd0.019925925322084467, 32'sd-0.035251307775194175, 32'sd0.0017913812729530483, 32'sd0.10804273112275242, 32'sd-0.09250208695845526, 32'sd0.05541053660182808, 32'sd0.05297640976846692, 32'sd0.05641780592960075, 32'sd0.06950586071187695, 32'sd0.09107978206653954, 32'sd0.06858007208201941, 32'sd0.006638562467040546, 32'sd0.013291224886886317, 32'sd-0.019529864516707893, 32'sd0.09325234215507652, 32'sd0.018097087652866117, 32'sd0.07292458594757002, 32'sd0.14855597907189483, 32'sd0.04955587911605834, 32'sd0.053416489474794285, 32'sd0.11689656936409137, 32'sd0.13248651121284108, 32'sd0.02305313399693789, 32'sd-0.04685227358881212, 32'sd-0.0008920322636979769, 32'sd0.007809994919786803, 32'sd0.10580360369733617, 32'sd-0.03134187952972173, 32'sd-0.013665251790822721, 32'sd0.07952408581435891, 32'sd-0.015766635404402565, 32'sd0.024641614994478176, 32'sd0.06048273550040584, 32'sd0.049781789934567625, 32'sd4.319320257084091e-118, 32'sd0.11774477740965691, 32'sd-0.0013169473194573466, 32'sd-0.03431228641802487, 32'sd0.03712365764901817, 32'sd0.1883892722087122, 32'sd0.05165707937465284, 32'sd0.07302978306799966, 32'sd-0.028473577968460166, 32'sd-0.06347988107624647, 32'sd0.06751465797725036, 32'sd-0.00461077514395401, 32'sd-0.06360394593152753, 32'sd0.040470367747656215, 32'sd0.09234290570951778, 32'sd0.0767431340581594, 32'sd0.09149143069712028, 32'sd0.025754526539363026, 32'sd0.1281518329348698, 32'sd0.029564405751533424, 32'sd0.069516568995491, 32'sd0.03711844646776197, 32'sd0.08181674361030944, 32'sd-0.012206560630402982, 32'sd0.034738327937270524, 32'sd0.09286100005052282, 32'sd-0.010843978359635666, 32'sd-1.1361860734326667e-116, 32'sd3.010064259990856e-128, 32'sd-8.492790196284544e-121, 32'sd0.04762025033123627, 32'sd0.02205205522127231, 32'sd-0.05902205754350639, 32'sd-0.05714059018419526, 32'sd0.05080501609994329, 32'sd0.11110984065430761, 32'sd0.006828745871845324, 32'sd0.010205150756777108, 32'sd-0.009594561213069425, 32'sd0.02826951324220858, 32'sd0.005637687349134428, 32'sd-0.042860389130130544, 32'sd0.10781899827824944, 32'sd-0.00047528030808681676, 32'sd-0.045724217883049256, 32'sd0.10298327095323083, 32'sd0.17014671176551593, 32'sd0.06656450127730985, 32'sd-0.06956408024735579, 32'sd-0.018847096099890024, 32'sd0.06044292638899234, 32'sd0.05151937215714339, 32'sd-0.02757604352371203, 32'sd-0.026230231394134013, 32'sd0.025679923669179382, 32'sd-1.276162038627306e-127, 32'sd-1.0229936049261528e-125, 32'sd1.7809845486889174e-117, 32'sd-0.0007499205169867555, 32'sd-0.02121610610908181, 32'sd0.013406227893428593, 32'sd-0.04753690594449954, 32'sd0.04348302011148966, 32'sd0.05663188692430748, 32'sd-0.01953842355395545, 32'sd0.026670191929967, 32'sd-0.02898939675688192, 32'sd0.11675332939232841, 32'sd0.03747754057846839, 32'sd0.21436423667049878, 32'sd0.018043592871562528, 32'sd-0.06596854335321804, 32'sd0.0969236009593321, 32'sd0.057948035027137676, 32'sd0.06065771503435075, 32'sd0.07410069653607515, 32'sd0.011947208614498479, 32'sd0.02442360771483028, 32'sd0.08286307694384343, 32'sd0.044541206076872154, 32'sd0.005455180917709656, 32'sd0.07053642426676042, 32'sd0.08366103854097724, 32'sd-3.547791431644072e-116, 32'sd-1.0465802856707858e-120, 32'sd2.1883568044594293e-124, 32'sd-5.126199347604704e-118, 32'sd0.11214337842974155, 32'sd0.04864964033754464, 32'sd-0.03843638463269173, 32'sd0.031419427256157824, 32'sd-0.02525167355391942, 32'sd0.020927982390064923, 32'sd0.009527039388621745, 32'sd0.01841139327417232, 32'sd0.03343079180373938, 32'sd0.0750416151525955, 32'sd0.09347433449957629, 32'sd0.0200721531056297, 32'sd0.08794855214500627, 32'sd0.04396687149563933, 32'sd-0.0008277240947530079, 32'sd-0.06784404399910465, 32'sd-0.10382689849414238, 32'sd0.012337108442962116, 32'sd-0.04187287960980067, 32'sd0.011879058071498512, 32'sd-0.05842202836938565, 32'sd0.08582267958312627, 32'sd0.07820292466909387, 32'sd-3.116682653232099e-125, 32'sd4.861647454797491e-127, 32'sd5.135653923126116e-121, 32'sd1.7940626055241652e-117, 32'sd-1.7933783537702205e-123, 32'sd-1.999559007362085e-127, 32'sd0.11920896369673387, 32'sd0.013069817393297012, 32'sd0.021840420629941383, 32'sd0.0893114837330482, 32'sd0.03115883170155575, 32'sd0.0439591788120705, 32'sd0.0972365439253439, 32'sd0.04684001142738819, 32'sd-0.0015089639324834614, 32'sd0.07921443025455852, 32'sd0.07091827037163029, 32'sd0.10921306247755277, 32'sd0.10734628350007502, 32'sd0.0650889368534927, 32'sd0.04830452793746682, 32'sd-0.04352309972535233, 32'sd0.06821370134647778, 32'sd0.008256738696547838, 32'sd-0.10561452038448012, 32'sd0.13262490578128244, 32'sd1.766348529945261e-126, 32'sd-6.007249221583761e-128, 32'sd-1.9328091417956054e-119, 32'sd1.0484762056942288e-119},
        '{32'sd-2.718604221830945e-125, 32'sd2.4187195571114205e-123, 32'sd-1.4362845798298787e-118, 32'sd4.869867385937299e-123, 32'sd3.2535864831962185e-120, 32'sd7.110943370636708e-120, 32'sd-1.6911849283416815e-117, 32'sd1.14873136813452e-117, 32'sd-4.882050268720733e-122, 32'sd-1.0487094034767105e-122, 32'sd-5.456377446607381e-115, 32'sd-7.41906303392845e-120, 32'sd-0.07931034954894427, 32'sd0.036647484107643805, 32'sd0.09835904087251061, 32'sd0.022861957456745297, 32'sd8.335874696561723e-124, 32'sd1.3006154217179211e-118, 32'sd3.3835415354659156e-120, 32'sd4.173342840409709e-118, 32'sd-3.8113155313256595e-120, 32'sd-6.244407623792348e-116, 32'sd-4.483393872412093e-123, 32'sd-3.675455530000432e-116, 32'sd-1.7951622276872987e-127, 32'sd2.7485657652650015e-122, 32'sd-1.2301769634281127e-124, 32'sd1.2447926730833575e-115, 32'sd4.35748229447777e-124, 32'sd2.5887301405716644e-124, 32'sd6.534890380999019e-126, 32'sd-6.586235139043038e-121, 32'sd-0.03221261988631944, 32'sd0.0003068462546269217, 32'sd-0.038222067169307976, 32'sd0.06288221981008725, 32'sd-0.10038578973171677, 32'sd0.05214361377727304, 32'sd0.08496488664379777, 32'sd-0.01714419341522216, 32'sd-0.0010715441089512341, 32'sd0.15736601298358602, 32'sd0.10125630987450052, 32'sd0.020492386734338577, 32'sd0.07979576385559037, 32'sd0.025548971210587492, 32'sd-0.021808206326942345, 32'sd-0.0459819076502885, 32'sd-0.04668538098999562, 32'sd-0.0442415614568923, 32'sd0.06612047808156633, 32'sd-0.019590454902244966, 32'sd-6.741605478928014e-124, 32'sd1.3256766751918406e-118, 32'sd-9.061274530840335e-123, 32'sd-1.1298780206376604e-119, 32'sd1.734972627071659e-125, 32'sd-3.788982294816552e-129, 32'sd0.031035094587454504, 32'sd-0.016006305389425983, 32'sd-0.03074959585149789, 32'sd0.07724097136136367, 32'sd-0.060570024043888705, 32'sd-0.0014850529536799013, 32'sd-0.013166749891738052, 32'sd0.08579534236715451, 32'sd0.046923843050702865, 32'sd0.07889127766718186, 32'sd0.002658663196906098, 32'sd-0.030795076616016433, 32'sd0.027322274937652918, 32'sd-0.02124476831302824, 32'sd-0.11071947970570122, 32'sd0.11363861982004406, 32'sd-0.020532687533138888, 32'sd-0.12009391956064197, 32'sd0.02475916809547202, 32'sd0.010294620166140623, 32'sd0.047869902795354, 32'sd0.022643808795441724, 32'sd0.012497823198028673, 32'sd-0.04444838140270689, 32'sd-1.2274422184413717e-125, 32'sd-6.739369504870084e-115, 32'sd-4.947764115611781e-118, 32'sd-7.046990686960161e-115, 32'sd-0.059587818048568726, 32'sd-0.025583313842390886, 32'sd0.052004363499974705, 32'sd0.0075183254447727405, 32'sd0.11797069118923609, 32'sd0.10375478621811848, 32'sd0.05665571886087625, 32'sd-0.04359311991439559, 32'sd0.09908456782851732, 32'sd0.038894538717080755, 32'sd0.017549777965843394, 32'sd0.04396858103001494, 32'sd-0.008073002675707427, 32'sd-0.004615573068987523, 32'sd-0.07577727551824819, 32'sd-0.04063157801185993, 32'sd-0.02331934904027427, 32'sd-0.021379802253850517, 32'sd0.023815388034312216, 32'sd-0.03441923864026444, 32'sd0.09465329023371766, 32'sd0.04921754309557724, 32'sd-0.0438491098066783, 32'sd0.03410852021461607, 32'sd0.0680683425866357, 32'sd1.0972493414078404e-122, 32'sd1.0442186944748869e-120, 32'sd0.07116440164862188, 32'sd0.06825294653206102, 32'sd0.012073252245345598, 32'sd0.015279293377904249, 32'sd0.05808467560273664, 32'sd-0.0773151738411018, 32'sd0.010836740926950441, 32'sd0.048854072718235754, 32'sd-0.06067043267453717, 32'sd0.18174235821272958, 32'sd0.07742523011705567, 32'sd0.06244708768784634, 32'sd-0.037620637969029806, 32'sd0.0929616892473016, 32'sd-0.09859257232532598, 32'sd0.008068263895737312, 32'sd0.1043895903124263, 32'sd0.039589033352403914, 32'sd0.07178532701374063, 32'sd0.002592112070234016, 32'sd0.03781975160348151, 32'sd0.018246255899473148, 32'sd0.009533251314918901, 32'sd0.10483880165453283, 32'sd0.019794936048557824, 32'sd0.05300904995644094, 32'sd-0.0031095549226554525, 32'sd1.7793414073227202e-121, 32'sd-0.006894699875414417, 32'sd0.08639888103406937, 32'sd0.10396580393166298, 32'sd0.024256860106718486, 32'sd0.029537114406235215, 32'sd-0.07449158279014975, 32'sd-0.01917548558061466, 32'sd0.0481248932835703, 32'sd-0.061045046599041204, 32'sd-0.011953696591384259, 32'sd0.04410698758718948, 32'sd0.10838660041776284, 32'sd0.21184062569020382, 32'sd0.15178661650464267, 32'sd-0.0019020961036220513, 32'sd0.07110393199145905, 32'sd-0.03686867749932599, 32'sd0.005048065965281098, 32'sd0.0017005541791973472, 32'sd0.022628593779329024, 32'sd-0.06406270031812393, 32'sd-0.08059170665557103, 32'sd-0.12293716757138129, 32'sd0.04496745184699596, 32'sd0.09680454021955129, 32'sd0.08322634810051767, 32'sd0.014835295061204854, 32'sd-1.2585745583373951e-125, 32'sd0.007164560901369814, 32'sd-0.0002677016377029517, 32'sd-0.08558966812598635, 32'sd-0.10424127404068531, 32'sd-0.059162462597185564, 32'sd0.024356063675483014, 32'sd0.06357701590428562, 32'sd0.09182007735564468, 32'sd0.03792894093025078, 32'sd0.03450257873549175, 32'sd0.06413859329362957, 32'sd0.1789574918207237, 32'sd0.23768865327226793, 32'sd0.14722822383349682, 32'sd0.11614084495244557, 32'sd-0.03861979218508677, 32'sd-0.07256219315029665, 32'sd-0.09961768641372855, 32'sd-0.08630934613702075, 32'sd-0.04573736690483551, 32'sd-0.024779299956063663, 32'sd-0.06854231122706446, 32'sd0.04053095921312592, 32'sd-0.12367952128963959, 32'sd-0.054536752354905946, 32'sd-0.03976672597190927, 32'sd-0.016764818258268793, 32'sd0.02444122878857302, 32'sd-0.037041715083704935, 32'sd0.05960766235810122, 32'sd-0.05580871837466767, 32'sd-0.0006651923900266346, 32'sd-0.0821044298518971, 32'sd-0.02795914389486081, 32'sd0.007927453329355445, 32'sd0.1218453249682225, 32'sd0.024132172231105583, 32'sd0.05296500340279072, 32'sd0.1369225203567366, 32'sd0.07913136408901983, 32'sd0.0887658918854922, 32'sd0.04271561696492061, 32'sd0.04586857532794235, 32'sd-0.074774441773611, 32'sd0.027003035901351766, 32'sd-0.07397290370034543, 32'sd-0.043256995311544574, 32'sd-0.029633117354397057, 32'sd0.01364453659033309, 32'sd0.001388954470533481, 32'sd0.04260299298993347, 32'sd-0.010964955997475542, 32'sd-0.042286132003860055, 32'sd-0.08872922226608762, 32'sd-0.026450218356786657, 32'sd-0.0009046982837877436, 32'sd-0.01631293497524179, 32'sd0.07663366967891866, 32'sd0.118970942898262, 32'sd0.10528427492231385, 32'sd0.08989993233177081, 32'sd0.002808626536062574, 32'sd0.02604069288792048, 32'sd0.10272633138947439, 32'sd0.02930589315134726, 32'sd0.1819133122001017, 32'sd0.12833281556429457, 32'sd0.12283324251088268, 32'sd0.06442190063964968, 32'sd-0.04791994254179659, 32'sd-0.036391864736045186, 32'sd0.04614010707097942, 32'sd1.570633162882056e-05, 32'sd-0.038058162121647914, 32'sd-0.09056438353103854, 32'sd-0.015781483858239572, 32'sd-0.012128722691586536, 32'sd-0.04891963158979464, 32'sd-0.04003496932525979, 32'sd-0.14712943383612082, 32'sd0.01834500651291771, 32'sd-0.022814576637888623, 32'sd0.02739508830575245, 32'sd-0.04568117191523577, 32'sd0.022769787847042155, 32'sd0.013360380016643494, 32'sd0.0506450902087692, 32'sd0.00887995767817712, 32'sd0.04624787410762654, 32'sd-6.945870876924266e-05, 32'sd0.05124666704215665, 32'sd-0.034445105155923125, 32'sd0.08418943925603001, 32'sd0.035593612532867434, 32'sd-0.11584101065872669, 32'sd-0.13342305582810365, 32'sd-0.046369729398553605, 32'sd0.06024413457112946, 32'sd-0.035799344360701556, 32'sd0.021005006085280716, 32'sd0.045660171447221266, 32'sd0.010108065651955387, 32'sd0.023295345504777316, 32'sd0.114629052539821, 32'sd-0.023578373935703247, 32'sd0.008335389130241132, 32'sd-0.02720307225741631, 32'sd-0.16105203031204, 32'sd-0.0891935687077537, 32'sd0.048353650378635205, 32'sd0.015244536660973614, 32'sd0.030782419898714858, 32'sd-0.0597328294174144, 32'sd-0.035491064461810794, 32'sd0.17276057012448243, 32'sd0.05169377036290796, 32'sd0.00808480985576575, 32'sd0.09410352394413495, 32'sd-0.10319430423465599, 32'sd-0.01619131438050254, 32'sd-0.01893484553866811, 32'sd-0.09692095895604734, 32'sd-0.1779703737169182, 32'sd-0.21738064444366625, 32'sd-0.17286077503095462, 32'sd0.010142216585396846, 32'sd0.03768492354250889, 32'sd0.15833952839434529, 32'sd0.1172449408523592, 32'sd0.07085108820255251, 32'sd-0.010605211547801106, 32'sd0.0783187508156365, 32'sd-0.06026385031140259, 32'sd0.02777093967985508, 32'sd-0.03854287087525173, 32'sd-0.11830888129384054, 32'sd-0.007851656458034305, 32'sd0.029881805492485133, 32'sd-0.07143993713959892, 32'sd-0.0008840177102119527, 32'sd0.012061214163840879, 32'sd0.06958554888233996, 32'sd0.10403397217288952, 32'sd0.001343879381060679, 32'sd-0.007824563195248192, 32'sd-0.022488470091074086, 32'sd-0.08771729425091673, 32'sd-0.07751132199873777, 32'sd-0.018210389679849205, 32'sd-0.032511471858129894, 32'sd0.05996138586401785, 32'sd-0.01284344586363655, 32'sd0.03509637498790176, 32'sd0.04804062705564021, 32'sd-0.04848298098041072, 32'sd0.10235964359197375, 32'sd0.11269364568300377, 32'sd0.051035283265761164, 32'sd0.0038443188998997057, 32'sd0.007810794981621179, 32'sd0.023274821065978196, 32'sd0.05599808860659438, 32'sd-0.13955732886830052, 32'sd-0.05146858195760412, 32'sd0.010614568935860881, 32'sd0.06826344624343654, 32'sd0.037987713008292436, 32'sd0.021711610481182194, 32'sd-0.045910333136828574, 32'sd-0.05746876107643776, 32'sd-0.013537989095287181, 32'sd0.07435160265585479, 32'sd-0.004418916751926128, 32'sd0.014882721573375238, 32'sd-0.07419327185996658, 32'sd-0.07875076415843349, 32'sd-0.02817632037194859, 32'sd-0.20599561675408226, 32'sd0.02894005513072947, 32'sd0.034818307552935454, 32'sd-0.04785461470696356, 32'sd0.009521856799781458, 32'sd0.09057290412882034, 32'sd-0.04024778276934933, 32'sd0.04493620659698554, 32'sd-0.08723747438732823, 32'sd0.12170698812463536, 32'sd-0.046472434118922476, 32'sd-0.01805203385718678, 32'sd-0.13182187729877298, 32'sd-0.1435519497011079, 32'sd-0.04710352936298163, 32'sd0.06546956782263691, 32'sd-0.05211320006825918, 32'sd-0.08198822224985147, 32'sd0.02158175312217789, 32'sd0.040762733129183396, 32'sd0.13157300012897494, 32'sd-0.11043823870155518, 32'sd-0.10141071794300559, 32'sd0.04576098459144395, 32'sd0.0028782062713756636, 32'sd-0.05768877131208149, 32'sd-0.07675703262852185, 32'sd-0.03405924165813329, 32'sd-0.06190601643315125, 32'sd0.016198899652483514, 32'sd-0.07209870203370022, 32'sd0.028489520047892354, 32'sd0.1236534487652374, 32'sd0.09550744539884616, 32'sd-0.05259676454027371, 32'sd-0.10917636579925058, 32'sd-0.07727890608545715, 32'sd-0.09941253201636542, 32'sd-0.04718330613456252, 32'sd-0.09807704053045178, 32'sd-0.11966344563776249, 32'sd-0.05510817968229643, 32'sd-0.06848889197673716, 32'sd0.054977832105748185, 32'sd-0.14643505481827182, 32'sd-0.006594909324862217, 32'sd0.0024304714087164283, 32'sd0.025358864519504035, 32'sd0.06973695284416202, 32'sd0.04204372494850254, 32'sd-0.1268636714908798, 32'sd0.0029342628673247268, 32'sd-0.1011788057096332, 32'sd-0.04632381588342136, 32'sd-0.13005431849042837, 32'sd-0.14108313538839198, 32'sd-0.11580246982146607, 32'sd0.05039361973477245, 32'sd0.011032469432190379, 32'sd0.07889202235028345, 32'sd0.2431126313308119, 32'sd0.141206957167927, 32'sd-0.050920385878990976, 32'sd-0.13109034261234123, 32'sd-0.13146260475739466, 32'sd-0.12075389206841913, 32'sd-0.07579504959071982, 32'sd-0.022925935790864327, 32'sd-0.18036940582020436, 32'sd-0.06144751141887327, 32'sd-0.1487083835121228, 32'sd0.0078033403569961034, 32'sd-0.012756552058222181, 32'sd0.04332001480247015, 32'sd-0.027290762242681756, 32'sd0.08194209940379132, 32'sd0.01244394601512171, 32'sd0.010712814420012104, 32'sd-0.1284217160749318, 32'sd0.043691726493407294, 32'sd0.028210802067309613, 32'sd-0.03742469523246236, 32'sd-0.04493226229453683, 32'sd-0.1703029442653491, 32'sd-0.17489587602248238, 32'sd0.11493732775636127, 32'sd0.170601244953965, 32'sd0.21006692400538815, 32'sd0.27504487969351443, 32'sd0.1479606209072313, 32'sd-0.014422623963434418, 32'sd-0.007524958966411285, 32'sd-0.03837744864275999, 32'sd-0.15314082345546237, 32'sd-0.10785424180553001, 32'sd-0.04179670522934942, 32'sd-0.1661964510537399, 32'sd-0.03678465943725774, 32'sd-0.031038649657017754, 32'sd0.02146422489792125, 32'sd-0.09870931750739839, 32'sd-0.039406226767183736, 32'sd-0.024113571791037174, 32'sd-0.015555693447812508, 32'sd0.06171999591686186, 32'sd0.027550472379337682, 32'sd-0.07471374036100244, 32'sd-0.06095031679859305, 32'sd0.011141839822231502, 32'sd-0.012126492841472896, 32'sd-0.029092553266043802, 32'sd0.024136783172628903, 32'sd0.009047533548545181, 32'sd0.057682609389659176, 32'sd0.024458183043600874, 32'sd0.1187303524078937, 32'sd0.18369973633629302, 32'sd0.010959311845687911, 32'sd0.05612571738603208, 32'sd0.0872079893266771, 32'sd0.01824858753456458, 32'sd-0.010775418650001827, 32'sd-0.004982559235476488, 32'sd-0.005215828001310717, 32'sd-0.10217311302900633, 32'sd0.05051187221414194, 32'sd0.017842790239870367, 32'sd0.04864617788739087, 32'sd0.03028886505705789, 32'sd0.03875035871442977, 32'sd3.17663165174133e-114, 32'sd-0.03336570040674855, 32'sd0.005207329580170174, 32'sd-0.011731930725896336, 32'sd-0.05600422895211382, 32'sd-0.13380622972468148, 32'sd0.013507451462962148, 32'sd-0.16432669883155834, 32'sd-0.1241559237139953, 32'sd0.011492001041527852, 32'sd-0.03839796735357578, 32'sd0.00962699894297147, 32'sd-0.004824023103125131, 32'sd0.12722365317795087, 32'sd0.0785291707945219, 32'sd0.050551431326651214, 32'sd-0.005878228646969383, 32'sd0.061247041829530294, 32'sd-0.026851356524245213, 32'sd-0.002749895257506137, 32'sd0.07918254836441632, 32'sd0.040921555686703, 32'sd0.022935392451046595, 32'sd0.02213240979609162, 32'sd0.12074316353074017, 32'sd0.0951037703825297, 32'sd-0.028670827241780366, 32'sd0.049937582257966094, 32'sd-0.009325904843660693, 32'sd-0.03340670727767906, 32'sd0.061983805030996056, 32'sd0.07694969942667379, 32'sd-0.03317006688228144, 32'sd-0.10332023590025571, 32'sd-0.06729674219562404, 32'sd-0.16390005727276177, 32'sd0.003618762079375903, 32'sd0.11263338675102502, 32'sd0.027585705898246826, 32'sd-0.0024727987905653393, 32'sd0.0734225647880093, 32'sd-0.10253313272699066, 32'sd-0.05428798777377844, 32'sd0.04463963974441356, 32'sd0.09702165611554693, 32'sd0.06536305891235623, 32'sd0.10285792790902705, 32'sd0.11260543531490656, 32'sd0.11844534780144282, 32'sd0.08604825130296943, 32'sd0.0778317595275922, 32'sd-0.017644654609703374, 32'sd-0.031401507575296445, 32'sd0.12310349502406584, 32'sd0.10920287022457191, 32'sd-0.006422046588023331, 32'sd0.0001433978263294199, 32'sd0.013462703047853191, 32'sd0.030743762577896717, 32'sd0.10775318081809025, 32'sd-0.1551841682520068, 32'sd-0.1755940382385227, 32'sd-0.20233104481156353, 32'sd0.03767077993180709, 32'sd0.07391528580064038, 32'sd0.09633640515854715, 32'sd0.11486676752289524, 32'sd-0.07402003998473322, 32'sd-0.1172238526809687, 32'sd-0.09468008717888567, 32'sd-0.07362335793768936, 32'sd-0.007445420097744071, 32'sd-0.0314990900531556, 32'sd-0.037067238170079876, 32'sd0.07652132607152339, 32'sd0.010618304278204923, 32'sd0.10672094271640374, 32'sd-0.030038860035354182, 32'sd0.04640727190790041, 32'sd-0.05840186295162968, 32'sd0.0324699966602454, 32'sd-0.03159515764223721, 32'sd0.06910978732701585, 32'sd-0.07670650454643788, 32'sd3.931860365463771e-118, 32'sd0.006407736636995936, 32'sd-0.04110095499279863, 32'sd-0.05235068707016105, 32'sd-0.08249130916748863, 32'sd-0.12538635401910675, 32'sd-0.13422220891647715, 32'sd0.0658777767923162, 32'sd0.13903870291329595, 32'sd0.14992993047423347, 32'sd0.14947049120153658, 32'sd0.023187710385916178, 32'sd-0.08899531236372343, 32'sd-0.0588149593231278, 32'sd-0.08419442538591801, 32'sd0.06548282691696994, 32'sd-0.06534089088108891, 32'sd-0.13909379500326866, 32'sd-0.06560568740486167, 32'sd0.05521608423063354, 32'sd0.11280549715206371, 32'sd-0.03512070495897816, 32'sd-0.052963581150197024, 32'sd0.09257592246462329, 32'sd0.07501685253421014, 32'sd-0.07414441480297236, 32'sd-0.1095962165864129, 32'sd-0.011592987112777375, 32'sd-0.01713320750457478, 32'sd0.028634854858666653, 32'sd0.05828872128312947, 32'sd0.09997281408835038, 32'sd0.002088980446233547, 32'sd-0.10462265343224132, 32'sd-0.019289303380645002, 32'sd0.025901180744837313, 32'sd0.12679953018514523, 32'sd-0.031702179197201426, 32'sd0.006155255419361204, 32'sd-0.05349070579385793, 32'sd-0.046607218338363614, 32'sd-0.010109777119953842, 32'sd-0.0036029071966856593, 32'sd-0.05424991716682184, 32'sd-0.0816209210472108, 32'sd-0.10945904515361102, 32'sd0.02856660631244121, 32'sd-0.0009799387943071106, 32'sd0.037711734334853725, 32'sd0.05320888420320879, 32'sd-0.005230630156918612, 32'sd0.08978943976584887, 32'sd-0.0003694272379359726, 32'sd-0.11696455789144973, 32'sd-0.12085865901791804, 32'sd0.0071437223580876645, 32'sd-0.0003011720697456821, 32'sd0.017438805227375655, 32'sd-0.01970670588803624, 32'sd0.12785315302999598, 32'sd-0.06317882022342347, 32'sd0.04979642126383424, 32'sd0.043201900771005504, 32'sd0.12544310015163315, 32'sd0.07748944630165126, 32'sd0.09042268765496712, 32'sd-0.06746629176239721, 32'sd-0.04875714218371183, 32'sd0.09911724660448681, 32'sd-0.005302491655452157, 32'sd0.014607714437035105, 32'sd0.1283476546559428, 32'sd0.04400245881702716, 32'sd-0.02497324230368132, 32'sd0.06219358544575469, 32'sd0.06828661108096047, 32'sd-0.04361297086079562, 32'sd0.01943220238376433, 32'sd0.027396974819798806, 32'sd0.10865829495645143, 32'sd0.05580173264177992, 32'sd-0.0039729948092940065, 32'sd-0.10794766663720128, 32'sd-0.03512790067143753, 32'sd-7.174603080370269e-127, 32'sd0.0360649077397703, 32'sd0.07771397809675101, 32'sd-0.04063562312640944, 32'sd0.02015764533640367, 32'sd0.04380023619418721, 32'sd0.04995223319840911, 32'sd0.12301846877489361, 32'sd0.0693264985273952, 32'sd0.13459858073268788, 32'sd-0.03411851743864284, 32'sd0.04732811136314951, 32'sd0.07314092573394962, 32'sd-0.049614714194358145, 32'sd0.037502027622752954, 32'sd0.02602441867158542, 32'sd0.01911747512439615, 32'sd0.114683515203764, 32'sd0.0853650900169824, 32'sd0.053962563707466216, 32'sd0.09911131214395325, 32'sd-0.07937993244162968, 32'sd0.07781959793680243, 32'sd0.07858258135345551, 32'sd-0.03872802012341033, 32'sd0.03305385216133065, 32'sd-0.08237251495792945, 32'sd1.167082799808512e-118, 32'sd-1.1014422979192064e-119, 32'sd-6.992328714881379e-117, 32'sd0.06812196202769273, 32'sd0.05752214754398148, 32'sd-0.008951827380244472, 32'sd-0.021493542439291007, 32'sd0.09531921282399268, 32'sd0.036280375837330694, 32'sd0.06583104685076292, 32'sd-0.004015502214549074, 32'sd-0.0704362407111168, 32'sd0.06150386698619943, 32'sd0.07447948775295503, 32'sd-0.04358343499748185, 32'sd-0.03120864212624019, 32'sd-0.0029261307428346105, 32'sd-0.0104050490167522, 32'sd-0.01848870066737355, 32'sd0.006658911340828964, 32'sd-0.08615733741585982, 32'sd-0.027198054760478804, 32'sd-0.04619073732449205, 32'sd0.07961531008102585, 32'sd-0.024302622457670828, 32'sd0.01004969152207395, 32'sd0.07190044857787248, 32'sd-0.04480619153727074, 32'sd1.8695840119680298e-119, 32'sd-9.364951468596204e-121, 32'sd-9.497400662464021e-128, 32'sd-0.01159538188567364, 32'sd0.02201412481099435, 32'sd0.06852798425138279, 32'sd0.023605177809732498, 32'sd0.031832583959847865, 32'sd0.07441126152820376, 32'sd-0.058902690143790015, 32'sd-0.10331461246754321, 32'sd-0.027949182165939876, 32'sd-0.07484494573121074, 32'sd-0.036960369590257704, 32'sd0.02914706446151055, 32'sd0.05637486469741467, 32'sd0.1341437356785315, 32'sd0.1183145373915038, 32'sd0.13618189221967072, 32'sd0.043395502705399915, 32'sd-0.08733496029819258, 32'sd0.00019662150844311737, 32'sd-0.031832929559938036, 32'sd-0.03329419266867559, 32'sd-0.03901948146951286, 32'sd-0.06479145266752082, 32'sd0.05967629485371137, 32'sd0.059605133998309696, 32'sd-3.0081880198857447e-124, 32'sd6.877786381514899e-126, 32'sd-5.056934604642698e-125, 32'sd2.344503479942566e-122, 32'sd-0.027670961108028476, 32'sd0.0357994437242473, 32'sd-0.011826235452608582, 32'sd-0.0032617404440058767, 32'sd-0.04598545042954351, 32'sd0.10298510763642847, 32'sd0.0712659979909304, 32'sd-0.045942230276168984, 32'sd-0.009197446975698255, 32'sd0.08842144877489821, 32'sd-0.013801703450346514, 32'sd-0.030826838767441484, 32'sd-0.01423063325365445, 32'sd0.016016949110408584, 32'sd0.0164649274523886, 32'sd0.07918095339174457, 32'sd0.03376952674254552, 32'sd-0.03171217588485288, 32'sd-0.01693089737445451, 32'sd0.06303090834593558, 32'sd-0.06290508908497712, 32'sd0.014357679531321445, 32'sd-0.03192129903760846, 32'sd1.1209852573512605e-122, 32'sd3.8061551381155014e-120, 32'sd1.0090358357436871e-119, 32'sd-9.570053616298516e-123, 32'sd7.315226780970439e-122, 32'sd6.763118955287852e-120, 32'sd0.0033497528230176975, 32'sd0.013152464973132568, 32'sd0.03354874600002072, 32'sd-0.0018706833887496695, 32'sd0.032797487278599644, 32'sd-0.03938076702088776, 32'sd-0.002066374911142938, 32'sd0.013780710798400014, 32'sd-0.009132923830621304, 32'sd-0.03906534087756661, 32'sd-0.06115546907657194, 32'sd-0.022238949581161863, 32'sd0.03386345490451823, 32'sd0.08601863437708843, 32'sd-0.01924147746014512, 32'sd0.0002316763356512564, 32'sd0.016967846375269758, 32'sd-0.1271896414145591, 32'sd-0.02210698752545228, 32'sd-0.03718380599971299, 32'sd-2.7512269307603688e-114, 32'sd-4.1013091347413924e-117, 32'sd1.5130353796357538e-127, 32'sd-1.1386234895475597e-119},
        '{32'sd-4.6297941586851995e-115, 32'sd1.4106095724369526e-127, 32'sd1.3150672392046345e-117, 32'sd-1.5992292367248726e-127, 32'sd-4.7016820834011516e-126, 32'sd9.741649957149401e-119, 32'sd-1.8971914914028571e-125, 32'sd-4.847473107840543e-122, 32'sd1.0707601470558152e-123, 32'sd-1.686676676018178e-122, 32'sd3.5782404093294077e-127, 32'sd9.249369952943909e-120, 32'sd-0.07781036488693824, 32'sd-0.006464937262484267, 32'sd-0.04869568497644652, 32'sd-0.0021401225318786517, 32'sd-6.888114219731479e-124, 32'sd1.1091336556592306e-121, 32'sd-1.8102474871019154e-126, 32'sd-1.2825197651412896e-118, 32'sd4.266704387038475e-118, 32'sd1.7874725225121756e-122, 32'sd-7.830641008709954e-121, 32'sd-1.9998526935936863e-117, 32'sd2.0140242560374537e-124, 32'sd-1.710027110435499e-120, 32'sd4.42257126341604e-125, 32'sd2.2609266899348017e-122, 32'sd3.685826660500752e-119, 32'sd2.656450491697081e-121, 32'sd1.6312075822220742e-115, 32'sd1.0594431845819736e-117, 32'sd0.09453739057529455, 32'sd0.007381588433924106, 32'sd-0.024123729666991105, 32'sd0.051813650188370725, 32'sd0.03618175486201162, 32'sd-0.030693829941776034, 32'sd-0.12600145645929586, 32'sd-0.12456993710601376, 32'sd-0.04164286064516909, 32'sd-0.048181146044499586, 32'sd0.05146328574133705, 32'sd-0.08964605235150405, 32'sd-0.1559931915450466, 32'sd-0.009563740635035789, 32'sd-0.11493655735151642, 32'sd0.04156148418371539, 32'sd-0.00310664441359295, 32'sd0.062112315206184175, 32'sd0.015572236096661422, 32'sd-0.028936254981808216, 32'sd-4.765740093190477e-123, 32'sd3.6477258149219305e-116, 32'sd-8.453176187236721e-131, 32'sd3.165297579247264e-123, 32'sd-7.560746074419927e-127, 32'sd6.977847704224558e-128, 32'sd-0.02575501512027719, 32'sd-0.08643480905021765, 32'sd-0.005264211971728867, 32'sd-0.03612267908892033, 32'sd-0.012614193306574291, 32'sd0.03556561189701911, 32'sd0.05448321693349566, 32'sd0.025449289230967485, 32'sd-0.10742080627128732, 32'sd0.07916584650907918, 32'sd0.07422118599796994, 32'sd0.10409077789451031, 32'sd0.1625931002289048, 32'sd0.06922563884264164, 32'sd-0.0537085310389527, 32'sd-0.027651445460694906, 32'sd0.030109265964178525, 32'sd-0.1411930298281155, 32'sd-0.017955650795803912, 32'sd-0.02450408395867945, 32'sd0.046849684242830016, 32'sd0.029927047549332418, 32'sd0.02551921118363747, 32'sd0.015338141256100364, 32'sd9.293079483588868e-123, 32'sd2.97279970367804e-122, 32'sd2.1169086981056975e-119, 32'sd-1.0998382656549795e-121, 32'sd-0.04328631799847505, 32'sd0.018887262814401815, 32'sd0.01733372512254885, 32'sd-0.010497947104653063, 32'sd-0.0016329797575946549, 32'sd0.06209082388360358, 32'sd-0.028524562071324772, 32'sd-0.10790168462386257, 32'sd-0.06268339856907953, 32'sd0.08283210113234865, 32'sd-0.004300560947058788, 32'sd0.0964828096469836, 32'sd0.18033354794829579, 32'sd0.13803028307888157, 32'sd0.18402299827657223, 32'sd0.005046714209710759, 32'sd0.035565981616608074, 32'sd-0.011669548121170424, 32'sd0.08124855508700118, 32'sd0.10270778444368278, 32'sd0.0032781187071486695, 32'sd0.039367148660006526, 32'sd-0.04404267983800382, 32'sd-0.10884185890785086, 32'sd0.03406290766127998, 32'sd1.8725130500161363e-117, 32'sd-6.575018716829093e-120, 32'sd-0.011042558143767214, 32'sd0.0019147861721981261, 32'sd0.00732686024187807, 32'sd0.0019385013545313193, 32'sd0.033235609114577847, 32'sd0.03928488362890881, 32'sd0.04723570489423056, 32'sd-0.08216491886819767, 32'sd0.03165602410005078, 32'sd0.0794356884530698, 32'sd-0.07214844865443228, 32'sd0.03592399928107034, 32'sd-0.058848166215068706, 32'sd0.03675540943090341, 32'sd0.14020193376644258, 32'sd-0.024274141544210922, 32'sd0.025012955670711184, 32'sd0.032882101743786495, 32'sd0.003381407147821698, 32'sd0.02981677401668327, 32'sd0.17418442995249275, 32'sd-0.07152094668952236, 32'sd0.10474381720007658, 32'sd0.12665682703466266, 32'sd-0.019667964418552213, 32'sd-0.1955613702829432, 32'sd0.01444138818945155, 32'sd1.0512962979748886e-129, 32'sd0.01515304610548346, 32'sd-0.0003859983810695552, 32'sd0.06484578213218209, 32'sd0.06358295089419903, 32'sd-0.007930014651135794, 32'sd0.13123112269275233, 32'sd-0.016302985294819276, 32'sd-0.15999720457631217, 32'sd-0.054659576022988786, 32'sd-0.05269882378515865, 32'sd-0.08889526552608842, 32'sd0.06370576622132514, 32'sd0.10324824595717948, 32'sd-0.007438067653964951, 32'sd-0.06874790386128662, 32'sd-0.099321538508887, 32'sd0.08246193639431826, 32'sd0.07985763373956348, 32'sd0.03671515080826701, 32'sd0.014661596381857009, 32'sd0.07625122225526997, 32'sd-0.05253914376688267, 32'sd0.08367194962402764, 32'sd0.09409156551176467, 32'sd-0.09399919143606564, 32'sd-0.09108593875634101, 32'sd-0.031218544187079342, 32'sd-7.615153086609165e-127, 32'sd0.05199831515675857, 32'sd0.053022259546385335, 32'sd-0.004943094598422997, 32'sd0.04724560313979584, 32'sd-0.07286815922924773, 32'sd-0.03826111742405208, 32'sd-0.026611680032630366, 32'sd0.00014229401794823546, 32'sd-0.054696314440222535, 32'sd-0.11073024852836433, 32'sd0.04581485315013738, 32'sd-0.04029434020903927, 32'sd-0.05575564049439156, 32'sd-0.058873377456728354, 32'sd-0.06492486327777484, 32'sd-0.03473511345679187, 32'sd0.09008139728136608, 32'sd0.0066689269537673485, 32'sd-0.04889031957257495, 32'sd-0.014928824353913387, 32'sd-0.03357357468202596, 32'sd0.1080196474767366, 32'sd0.07637478143971607, 32'sd0.08084600217029235, 32'sd0.06825296791382528, 32'sd-0.034106021380757696, 32'sd-0.012577897527009945, 32'sd-0.032167073361327826, 32'sd0.03348980243560419, 32'sd0.0038779862156215167, 32'sd-0.057987934270145536, 32'sd-0.05821187859805512, 32'sd-0.13620544600587545, 32'sd-0.012986460423101365, 32'sd-0.09672696427723894, 32'sd-0.052508524051250526, 32'sd-0.12254429128084589, 32'sd-0.008190268188905583, 32'sd0.08065699582051847, 32'sd0.02890177362986581, 32'sd-0.07687547753073269, 32'sd0.0173428446418092, 32'sd0.04983607197057342, 32'sd0.0667617429363062, 32'sd0.10203604902027061, 32'sd-0.05858803905569207, 32'sd-0.1461912282492964, 32'sd-0.023405833283023376, 32'sd-0.057848617530202526, 32'sd0.1375371941401287, 32'sd-0.034990639846483707, 32'sd0.14410958032172452, 32'sd0.12288521612070254, 32'sd-0.08509164817685552, 32'sd-0.06882778967939963, 32'sd-0.03222082265832945, 32'sd0.045643358386641096, 32'sd-0.019061264102767088, 32'sd-0.1710711433547027, 32'sd-0.11170839962015586, 32'sd-0.12093120956078819, 32'sd0.03627364996386843, 32'sd-0.05744730266259238, 32'sd-0.04184288553236371, 32'sd-0.0014476947204516608, 32'sd-0.06600023173591525, 32'sd-0.12299770433687693, 32'sd-0.023916310079671856, 32'sd0.031589575229181314, 32'sd0.10686348105823552, 32'sd-0.027020904334334104, 32'sd0.07280697201269443, 32'sd-0.027010243984803964, 32'sd-0.07857139470921376, 32'sd-0.09049623914627157, 32'sd-0.15938063433542715, 32'sd-0.04040148967259757, 32'sd-0.10280631922945359, 32'sd-0.0609457330540141, 32'sd0.02659079776862363, 32'sd0.10355155492312765, 32'sd-0.0017176622068008878, 32'sd0.021269821635237374, 32'sd-0.011459858264031416, 32'sd0.0521493761632506, 32'sd0.04747362355472718, 32'sd-0.11945585223248792, 32'sd-0.01262480185284025, 32'sd0.017262575602069858, 32'sd0.022858629603085476, 32'sd0.004618043101994258, 32'sd-0.11318852615244468, 32'sd-0.1142782400538107, 32'sd-0.19041611767483166, 32'sd-0.06354158219337835, 32'sd0.08935299097706793, 32'sd0.0323799598728349, 32'sd-0.03962021831638573, 32'sd-0.11704719001185158, 32'sd0.045956860512299934, 32'sd0.06488430148693422, 32'sd-0.05156817035172996, 32'sd0.021912827286903174, 32'sd-0.0647736835785223, 32'sd0.07765591169095343, 32'sd-0.1652191653501355, 32'sd-0.08379892355885624, 32'sd-0.08858313131910611, 32'sd0.038214921488749956, 32'sd-0.08949367782149562, 32'sd-0.06488849214225986, 32'sd-0.027368957259399865, 32'sd0.04844770101175204, 32'sd-0.05522809288863464, 32'sd0.006181780271101413, 32'sd0.09249752794156933, 32'sd0.15149372095150473, 32'sd0.044265088461139274, 32'sd-0.021487643054518897, 32'sd-0.07431057650884944, 32'sd0.020974232771565914, 32'sd-0.0634890320156808, 32'sd-0.05761038562538055, 32'sd-0.08283794977521844, 32'sd-0.1397401182621715, 32'sd-0.0931683445247105, 32'sd-0.1818450903794426, 32'sd-0.08866386636238481, 32'sd-0.050082029814558456, 32'sd-0.02893756233645006, 32'sd-0.0553537413346856, 32'sd-0.09771081021641143, 32'sd-0.07943486071833479, 32'sd-0.12890307147572672, 32'sd-0.04813243651934079, 32'sd-0.0005097246882310396, 32'sd-0.012986767351477175, 32'sd-0.042528768076404364, 32'sd-0.007615632076815943, 32'sd-0.046439819174056436, 32'sd-0.0012575499116689278, 32'sd0.05667904161236499, 32'sd0.07314620185201114, 32'sd-0.0331243269092401, 32'sd-0.02182849226979256, 32'sd0.11485246411681418, 32'sd0.08323804105900115, 32'sd0.07156531887972055, 32'sd-0.0030549469002255883, 32'sd-0.016621848523062442, 32'sd-0.06625010883824112, 32'sd-0.19586961732070401, 32'sd-0.2633735817228527, 32'sd-0.17643080408762424, 32'sd-0.14309413569476945, 32'sd-0.06749305620286136, 32'sd-0.07992742545232993, 32'sd-0.033822709883584115, 32'sd-0.008261670282446544, 32'sd0.06603032292328925, 32'sd-0.019224605057967435, 32'sd-0.18228385259386962, 32'sd-0.1258540347239649, 32'sd-0.16272257121663714, 32'sd-0.0997408482428582, 32'sd-0.06743031509972376, 32'sd-0.04733123543214667, 32'sd0.003289684025130058, 32'sd-0.04329414355980569, 32'sd0.018614342747152273, 32'sd-0.0317992785470977, 32'sd-0.043302902793383474, 32'sd0.039643942910608694, 32'sd0.08807932073267488, 32'sd-0.03869245941861964, 32'sd0.05901208668499676, 32'sd0.01965075332274631, 32'sd0.13688506539290687, 32'sd-0.04999703852796389, 32'sd-0.15804402898332648, 32'sd-0.12819318162248802, 32'sd-0.10906988873072022, 32'sd-0.10751174989413854, 32'sd-0.034900356605906395, 32'sd-0.0775353350679953, 32'sd0.03800454140654046, 32'sd0.04146813322491193, 32'sd-0.10391743506475458, 32'sd-0.13086259601400155, 32'sd-0.03482902671133486, 32'sd0.017437239179585798, 32'sd-0.009891452990926518, 32'sd0.06768544969297924, 32'sd0.011683654481724846, 32'sd-0.060610937291585794, 32'sd0.009071454104562095, 32'sd0.03362038426326272, 32'sd-0.05882198642398084, 32'sd0.08018887695160076, 32'sd-0.02366782651853718, 32'sd-0.07025402996380314, 32'sd0.04754042842250362, 32'sd-0.02071850871395986, 32'sd0.0047584560873957515, 32'sd0.1472780195701832, 32'sd0.2569385662787918, 32'sd0.07086225951132609, 32'sd-1.9216059702502924e-05, 32'sd-0.07838488270443034, 32'sd-0.055794486089596064, 32'sd-0.06971669530140677, 32'sd0.1160176061024269, 32'sd0.007301436056987871, 32'sd-0.09321077330234823, 32'sd0.023336897745206153, 32'sd-0.03361222297301813, 32'sd-0.07268969083464463, 32'sd-0.0568805279969852, 32'sd-0.11885882569832902, 32'sd0.009830014804179773, 32'sd-0.07659411871450576, 32'sd0.032099498642063885, 32'sd-0.0019625078691462242, 32'sd0.006003393516543059, 32'sd0.008705935245455121, 32'sd0.017988932823072235, 32'sd0.07931044362325775, 32'sd-0.059459907227632926, 32'sd0.0011819685186462202, 32'sd0.08484804293092872, 32'sd0.02144918248308455, 32'sd0.05034892562253159, 32'sd0.018256345950706732, 32'sd0.07571259006126854, 32'sd0.09618433362329847, 32'sd0.12083203516417662, 32'sd0.1310998094616179, 32'sd0.030161223672488226, 32'sd0.03680379108002908, 32'sd0.1005894067811378, 32'sd0.08505828806120717, 32'sd-0.06941825944994008, 32'sd-0.06110413745473872, 32'sd-0.1331500437440967, 32'sd-0.07299339507862157, 32'sd-0.056432513538418265, 32'sd-0.027206356145502677, 32'sd-0.03912989002787317, 32'sd0.007880626457573382, 32'sd0.05575386344542672, 32'sd-0.03582997789703694, 32'sd-0.048746674107187166, 32'sd-0.022695565546527047, 32'sd-0.06668199421921184, 32'sd0.0803396864453166, 32'sd0.002135544132890572, 32'sd0.005772171227852098, 32'sd0.06756813078476229, 32'sd0.08260701975108493, 32'sd0.09228243166201053, 32'sd0.05276843526559199, 32'sd0.057254613356106175, 32'sd0.048706065477356335, 32'sd0.11804896198373127, 32'sd0.12873265136410178, 32'sd0.0943856230375377, 32'sd0.15070189337794643, 32'sd0.20815003408996313, 32'sd-0.010775147821285767, 32'sd-0.10429263462351648, 32'sd-0.062415827296620596, 32'sd-0.13987081085414674, 32'sd-0.051036401850707076, 32'sd0.05992699504353351, 32'sd0.05240592307521507, 32'sd0.044930285171895276, 32'sd-0.03784626805147346, 32'sd0.012234175220660335, 32'sd-0.010503993304419944, 32'sd0.049948999058588475, 32'sd0.035266798050039544, 32'sd-0.0056477503616067844, 32'sd0.012082256175580439, 32'sd0.02921515307134818, 32'sd0.04789284388746117, 32'sd0.15156970469772327, 32'sd0.17058205517620964, 32'sd0.1522641879601995, 32'sd0.07860084543045126, 32'sd0.03970247499493364, 32'sd0.11593636833507842, 32'sd0.2323238157703704, 32'sd0.16030048882124234, 32'sd-0.017348114274361698, 32'sd0.08639675032903683, 32'sd0.08622558674534765, 32'sd0.09036627368021949, 32'sd-0.049781277441938006, 32'sd0.034702531516070674, 32'sd-0.0038840957799543903, 32'sd-0.07055185238168679, 32'sd0.020790292120243622, 32'sd-0.020464744411997676, 32'sd-0.0276561426993146, 32'sd0.003092055579750906, 32'sd0.05021098694232478, 32'sd0.00863501741709157, 32'sd1.775239710215065e-123, 32'sd0.06537279602251124, 32'sd0.01149562788884564, 32'sd0.10143944906075231, 32'sd-0.06748059930526952, 32'sd0.0275630877555991, 32'sd0.04810302229350316, 32'sd0.05460286020053189, 32'sd0.05950122980918815, 32'sd0.1234137302738968, 32'sd0.2157773155772312, 32'sd0.09194588989331738, 32'sd0.16260712079234896, 32'sd0.057968318750854474, 32'sd-0.03086405845395254, 32'sd-0.005518152160511978, 32'sd0.06459927786616303, 32'sd0.04382998001076306, 32'sd-0.12277459561347634, 32'sd-0.014515160721255223, 32'sd-0.046454704717315984, 32'sd0.029443656024195516, 32'sd-0.0805009756921665, 32'sd-0.03972531205181198, 32'sd0.05502637403129064, 32'sd-0.015984696694117, 32'sd-0.03802185466051911, 32'sd-0.04757386982281618, 32'sd-0.0026061095066167903, 32'sd-0.1012543934868637, 32'sd-0.08811840236837946, 32'sd0.07003882337110771, 32'sd-0.04845570641030268, 32'sd-0.17004379138109382, 32'sd-0.03096035646179631, 32'sd0.1021819295824631, 32'sd0.1889757513249384, 32'sd0.17442234122032577, 32'sd0.010681572209676488, 32'sd0.12911096554041396, 32'sd0.14541008087168486, 32'sd0.12756254892407304, 32'sd-0.053741078454384306, 32'sd0.07294019815737177, 32'sd0.024336600707979043, 32'sd0.016765162391492165, 32'sd-0.05114516483795899, 32'sd-0.07845940951414634, 32'sd-0.06003479860760887, 32'sd-0.03385821925750722, 32'sd-0.017511695774800974, 32'sd0.03769436085634716, 32'sd0.10834229479899796, 32'sd0.10225003193324855, 32'sd-0.16440542285850973, 32'sd-0.058694692220834295, 32'sd0.05369349535108508, 32'sd-0.04884590107449849, 32'sd-0.1225991831203311, 32'sd0.04417271903957183, 32'sd0.09470695213440657, 32'sd-0.021227181908727438, 32'sd-0.12698788793809393, 32'sd-0.05237964234449355, 32'sd-0.04851510535617479, 32'sd-0.05653715250355692, 32'sd-0.08753599301983016, 32'sd-0.0429488805198771, 32'sd0.10334740181515517, 32'sd0.08859760863345242, 32'sd0.024494144257664007, 32'sd0.005047952295988828, 32'sd0.04292771231457077, 32'sd0.12639898803623134, 32'sd-0.007333056424495475, 32'sd-0.02595707811872226, 32'sd-0.11322818121148202, 32'sd0.051435422648275254, 32'sd-0.013449527973624762, 32'sd0.02297933799502699, 32'sd0.0829718004509007, 32'sd0.053507179290584704, 32'sd0.0064440341792824435, 32'sd-0.07165176548262553, 32'sd3.8793624547786746e-125, 32'sd0.046334209472639463, 32'sd0.03960117774514167, 32'sd0.0031479610064691515, 32'sd-0.1668042598206007, 32'sd-0.13977187953849535, 32'sd-0.09975760945188104, 32'sd-0.035089477882360665, 32'sd-0.0037261598276939483, 32'sd0.01849560863432822, 32'sd-0.1393433454567541, 32'sd-0.08224688199824949, 32'sd-0.05887386887445116, 32'sd0.06805645077446848, 32'sd0.0777779569701611, 32'sd0.010124829624763548, 32'sd-0.0511133454530921, 32'sd0.10010216020915841, 32'sd0.13007295466054275, 32'sd-0.05203857340472038, 32'sd0.05407853411291561, 32'sd0.028384532889961997, 32'sd0.05941878734653629, 32'sd-0.08143192101139887, 32'sd0.025708508749670605, 32'sd-0.03195722740096397, 32'sd-0.006583021599410211, 32'sd0.024539166703964006, 32'sd-0.04198069068396032, 32'sd0.08622580815628093, 32'sd0.012374508283806054, 32'sd-0.010792795919502522, 32'sd-0.12563960075319078, 32'sd-0.059250263834687, 32'sd-0.07838476256289724, 32'sd-0.10817060628604779, 32'sd-0.022444142432713855, 32'sd0.0019078243114028961, 32'sd-0.027357566457524084, 32'sd-0.09173804749424695, 32'sd-0.054479244460324025, 32'sd0.13363131625760732, 32'sd-0.04626121501121352, 32'sd0.06847871178502037, 32'sd-0.010221996067340625, 32'sd0.12727378110731202, 32'sd0.14195100470626618, 32'sd0.011962295238718133, 32'sd0.004683052259721946, 32'sd-0.05106947716893374, 32'sd0.08014391797991614, 32'sd0.016448951226345702, 32'sd-0.10851109714023272, 32'sd-0.0858040671270105, 32'sd-0.05262787557481366, 32'sd0.03782852880613336, 32'sd0.013153426745948958, 32'sd-0.007324102822833622, 32'sd0.008490204666078808, 32'sd0.08859711356587897, 32'sd0.02664456997651075, 32'sd-0.030390348145114984, 32'sd-0.21581395280544668, 32'sd-0.15880473038487808, 32'sd-0.12183286288310596, 32'sd0.004468425976773402, 32'sd0.027540014428856667, 32'sd0.038945662836765246, 32'sd-0.02002665314949798, 32'sd-0.0005598204842699285, 32'sd-0.06019866007427211, 32'sd0.10217390868746885, 32'sd0.18601734782752016, 32'sd0.04212580317525311, 32'sd0.16846919149273648, 32'sd0.0965450321816863, 32'sd0.11100709707950975, 32'sd0.08670009936431426, 32'sd0.02753267390007012, 32'sd-0.14584854733967748, 32'sd-0.04336571538101943, 32'sd-0.07289876557198148, 32'sd0.022381019508297437, 32'sd-0.017743370668313885, 32'sd4.246983721848622e-121, 32'sd0.06695858131598478, 32'sd-0.029101204538956163, 32'sd0.11538926611368741, 32'sd0.04092358767829025, 32'sd0.006193866414261251, 32'sd-0.05162823649312605, 32'sd-0.21923410148331812, 32'sd-0.03608429248533859, 32'sd-0.04075046606515015, 32'sd0.05496072218238208, 32'sd-0.014396604839100798, 32'sd-0.06987874288821959, 32'sd-0.12345056361606237, 32'sd0.018650339360238063, 32'sd0.1203282194219444, 32'sd-0.01971588507301023, 32'sd0.07175915339016746, 32'sd0.08878271621017755, 32'sd0.1089248423334243, 32'sd0.050404788554746505, 32'sd0.06246822374434035, 32'sd-0.010471781816130333, 32'sd-0.022533207886767864, 32'sd-0.02022610686320697, 32'sd-0.09002287239243449, 32'sd-0.023083208960389803, 32'sd-5.485906747378311e-124, 32'sd6.7021922918541306e-127, 32'sd-3.495104945149166e-122, 32'sd-0.061603503911534685, 32'sd-0.04231386388699802, 32'sd-0.14097795897946364, 32'sd-0.09531232561072792, 32'sd0.02497780632075025, 32'sd-0.008729669048788464, 32'sd0.06530306094211549, 32'sd-0.01627206404993918, 32'sd-0.01615053234130029, 32'sd0.15428994017938424, 32'sd-0.022821970018065425, 32'sd0.07022098356403361, 32'sd0.09566902603157294, 32'sd-0.025850623098622107, 32'sd0.029904999556944468, 32'sd-0.11723915981809352, 32'sd-0.02292533013729025, 32'sd0.0902659604379013, 32'sd0.14969871325878228, 32'sd-0.03902635128277502, 32'sd-0.008013971908078978, 32'sd0.06492336067349834, 32'sd-0.09451723292444862, 32'sd0.014401580078967332, 32'sd0.05523010927100406, 32'sd-7.408043009839419e-118, 32'sd3.0487898748521816e-124, 32'sd-5.954611173190094e-125, 32'sd-0.030218398992368677, 32'sd-0.032650323175229395, 32'sd-0.05312454473191595, 32'sd0.0656297885126433, 32'sd-0.02671001912666308, 32'sd-0.0010847890560446165, 32'sd-0.07652756299074413, 32'sd0.02064797243032818, 32'sd-0.055350621757596676, 32'sd0.04838119227985096, 32'sd0.16201424534869993, 32'sd0.10472098004820192, 32'sd-0.09741522042639585, 32'sd-0.09566586093035553, 32'sd-0.12445956355207675, 32'sd-0.11754955774643645, 32'sd0.03885588326520841, 32'sd0.11125889703341536, 32'sd0.07117823227527517, 32'sd-0.07954458590676139, 32'sd-0.03514162837998294, 32'sd-0.06753711972971907, 32'sd-0.01560190188152464, 32'sd0.07928931709947545, 32'sd0.01956806205997161, 32'sd-2.560680750705505e-120, 32'sd-1.142987267347651e-123, 32'sd2.3594790498369915e-118, 32'sd-8.615622230110274e-126, 32'sd0.020095601842587497, 32'sd0.04376892421452022, 32'sd0.03994876685936016, 32'sd0.0919834562317019, 32'sd0.03536153383068195, 32'sd0.003094009941691667, 32'sd-0.052901999929997084, 32'sd-0.11935855281649835, 32'sd0.030354899256468955, 32'sd0.05760739113926329, 32'sd0.09296807218162824, 32'sd0.057673962309365605, 32'sd0.02872347047416432, 32'sd0.011602211415959029, 32'sd-0.10870912002230171, 32'sd-0.010725096321717946, 32'sd-0.031262356605932705, 32'sd-0.05200096498135348, 32'sd0.047248006711638625, 32'sd0.04647813289892214, 32'sd-0.01971661269978226, 32'sd0.08105189910555077, 32'sd-0.03152047992574606, 32'sd9.659587974363775e-122, 32'sd4.0586418578243103e-115, 32'sd-4.167683499824437e-118, 32'sd2.940787819145885e-121, 32'sd1.0924048960528752e-121, 32'sd-1.2993719922276303e-125, 32'sd-0.0402085828019228, 32'sd-0.044459957772449855, 32'sd-0.036593271337358554, 32'sd0.053266241217720035, 32'sd0.07022209436257439, 32'sd-0.00649230007484732, 32'sd0.04363036389838075, 32'sd0.048483750933026024, 32'sd0.09233137404595612, 32'sd0.007855676213710465, 32'sd0.0617321232955392, 32'sd0.0465468637833321, 32'sd0.0057080658723181535, 32'sd-0.01506555936833644, 32'sd-0.06744598196017601, 32'sd0.028624539028130568, 32'sd0.05163211548448608, 32'sd0.04067016573418661, 32'sd0.03360441044604608, 32'sd0.0005655325284959753, 32'sd1.8433888295200474e-120, 32'sd-4.674645066405005e-118, 32'sd-4.914367719594069e-120, 32'sd-7.348494013207921e-115},
        '{32'sd1.640079518399767e-116, 32'sd4.311414554410861e-125, 32'sd-1.3611581143330544e-126, 32'sd-8.61713267948596e-117, 32'sd-3.403782891747188e-125, 32'sd-4.766617931593875e-126, 32'sd1.0245743846416209e-115, 32'sd-3.289410324429303e-121, 32'sd-1.3221951878250814e-124, 32'sd-3.0158090737704277e-120, 32'sd2.183680201630986e-122, 32'sd-2.1362294002061042e-122, 32'sd0.133073787070603, 32'sd0.05979700745184205, 32'sd0.1002764569535098, 32'sd0.03705655299184246, 32'sd-3.735093522930128e-120, 32'sd-3.3890393287202e-122, 32'sd-2.1179993235250936e-119, 32'sd-1.0333352927850474e-116, 32'sd1.0768907895658592e-124, 32'sd-3.6401904901742593e-122, 32'sd9.906850318488642e-123, 32'sd9.61311545379454e-123, 32'sd5.298436991930494e-118, 32'sd-2.3871889963749115e-122, 32'sd-7.589202516718341e-126, 32'sd6.524879189045635e-126, 32'sd1.069489677224011e-121, 32'sd-2.9625222233393252e-118, 32'sd3.6298594128180227e-115, 32'sd3.766046315207982e-126, 32'sd0.027101206775146106, 32'sd0.027285498163683513, 32'sd-0.004472685285863839, 32'sd0.14961199642404752, 32'sd0.1350617911573765, 32'sd0.06959261192066238, 32'sd0.012951108437085487, 32'sd0.042308963496269864, 32'sd0.11249772610493218, 32'sd0.05032607444322446, 32'sd-0.005377380892304511, 32'sd0.06398373407634618, 32'sd0.047767849576857514, 32'sd0.0010672146773690004, 32'sd-0.0827861692219993, 32'sd0.05346520021158061, 32'sd0.05005395816039865, 32'sd0.09800819403248281, 32'sd0.024264070092080887, 32'sd0.01889430772626745, 32'sd1.3916945487371956e-127, 32'sd3.85198522695809e-115, 32'sd1.2155881958276004e-117, 32'sd1.73264820257255e-125, 32'sd6.782678751111303e-124, 32'sd4.1277080072332707e-122, 32'sd0.05280787425482569, 32'sd0.0910922888426257, 32'sd0.0003876792105961591, 32'sd-0.0046401644616196076, 32'sd0.0598528114636204, 32'sd-0.02704293543393837, 32'sd0.10906125112909686, 32'sd0.13175681288352165, 32'sd0.0196024869942899, 32'sd0.02313265752166656, 32'sd0.09456301657438736, 32'sd0.0821446373234339, 32'sd0.04304798626462648, 32'sd0.08881918904111832, 32'sd0.059805276115329445, 32'sd0.102226053526293, 32'sd0.026865535472362326, 32'sd0.03269762464940796, 32'sd0.08390902486838679, 32'sd0.07721491205651214, 32'sd0.08000402668842313, 32'sd0.07090832694293506, 32'sd-0.010725147500540115, 32'sd0.08307619102839175, 32'sd3.1108364769100204e-125, 32'sd2.6843144796899164e-124, 32'sd8.126915528722594e-122, 32'sd6.277941732682105e-119, 32'sd0.07458549380796765, 32'sd0.0993406587914086, 32'sd0.03646616834052056, 32'sd0.026400396145668494, 32'sd-0.00030983404523518874, 32'sd0.1081667201118406, 32'sd0.08152048146101133, 32'sd0.15821297743032756, 32'sd0.0015968639185127216, 32'sd0.07862868244092501, 32'sd-0.09381110414208006, 32'sd0.030187322903038043, 32'sd0.030048793268652885, 32'sd-0.01736715778072254, 32'sd0.008752088707287732, 32'sd-0.07567476667621041, 32'sd-0.09717523225709702, 32'sd-0.10155763645251226, 32'sd-0.13804806994761343, 32'sd0.027994368919003393, 32'sd-0.05670444297300537, 32'sd0.028351798287783267, 32'sd0.015771944970178895, 32'sd0.007677692870182676, 32'sd0.09985004137833152, 32'sd2.3847564829251327e-124, 32'sd5.415352633410414e-115, 32'sd0.0469601128601678, 32'sd0.06391249629759164, 32'sd-0.01887556464845246, 32'sd0.047992771504027754, 32'sd0.07962545682860342, 32'sd-0.056700555607219136, 32'sd0.020116115973670072, 32'sd0.04650578512183264, 32'sd-0.03310316100740729, 32'sd0.06328433548597603, 32'sd-0.07185458702897571, 32'sd0.018589750439259613, 32'sd-0.08023035547083207, 32'sd-0.0122156734265321, 32'sd0.08231960516052798, 32'sd0.11348203947287723, 32'sd0.029327648443221017, 32'sd-0.057388190332168985, 32'sd-0.013058666711255938, 32'sd-0.0014331769100306953, 32'sd0.031459579658820125, 32'sd0.15751865371869853, 32'sd-0.030965679327883258, 32'sd-0.061687150843999186, 32'sd-0.12216420491793409, 32'sd0.04361011934747563, 32'sd0.0363935949058683, 32'sd1.1988448347169176e-122, 32'sd0.07124639846562715, 32'sd-0.08811179382283008, 32'sd0.02577878348513496, 32'sd0.08126125758518475, 32'sd-0.0020655275427055144, 32'sd-0.014969708364300529, 32'sd0.017113872923585623, 32'sd0.023870593608693355, 32'sd-0.04541584404074478, 32'sd-0.1691171623385157, 32'sd-0.13204433962708248, 32'sd-0.054279067377346495, 32'sd-0.12751759691436002, 32'sd0.0035834481755374053, 32'sd0.022075721143662422, 32'sd-0.008551908995530414, 32'sd0.05397295501742701, 32'sd-0.10102407449860538, 32'sd-0.030961030548316778, 32'sd-0.013392875314751616, 32'sd0.046941562129666534, 32'sd0.09901851606573345, 32'sd0.17099049073261952, 32'sd-0.0776182100427041, 32'sd-0.021482314148289897, 32'sd-0.19875510478491754, 32'sd0.0029739932679217073, 32'sd-3.673672021338075e-116, 32'sd0.04137163894516794, 32'sd-0.0003015670062110312, 32'sd-0.0693416622784735, 32'sd0.036604803205580294, 32'sd0.09252441692718164, 32'sd0.04943167418546383, 32'sd0.0866997932180474, 32'sd0.1647710232317891, 32'sd0.05117489084711875, 32'sd-0.23706364791263784, 32'sd-0.12431014517179452, 32'sd-0.19477007714997235, 32'sd-0.24162927350274063, 32'sd-0.15385672280819865, 32'sd-0.02363802348760945, 32'sd0.0485995563070802, 32'sd-0.02324543140213992, 32'sd0.03437710586355476, 32'sd0.021481042089348534, 32'sd-0.024745825272461476, 32'sd-0.013682557313231019, 32'sd0.008563314559683429, 32'sd-0.036740131430022284, 32'sd0.03767274681408896, 32'sd-0.048250800417729854, 32'sd0.020966718530581387, 32'sd-0.07836529933369367, 32'sd0.11308774938457422, 32'sd-0.07940300948769165, 32'sd-0.10215689693243954, 32'sd-0.009355116268755934, 32'sd0.06974812913747405, 32'sd0.010925600156490748, 32'sd0.0002069345028828234, 32'sd0.016451833775116248, 32'sd0.02475713899494597, 32'sd-0.15101266882077544, 32'sd-0.13664846473532888, 32'sd-0.15632728790411896, 32'sd-0.11685907537090917, 32'sd-0.11922017658479062, 32'sd-0.06892267087884049, 32'sd0.013824938118598059, 32'sd0.12940658825461301, 32'sd-0.013943597624311351, 32'sd-0.14344881116445837, 32'sd0.13867325797335503, 32'sd0.10399284167338446, 32'sd0.0019491258633138042, 32'sd-0.09246356317953462, 32'sd-0.043625570561863516, 32'sd-0.01554639209788226, 32'sd-0.025641389590427617, 32'sd0.008795584214850048, 32'sd0.041518833289648525, 32'sd-0.012896279995296099, 32'sd-0.061335668361304954, 32'sd-0.014014275169458391, 32'sd-0.058659027594660955, 32'sd0.05319862831569931, 32'sd-0.019956990759701313, 32'sd0.12968564033832383, 32'sd0.00570185405909212, 32'sd-0.0037128838193597534, 32'sd-0.10910261637509241, 32'sd-0.05152555949674608, 32'sd-0.03530011720739054, 32'sd-0.03511466047943039, 32'sd-0.10725952845155036, 32'sd0.12881199626663972, 32'sd0.013893497449848451, 32'sd0.061640893591060994, 32'sd-0.08736946226745275, 32'sd-0.06838039771164478, 32'sd0.08538218354153636, 32'sd0.047103073582504255, 32'sd-0.01906944455420026, 32'sd-0.05045517293160877, 32'sd-0.13520718062168582, 32'sd0.004110498097110213, 32'sd-0.001920395053928028, 32'sd0.05142304392380966, 32'sd0.06410087258351449, 32'sd0.04269672394981501, 32'sd-0.004031627588489348, 32'sd0.0016378677960400994, 32'sd0.007982240858867826, 32'sd0.02084190881279486, 32'sd0.020543809297657565, 32'sd0.1026762053608207, 32'sd0.04294313989811178, 32'sd-0.03992738797614429, 32'sd0.001579027569591236, 32'sd0.067419200002036, 32'sd-0.09286337607972107, 32'sd-0.10393901184303243, 32'sd-0.1539311879301524, 32'sd0.012083425774176253, 32'sd0.0781066251477933, 32'sd0.08860794558734716, 32'sd-0.03782191735412064, 32'sd-0.08488233963095056, 32'sd-0.0433385195124518, 32'sd-0.05468866588510533, 32'sd0.09149701626321709, 32'sd-0.0857037035851144, 32'sd-0.04264503741510351, 32'sd-0.045128593067517216, 32'sd-0.004075889815283914, 32'sd0.047266517054167984, 32'sd0.07597674918350487, 32'sd0.015633355313802437, 32'sd0.0851878917451399, 32'sd-0.06653296630946139, 32'sd-0.011727168614114257, 32'sd-0.03642720068007177, 32'sd0.019626359340345918, 32'sd-0.033149867588464346, 32'sd0.031483244524283936, 32'sd-0.057053399653600595, 32'sd0.05222278566847917, 32'sd0.020464908614076897, 32'sd-0.11113926839504024, 32'sd-0.20621484411928445, 32'sd-0.08810193871236803, 32'sd-0.001394847335351589, 32'sd0.06701226326138668, 32'sd-0.019155656296035894, 32'sd-0.028160273504017255, 32'sd-0.02396373065417713, 32'sd-0.012073504270478578, 32'sd-0.11705602634477522, 32'sd-0.007287361324695098, 32'sd-0.01468143073259783, 32'sd-0.05659325798082357, 32'sd-0.01578206906960684, 32'sd-0.06180133115815641, 32'sd-0.04694531481422763, 32'sd0.0784765543283434, 32'sd0.00021914665128770108, 32'sd0.009020868830294914, 32'sd0.04462005639484912, 32'sd-0.01333197013404467, 32'sd0.023132894392971972, 32'sd-0.06960012251014802, 32'sd0.04456168674310161, 32'sd-0.05758954156465331, 32'sd0.0866532433887056, 32'sd0.18595498519401438, 32'sd0.039562992876228865, 32'sd-0.0969950935430148, 32'sd-0.13004624779851076, 32'sd-0.15454320260609808, 32'sd0.04576534444520709, 32'sd-0.03347232151321131, 32'sd0.047747837047838096, 32'sd-0.13854234718026198, 32'sd-0.10202177555423803, 32'sd0.04197652750147716, 32'sd-0.1370364519967906, 32'sd-0.022689787942024184, 32'sd-0.11966524807186191, 32'sd0.05491495096432997, 32'sd-0.1245480444450734, 32'sd-0.041798478034329, 32'sd0.021768161059736627, 32'sd-0.001342494370764471, 32'sd0.049895144819605594, 32'sd-0.02403947562824349, 32'sd0.04913431588470642, 32'sd0.025235607697338763, 32'sd-0.015152372751872378, 32'sd0.007669449165110889, 32'sd-0.06891214664964321, 32'sd-0.0027096956087215786, 32'sd0.11358059971845602, 32'sd0.0990960530621688, 32'sd0.03300653422196764, 32'sd-0.09685360005927728, 32'sd0.055435992066673136, 32'sd-0.010939194398980277, 32'sd-0.021173069023371845, 32'sd-0.05758738420676154, 32'sd0.010666686614067453, 32'sd-0.06658390252629458, 32'sd-0.007552544236140566, 32'sd-0.0484835985258454, 32'sd-0.0643300501939768, 32'sd-0.02222587697826886, 32'sd-0.009611988350070187, 32'sd-0.044287600400309775, 32'sd-0.06529090627067172, 32'sd0.04100515788972107, 32'sd-0.045389146965861084, 32'sd-0.003290739743664521, 32'sd0.03228736580946728, 32'sd0.02186648389478206, 32'sd-0.0068841750018260916, 32'sd-0.10448972121075978, 32'sd-0.12725715689043035, 32'sd-0.020872196504476075, 32'sd-0.07988701891400816, 32'sd0.0817110822202509, 32'sd0.09629013450136478, 32'sd0.20734603002832733, 32'sd0.13395492591362498, 32'sd-0.04372843163683649, 32'sd0.014098593436181582, 32'sd-0.061012112934188484, 32'sd-0.0438931881917671, 32'sd0.11687047584835675, 32'sd0.0025139091681294, 32'sd0.019036228340489913, 32'sd0.06266283307812935, 32'sd-0.044500787277178044, 32'sd-0.08375830457956346, 32'sd-0.029229568070978925, 32'sd0.005094264136834772, 32'sd-0.013390242625523055, 32'sd-0.029918333872693062, 32'sd-0.02695702524067569, 32'sd-0.022298079282487684, 32'sd0.10318834887042293, 32'sd0.06263559815678739, 32'sd0.0219040263097978, 32'sd0.03335647696897702, 32'sd0.02471809735139073, 32'sd-0.05463906550276617, 32'sd-0.03316005952498127, 32'sd-0.06276358477223373, 32'sd0.0032437464338439773, 32'sd0.10435375132548684, 32'sd0.05741645774886764, 32'sd0.06996979743813068, 32'sd-0.038615734975749515, 32'sd-0.10316814343921889, 32'sd-0.03163322443250708, 32'sd0.1310334024874171, 32'sd0.08058745992986638, 32'sd0.16093208335483, 32'sd0.028708695006634626, 32'sd0.0314311493077506, 32'sd0.005204640747855232, 32'sd-0.030272015158353018, 32'sd-0.12604201178249874, 32'sd-0.037696999175765716, 32'sd-0.008272547011797386, 32'sd0.08083847213494058, 32'sd-0.024949028335331646, 32'sd0.02687897639770179, 32'sd0.15870591249599195, 32'sd-0.07733786848121402, 32'sd0.057571501694898046, 32'sd-0.010532092705879743, 32'sd0.045610267876561784, 32'sd0.0066364923531264455, 32'sd0.10562542451681575, 32'sd-0.003552647322628455, 32'sd-0.006524348941708732, 32'sd0.06740804190344339, 32'sd0.03745063122178077, 32'sd0.008036497828696974, 32'sd-0.06697764865945452, 32'sd-0.08865868490167457, 32'sd0.0063682364506693545, 32'sd0.11491870711073565, 32'sd-0.02699018572344451, 32'sd0.0703928712334902, 32'sd0.07652727005631302, 32'sd0.007967027959359583, 32'sd-0.08912663826189762, 32'sd0.07572958295946701, 32'sd-0.06385425827165178, 32'sd0.02479664660999119, 32'sd0.07275248212709265, 32'sd0.07732017750526414, 32'sd-0.11096437150477002, 32'sd-0.13528369697666012, 32'sd0.0794934713481646, 32'sd0.027136135257531627, 32'sd-0.09675973835846137, 32'sd-0.015058561356898655, 32'sd-0.02410905549311607, 32'sd-0.07055425545422428, 32'sd0.00669721498128863, 32'sd-0.011702680103636374, 32'sd-0.018405545801339653, 32'sd-0.001369943795293368, 32'sd0.02244753905521141, 32'sd0.030686466630506393, 32'sd-0.02723696736004879, 32'sd0.011223545206370878, 32'sd0.008751051035191441, 32'sd-0.05299767365897972, 32'sd0.16149185902326466, 32'sd0.13017126811965324, 32'sd-0.015167921370959625, 32'sd0.033061317564374325, 32'sd-0.007438263921501843, 32'sd0.04675402532463377, 32'sd0.06935991408066854, 32'sd0.03614592332378071, 32'sd-0.027904189197221776, 32'sd0.02943560875344629, 32'sd0.07439809024860092, 32'sd0.008288250935344495, 32'sd0.06913477607499154, 32'sd2.518567060650645e-121, 32'sd-0.05632244844047593, 32'sd-0.021535073839027294, 32'sd-0.049218902209932476, 32'sd5.421243585742523e-05, 32'sd0.07926112484368904, 32'sd-0.03569818760774969, 32'sd0.026194080072712036, 32'sd0.05999674187681422, 32'sd-0.12159525757741864, 32'sd-0.022096334024067375, 32'sd-0.08395192520934139, 32'sd-0.07744274781708772, 32'sd0.017868197490026935, 32'sd0.11516850635416963, 32'sd0.17651884344830235, 32'sd0.1666698624094347, 32'sd0.014014368018780862, 32'sd-0.04964913872201173, 32'sd-0.10971474003232129, 32'sd-0.14695417739473887, 32'sd-0.040664045738619016, 32'sd0.15117281519381662, 32'sd0.014373477951547206, 32'sd-0.09380542167106413, 32'sd-0.027600582503566763, 32'sd-0.05999080359138831, 32'sd-0.029794996967995032, 32'sd0.044639509417858346, 32'sd0.05903056053019521, 32'sd-0.10353328099923507, 32'sd0.10194978990474533, 32'sd-0.03008716051168502, 32'sd-0.006198281231419645, 32'sd-0.1032043552601324, 32'sd-0.035721858530235455, 32'sd0.0035611956586593875, 32'sd0.01838551228393072, 32'sd-0.0470310703217083, 32'sd-0.008476207848187898, 32'sd0.09046795623954146, 32'sd0.09724647043751954, 32'sd0.1850039910203819, 32'sd0.09088814447077535, 32'sd-0.013949575395248902, 32'sd0.01232185702889908, 32'sd-0.030207433465051815, 32'sd-0.0627108704323838, 32'sd-0.10804087551718816, 32'sd-0.09376538622147518, 32'sd0.04442868178216926, 32'sd-0.10983705719823222, 32'sd-0.11013593839890062, 32'sd-0.06821481266240485, 32'sd-0.07982104529869123, 32'sd0.04344837966372968, 32'sd0.06408996845738087, 32'sd-0.030495141929643005, 32'sd-0.08755583403061074, 32'sd0.10419003953627409, 32'sd0.013712783684704818, 32'sd-0.01898628658906995, 32'sd-0.03876007308528142, 32'sd0.0036758701963675116, 32'sd-0.034074365424652656, 32'sd-0.07697781298274782, 32'sd0.028728320722517586, 32'sd0.09165609950064459, 32'sd0.13601831423344168, 32'sd0.14735451803144603, 32'sd0.18385791232147383, 32'sd0.08494839236767318, 32'sd0.08487354175836115, 32'sd-0.060508848340975745, 32'sd-0.04373041567959722, 32'sd-0.04254978548023207, 32'sd-0.01820931278951901, 32'sd-0.0910937127217187, 32'sd-0.02879233157787, 32'sd-0.04734843950645033, 32'sd-0.13387238175706628, 32'sd0.014391703917764412, 32'sd-0.02634394132955782, 32'sd0.007808918268121684, 32'sd2.030829008018263e-123, 32'sd0.007833688807670592, 32'sd-0.0739413219388955, 32'sd0.07039007778643909, 32'sd0.020543477271714232, 32'sd-0.08154872193103359, 32'sd-0.12141075016233989, 32'sd-0.0334286460719983, 32'sd-0.01601007999019564, 32'sd-0.037937006032365946, 32'sd-0.036829190749563354, 32'sd0.10323428909782832, 32'sd0.09268815503726432, 32'sd0.017487723768319564, 32'sd0.22224231491188065, 32'sd0.10373257117498431, 32'sd0.1764541676879662, 32'sd-0.0020026305831247104, 32'sd0.011800404381767536, 32'sd-0.04050743459196017, 32'sd-0.08756199245540781, 32'sd-0.13137448202009508, 32'sd-0.16347405304138646, 32'sd-0.08207463631048001, 32'sd0.031136590088131914, 32'sd0.07757998112597453, 32'sd-0.05606634549713415, 32'sd-0.015110904255446764, 32'sd0.09839110634216347, 32'sd0.026576911070237928, 32'sd0.04806821166044609, 32'sd0.05925825966366282, 32'sd0.03450644228074248, 32'sd-0.06279895696776325, 32'sd-0.1406936759384931, 32'sd-0.1150207982388785, 32'sd-0.12267917455286131, 32'sd-0.02793570149019538, 32'sd-0.04707721392843873, 32'sd-0.05448294010687928, 32'sd-0.07411657462819231, 32'sd0.07968710890990609, 32'sd0.07850343290307188, 32'sd-0.021981618922610892, 32'sd-0.003963717084979327, 32'sd0.009461720170517137, 32'sd0.10140345432972227, 32'sd0.06616859836642885, 32'sd-0.05942351801832728, 32'sd-0.0682605229223762, 32'sd0.02676801367077611, 32'sd0.05668187155289974, 32'sd0.03330735887513346, 32'sd0.0852693507999954, 32'sd-0.09619004494658012, 32'sd-0.05111027899968988, 32'sd0.102786051869671, 32'sd0.09107086495509038, 32'sd0.017547310697067022, 32'sd-0.0366846031429478, 32'sd0.030734898637527017, 32'sd0.024534724709179476, 32'sd-0.04814318667385447, 32'sd-0.07003995453846486, 32'sd-0.12366126661289827, 32'sd-0.06573734113637252, 32'sd-0.0021715155219685068, 32'sd0.022247905951832608, 32'sd-0.07791818682480321, 32'sd0.09959808699164194, 32'sd0.10550364198727573, 32'sd-0.05902328973468661, 32'sd0.002241144725823848, 32'sd-0.016577770042868804, 32'sd0.15338132105989077, 32'sd0.13722681714300497, 32'sd0.1131374692543473, 32'sd0.14403650545573482, 32'sd0.06100635397961681, 32'sd-0.020351672622879537, 32'sd-0.08893896289393703, 32'sd-0.027171425866086018, 32'sd0.039886472432128735, 32'sd0.06035561581790192, 32'sd1.1063351205608225e-121, 32'sd0.07505739574847409, 32'sd0.032387994615133114, 32'sd0.023661184789966025, 32'sd-0.017627709236912585, 32'sd-0.09178578683615182, 32'sd-0.07362577091135335, 32'sd-0.057557524064184504, 32'sd-0.0697536930284773, 32'sd-0.031258231300310496, 32'sd0.035059273447823884, 32'sd-0.05382942031173637, 32'sd0.11611460374382332, 32'sd0.11886169963765905, 32'sd0.14933545431544487, 32'sd-0.07356381244946683, 32'sd0.07532079640503396, 32'sd0.02699376556439823, 32'sd0.1361999840778524, 32'sd0.005043253535540088, 32'sd0.09468390208337987, 32'sd0.08595871978814562, 32'sd0.053848196929429326, 32'sd-0.09625893553586863, 32'sd-0.07993034833712857, 32'sd0.04816924006911217, 32'sd0.026814665437907267, 32'sd-7.480516394455098e-122, 32'sd-3.416487666150987e-114, 32'sd3.106925582375998e-124, 32'sd-0.06869022223762203, 32'sd-0.05077200690779725, 32'sd-0.08711629499934796, 32'sd-0.021105921902002642, 32'sd-0.009914107972720122, 32'sd0.09295432094384692, 32'sd0.048031836098441506, 32'sd-0.0518683755167245, 32'sd-0.011140161189453561, 32'sd-0.07009956201897914, 32'sd0.041887352011544705, 32'sd0.018726328138214517, 32'sd0.09523858409997002, 32'sd0.09029356608543292, 32'sd-0.060418982013772236, 32'sd-0.08479194572032359, 32'sd0.05718944492729132, 32'sd0.03223042924143643, 32'sd0.08828482847877188, 32'sd-0.023439037692154007, 32'sd-0.07556128184410327, 32'sd-0.058526886637344656, 32'sd-0.004416335608355688, 32'sd0.02515427578036297, 32'sd0.10251898622478943, 32'sd7.577597468231644e-121, 32'sd1.3405677212590374e-122, 32'sd-1.0607900789682562e-126, 32'sd0.06305567270737401, 32'sd0.06484113637835649, 32'sd-0.03612950377278483, 32'sd0.026962105166439532, 32'sd-0.08046349716277051, 32'sd0.000878962325114912, 32'sd0.008980959322866309, 32'sd0.03363045221272634, 32'sd-0.11273444460200616, 32'sd-0.00604589089989944, 32'sd0.10847300951149753, 32'sd0.07644879012856007, 32'sd0.09536653875842735, 32'sd0.046462882602993597, 32'sd0.01079184351365887, 32'sd-0.07802058839166472, 32'sd-0.06851351108469991, 32'sd0.0004487432259842102, 32'sd0.024077465303178225, 32'sd0.06661638043844519, 32'sd0.023528572990066932, 32'sd0.01628548044472779, 32'sd0.009987324776258556, 32'sd0.062100780808031754, 32'sd-0.05303971802803926, 32'sd-4.18192624451208e-125, 32'sd-8.632572886154118e-117, 32'sd9.268289116889334e-125, 32'sd8.369954688679039e-127, 32'sd0.08340252064168988, 32'sd0.053378361520316005, 32'sd-0.006774767057645374, 32'sd0.015519255676583575, 32'sd-0.06784535381608346, 32'sd-0.05911687269106096, 32'sd-0.09273984307385535, 32'sd0.033464511644656386, 32'sd0.004112085040180901, 32'sd-0.08172734196041156, 32'sd-0.14503673852573862, 32'sd-0.0029699116011401685, 32'sd-0.07297047000638177, 32'sd0.02285876791666702, 32'sd0.027170345175693392, 32'sd0.08759218163890593, 32'sd0.08427996355160114, 32'sd-0.08407912923086722, 32'sd-0.08895941981261166, 32'sd-0.13004851068338136, 32'sd0.0677399238110818, 32'sd0.04203522532640329, 32'sd0.04202259892383454, 32'sd-2.165178732869224e-126, 32'sd-4.834199442255641e-123, 32'sd3.920240786951624e-125, 32'sd-8.549729687527739e-122, 32'sd-2.429129592447266e-119, 32'sd-6.520370531668294e-120, 32'sd0.06721554806744295, 32'sd0.02118307496890751, 32'sd0.05329255562242501, 32'sd-0.008413265515687997, 32'sd-0.0602369507266147, 32'sd-0.005417511152642004, 32'sd-0.0024072310025583864, 32'sd-0.03589403041279058, 32'sd0.01912833963397459, 32'sd-0.027891825728919913, 32'sd-0.06018382929514521, 32'sd0.050787627032432794, 32'sd-0.06168438289132207, 32'sd0.02438751518268992, 32'sd0.02772366578736964, 32'sd0.003838131373113568, 32'sd-0.07964418881463711, 32'sd0.06671356951337111, 32'sd0.05116690165114504, 32'sd0.001714686617496533, 32'sd-7.10530863469679e-122, 32'sd-3.209266763135981e-120, 32'sd-1.4944397001463442e-123, 32'sd2.9799607273254478e-117},
        '{32'sd-4.286752715092232e-123, 32'sd-4.241469699168677e-115, 32'sd5.8883508278024235e-115, 32'sd3.356611322885337e-126, 32'sd-1.1928743967076328e-118, 32'sd-1.0821138356259666e-121, 32'sd6.934831678822231e-123, 32'sd-8.903820905952488e-127, 32'sd1.951266232176744e-121, 32'sd2.8620951667008615e-118, 32'sd-3.29681752591981e-115, 32'sd-2.344130316165502e-116, 32'sd0.07744880293750578, 32'sd0.08124922354081181, 32'sd0.043516426240193855, 32'sd0.0551564877220129, 32'sd2.199250840559445e-114, 32'sd1.3554357576120832e-118, 32'sd-7.583461399093367e-124, 32'sd-1.676690014740306e-126, 32'sd1.5740971976138023e-116, 32'sd5.601114066804496e-117, 32'sd9.633405164717598e-121, 32'sd-2.1707076934632123e-127, 32'sd5.551844633376518e-124, 32'sd1.357389423128701e-121, 32'sd3.313936987505172e-122, 32'sd-8.843761595915278e-121, 32'sd-9.782720134338609e-116, 32'sd-4.18560271119056e-121, 32'sd4.087340367424132e-126, 32'sd-3.1571067950631665e-127, 32'sd0.10039507188186636, 32'sd-0.07633467923446935, 32'sd0.037437181153045555, 32'sd0.05242596526099427, 32'sd0.0328105791892893, 32'sd-0.004066356869423754, 32'sd0.000723339768767097, 32'sd0.048264284923181515, 32'sd0.034817839318279475, 32'sd0.021797183297168683, 32'sd0.04879266687303573, 32'sd-0.054400628034307244, 32'sd0.06683771025579749, 32'sd0.03155051525185686, 32'sd0.11870810277271285, 32'sd0.009005371772182606, 32'sd-0.03155521990696499, 32'sd0.004863223703355511, 32'sd0.006148688765917705, 32'sd0.06567642487898756, 32'sd1.646824190263862e-116, 32'sd-6.856743262376417e-119, 32'sd9.471508587137424e-120, 32'sd-3.048447990522087e-116, 32'sd-2.495660097173357e-118, 32'sd-6.796607381463793e-121, 32'sd0.035192509532417635, 32'sd0.027899410922637688, 32'sd0.044957091007555364, 32'sd0.0425110087113891, 32'sd0.051368835457619715, 32'sd-0.08908389258996798, 32'sd0.025941854570840157, 32'sd0.0162080549234635, 32'sd0.04964913856004257, 32'sd0.034831729252457595, 32'sd-0.0650226490539067, 32'sd-0.022578029940412678, 32'sd0.034396225933051444, 32'sd-0.11139150762660915, 32'sd-0.17643554688290572, 32'sd-0.04008226662120368, 32'sd-0.026954418768475315, 32'sd0.0046079984603097915, 32'sd0.007146967187566037, 32'sd0.09389287589812226, 32'sd0.05039997580518808, 32'sd-0.08694681369562289, 32'sd0.0632346211311668, 32'sd0.04582741685456745, 32'sd-1.630245137372166e-123, 32'sd3.0087620633667426e-117, 32'sd7.535768845261557e-115, 32'sd5.585846281648499e-126, 32'sd-0.0035077305080552495, 32'sd0.024179975515736432, 32'sd0.03609331736960999, 32'sd0.04095236530769636, 32'sd0.10423109664840928, 32'sd0.03509539393406377, 32'sd-0.06836481019110217, 32'sd-0.0031720340597737964, 32'sd-0.03706574577859072, 32'sd-0.05985666295773777, 32'sd-0.114327659883724, 32'sd-0.17610557505749228, 32'sd-0.06337620115096272, 32'sd-0.10345223011671381, 32'sd-0.09398640878911818, 32'sd-0.06837380055854742, 32'sd-0.21237069619851368, 32'sd-0.05185203929522429, 32'sd-0.1281043907667175, 32'sd-0.09213639034201457, 32'sd-0.020245153117097722, 32'sd0.016756775572112786, 32'sd0.0827443844841379, 32'sd0.006854917785236206, 32'sd-0.04604301690508277, 32'sd1.5742543784947992e-123, 32'sd-9.260088559781603e-122, 32'sd0.06462971967160797, 32'sd0.032297313179158293, 32'sd-0.022873022460073257, 32'sd0.021077292696353885, 32'sd0.031246167507482634, 32'sd-0.0067037054505071, 32'sd0.06688614380466511, 32'sd0.1504698911179327, 32'sd0.043194085365631955, 32'sd0.01835383316061811, 32'sd-0.07602646419642817, 32'sd-0.00803553221946248, 32'sd0.06146335331259921, 32'sd-0.12577870673748517, 32'sd-0.16075041093505046, 32'sd-0.1806825464114675, 32'sd-0.059535718106050114, 32'sd-0.07726392556948722, 32'sd-0.07204448283258848, 32'sd-0.004073983833617229, 32'sd-0.0028358567175405885, 32'sd0.11956328771660373, 32'sd0.09115428155782375, 32'sd-0.05785977921055858, 32'sd-0.011582415188135086, 32'sd-0.029198462483400182, 32'sd0.10097449499883746, 32'sd-1.613611657067355e-115, 32'sd0.040141376571397006, 32'sd0.12513357909890893, 32'sd0.028540378212703568, 32'sd0.03178142776407159, 32'sd0.11929099912254192, 32'sd0.10197585136853064, 32'sd0.037450845814818015, 32'sd0.11307185959715134, 32'sd0.10878723589481958, 32'sd0.05073687216930213, 32'sd-0.056100211711622994, 32'sd-0.14857635649514114, 32'sd-0.19481652810397787, 32'sd-0.13399943920888494, 32'sd-0.08713018300537885, 32'sd-0.04724835480229851, 32'sd-0.015301753793195275, 32'sd-0.07707302287216794, 32'sd-0.08398162643739912, 32'sd-0.08701793462131271, 32'sd0.01082181887943558, 32'sd0.07042988973637324, 32'sd0.11621858226844446, 32'sd-0.03290688814676262, 32'sd-0.008571040201150931, 32'sd-0.011776940200256757, 32'sd-0.0013683413040753594, 32'sd1.0874138882239174e-121, 32'sd-0.023160794759271627, 32'sd-0.03895239685312945, 32'sd-0.0019849920196296, 32'sd0.05905857619132217, 32'sd0.003024678233582261, 32'sd-0.12500304950828028, 32'sd-0.001203221030463828, 32'sd0.08027820310681338, 32'sd0.05177392777069203, 32'sd0.005741882493691574, 32'sd-0.08498938009035754, 32'sd-0.06701986957980798, 32'sd-0.20834376650898498, 32'sd-0.19471643930003116, 32'sd-0.17496808297463953, 32'sd-0.1305143354994106, 32'sd-0.11496213757171553, 32'sd-0.06275844747245884, 32'sd-0.013672720082276355, 32'sd0.013768281758338895, 32'sd-0.09308138125364387, 32'sd-0.13175169059429906, 32'sd-0.062185984869990954, 32'sd-0.04837020910068837, 32'sd-0.07727736826398289, 32'sd0.10459253402332529, 32'sd0.019525856728241423, 32'sd0.03455520405303354, 32'sd0.04531034661798795, 32'sd-0.06440239547978643, 32'sd-0.14207229266166538, 32'sd-0.010889252858652661, 32'sd0.034229702504772815, 32'sd-0.1307756458299639, 32'sd0.07487276252839468, 32'sd0.08005232425715364, 32'sd0.16131411560981612, 32'sd-0.014142403555690707, 32'sd-0.03158851866956722, 32'sd-0.06803625961357508, 32'sd-0.21950868489393932, 32'sd-0.259895909581859, 32'sd-0.17637049085727471, 32'sd0.00047886217996710365, 32'sd-0.07902290181253858, 32'sd-0.1413274443130272, 32'sd-0.11340029743355969, 32'sd0.0391457759497889, 32'sd-0.1259103863225742, 32'sd-0.07518973813766079, 32'sd-0.12137050413726129, 32'sd0.048637089978537544, 32'sd-0.005926769761806992, 32'sd-0.014060413423306096, 32'sd-0.05930158413199589, 32'sd0.046598501887431185, 32'sd-0.006200774732537787, 32'sd-0.04001580198251091, 32'sd-0.05798325321585621, 32'sd0.12955822399683642, 32'sd0.0259664251306739, 32'sd-0.007154611262806697, 32'sd0.0854206561416223, 32'sd3.565511325710821e-05, 32'sd0.10178592066213243, 32'sd0.05638370110915916, 32'sd0.051555891857465466, 32'sd-0.11694464056743398, 32'sd-0.1992470276351128, 32'sd-0.17908084720099285, 32'sd-0.10378389001735729, 32'sd-0.0069528841630976945, 32'sd0.004642639540025635, 32'sd-0.04088473813930888, 32'sd-0.04383659355421763, 32'sd-0.02347465205913887, 32'sd-0.10054199020801795, 32'sd-0.02824753867129127, 32'sd-0.02267470246547592, 32'sd0.1065094931871349, 32'sd-0.009512631410004399, 32'sd0.017863546814621684, 32'sd-0.08973692868733864, 32'sd0.07242738565539852, 32'sd0.04851246690292791, 32'sd0.08282352119728396, 32'sd0.031120311136331943, 32'sd0.020584595822776625, 32'sd-0.13267514688357337, 32'sd-0.12953477870166913, 32'sd-0.029433286724039137, 32'sd-0.015061487052991259, 32'sd0.03828576242502854, 32'sd0.09237297643693917, 32'sd0.04091018916805619, 32'sd-0.1615351500787833, 32'sd-0.28453137629886543, 32'sd-0.21605501477200634, 32'sd-0.09685586319251388, 32'sd0.08766045723890951, 32'sd0.10286462871690348, 32'sd0.01054174707612557, 32'sd0.06593204533208427, 32'sd0.020984216397666254, 32'sd0.08896140570637813, 32'sd-0.07181683117435005, 32'sd-0.024045465463770194, 32'sd0.026218966095145815, 32'sd-0.04283708462551971, 32'sd0.0276265263175629, 32'sd0.07429997229488838, 32'sd0.030050325257328443, 32'sd0.04318179214383326, 32'sd0.11807373135318341, 32'sd-0.04111877616486702, 32'sd-0.07358704742286738, 32'sd-0.09077968670334799, 32'sd-0.10351752843241356, 32'sd0.038082415268263024, 32'sd0.05944694702579315, 32'sd0.051457462068223776, 32'sd0.04631612662202638, 32'sd0.0476446201423073, 32'sd-0.16945050691205568, 32'sd-0.18345107279102651, 32'sd-0.1868628130297932, 32'sd0.09418668498586914, 32'sd0.09426744082548201, 32'sd0.06795201442192182, 32'sd0.03107628830424762, 32'sd0.01476335997747252, 32'sd-0.103815215694564, 32'sd0.03550805534181986, 32'sd0.008128198341424153, 32'sd-0.04477013162377805, 32'sd0.16135724434960597, 32'sd0.06924270878488586, 32'sd0.08844742871371138, 32'sd-0.02511007090534445, 32'sd0.03703238310283555, 32'sd0.11179454180573851, 32'sd-0.063548549280047, 32'sd-0.0447087779884121, 32'sd0.003329214171930155, 32'sd0.07044792360600476, 32'sd0.016431792677865757, 32'sd-0.0007319611284334699, 32'sd-0.04326605502960228, 32'sd0.013158674342197037, 32'sd-0.03371207584205551, 32'sd-0.01963732531807743, 32'sd-0.11196844309770744, 32'sd-0.17063364070904777, 32'sd-0.08514165104117441, 32'sd0.09951359474322247, 32'sd-0.02010649416740569, 32'sd-0.07874790322924187, 32'sd-0.009890060291011927, 32'sd0.07533785270334416, 32'sd-0.005915776783476615, 32'sd0.029958312505570104, 32'sd-0.001969954620787522, 32'sd0.03611376318843579, 32'sd0.09167735924842044, 32'sd-0.006660414931150165, 32'sd-0.06791740087096214, 32'sd-0.00023896189308822644, 32'sd0.0864638615843921, 32'sd0.010558938278465824, 32'sd0.0038442791614166586, 32'sd-0.0060240660803824765, 32'sd0.009405671532013877, 32'sd-0.036032533545812276, 32'sd-0.04407339529546153, 32'sd-0.05513319354471508, 32'sd-0.09758609495238764, 32'sd-0.08924023558410085, 32'sd0.03520630537436255, 32'sd-0.04007913504852887, 32'sd-0.008753108602611656, 32'sd0.030800776657468307, 32'sd0.11756069470116357, 32'sd0.12681493598340313, 32'sd0.15952630440367954, 32'sd-0.04635151428638479, 32'sd-0.09883883135646146, 32'sd0.03594846592481643, 32'sd0.11152510920933993, 32'sd0.10157097163230314, 32'sd0.11819022120488736, 32'sd-0.0017883226657076404, 32'sd-0.027791533064181702, 32'sd0.10196745882771055, 32'sd-0.028688354319975427, 32'sd0.009193742811837533, 32'sd0.029291211540189488, 32'sd0.1134091575473941, 32'sd-0.04937252260051934, 32'sd-0.02784467034702626, 32'sd-0.010820929282081178, 32'sd0.03421535611960207, 32'sd-0.08064949771977391, 32'sd0.03144767415754671, 32'sd0.05347335200400956, 32'sd-0.025695630525446052, 32'sd0.07488605413664959, 32'sd-0.004210304589179268, 32'sd-0.05557414420489153, 32'sd0.013426697895344938, 32'sd0.09315876626715539, 32'sd0.07981027292279996, 32'sd-0.012622280141822933, 32'sd0.06498444783221159, 32'sd0.05349445259531728, 32'sd0.18397098533598338, 32'sd0.17009646691579494, 32'sd0.15226327804789874, 32'sd0.1515435286821969, 32'sd0.10938178891097582, 32'sd-0.005665995289626283, 32'sd-0.018447482489306468, 32'sd0.035300913501678396, 32'sd-0.07860006675361837, 32'sd0.025826362186285735, 32'sd0.013559161987479213, 32'sd0.011562567870883196, 32'sd-0.10564629869962638, 32'sd0.10577773568062825, 32'sd0.1529878776305517, 32'sd0.067676947062601, 32'sd0.14864015211836604, 32'sd0.07075422087263751, 32'sd0.09381672182610747, 32'sd0.04752457159515539, 32'sd0.002350374126711942, 32'sd0.1940217556335664, 32'sd0.16311882477016948, 32'sd0.06264715814778112, 32'sd-0.009685296183935514, 32'sd0.05238902973139906, 32'sd0.08544221047922626, 32'sd-0.020841357664002275, 32'sd0.16644027560574803, 32'sd-0.0005794171419693991, 32'sd0.04494598403275787, 32'sd0.07086212825424802, 32'sd0.05072914858105002, 32'sd0.11948847993966188, 32'sd0.05499639733954572, 32'sd-0.05675608328631058, 32'sd0.04718886251170686, 32'sd-0.022247182559063106, 32'sd-0.015563386034993243, 32'sd0.022066312162120173, 32'sd0.05891259345614389, 32'sd-0.038079484051655725, 32'sd0.06605957339426032, 32'sd0.04790476803653087, 32'sd0.1751193961364624, 32'sd0.11424787251909, 32'sd0.06449238573766511, 32'sd0.16928007822839888, 32'sd0.11122634435017831, 32'sd0.1192794525791358, 32'sd0.18668047627213208, 32'sd0.15025431267700798, 32'sd0.012812623551236173, 32'sd-0.006759743305179537, 32'sd0.10852049696347588, 32'sd-0.03922687110001565, 32'sd0.036127288464144265, 32'sd0.050525528727836166, 32'sd-0.07870254125453273, 32'sd0.0932210803563904, 32'sd-0.00046805294962376927, 32'sd0.03170426391991948, 32'sd0.0979624330736931, 32'sd-0.04865611029454305, 32'sd0.06984466696208308, 32'sd0.027038649262634842, 32'sd0.11607362204923799, 32'sd-0.037562209413664734, 32'sd0.009808312283252825, 32'sd-0.08031514412610871, 32'sd0.05367227439473612, 32'sd0.07902088143737797, 32'sd0.10095754326851547, 32'sd0.05603857814233978, 32'sd-0.019007812033461274, 32'sd0.008118640612558937, 32'sd0.011009966061999757, 32'sd0.07630984673996721, 32'sd-0.037035264502246625, 32'sd-0.03692582590776942, 32'sd0.20340930771385518, 32'sd0.018719325163498807, 32'sd0.053352648545083724, 32'sd0.11098019645185357, 32'sd0.07202525028993112, 32'sd0.10036068064029975, 32'sd0.025722205505366375, 32'sd-0.040917632139420484, 32'sd-0.061776537472058635, 32'sd-0.1781343682842537, 32'sd-0.06006258154057339, 32'sd-0.06652643316926163, 32'sd0.04157199042742492, 32'sd4.103704027121591e-121, 32'sd0.029618781800326746, 32'sd-0.047186965095612994, 32'sd-0.024566021042593558, 32'sd-0.037766222784848216, 32'sd0.09528428658345744, 32'sd0.03404343476470664, 32'sd0.014465922497135625, 32'sd0.059879254311258144, 32'sd-0.010279547770606821, 32'sd0.07699184821548052, 32'sd-0.016495499326863484, 32'sd0.006566434755657947, 32'sd0.005122837525810473, 32'sd0.07984505002226994, 32'sd0.07681306423741832, 32'sd-0.002106308648819039, 32'sd-0.013004423293547627, 32'sd-0.005465764493918457, 32'sd0.02417694751716284, 32'sd0.10591550922402264, 32'sd0.05431591296363535, 32'sd-0.012295255176114869, 32'sd-0.023709269440392616, 32'sd-0.13164478790375994, 32'sd-0.03760910427002806, 32'sd-0.014255601076133408, 32'sd-0.05326291447617027, 32'sd0.007181473850342237, 32'sd0.05155131046604408, 32'sd-0.05674457162425011, 32'sd0.05037643672784893, 32'sd0.0015134350771033316, 32'sd-0.004804109728264389, 32'sd0.08196673938080175, 32'sd-0.06765987979287189, 32'sd-0.03854932764369421, 32'sd0.07142676891063314, 32'sd0.038952042255020004, 32'sd0.12520916155559686, 32'sd0.028033750139352075, 32'sd0.01138094179960613, 32'sd0.14444715145191886, 32'sd0.04805488020990757, 32'sd-0.0061220563822216075, 32'sd0.031202137954938654, 32'sd0.09504529487067763, 32'sd0.08877597870731607, 32'sd0.1356897996999753, 32'sd0.05611904947661599, 32'sd-0.033233709723338466, 32'sd-0.10334676910485598, 32'sd-0.0523735802154817, 32'sd0.021756840435472775, 32'sd0.020907059220694937, 32'sd0.09057888415864913, 32'sd0.02725377887305315, 32'sd0.03587041502050211, 32'sd0.031932240205273243, 32'sd0.07760017158928724, 32'sd0.07616924352175836, 32'sd0.07888591840977292, 32'sd0.10718361637711495, 32'sd0.07819261602311459, 32'sd0.05253214484574716, 32'sd0.03983468870402865, 32'sd0.06279091632955157, 32'sd-0.001304547876225797, 32'sd-0.14014882786286617, 32'sd-0.08204654561192405, 32'sd-0.048466014269919686, 32'sd0.024548753156629476, 32'sd0.05466447597662494, 32'sd-0.05506974750562935, 32'sd0.04977519150197175, 32'sd-0.10704070845628352, 32'sd-0.00396314108449744, 32'sd0.05190477599452428, 32'sd-0.026172088894083838, 32'sd-0.0005973837180751734, 32'sd-0.11473347178729401, 32'sd-0.0928809371824912, 32'sd-0.06139976806571934, 32'sd0.02814618510504762, 32'sd-7.671405576010666e-125, 32'sd0.03091808273843216, 32'sd-0.022390754583129457, 32'sd0.05378130540051167, 32'sd0.07488247334645674, 32'sd0.02513227310498664, 32'sd0.14956912338873476, 32'sd0.07276703546400272, 32'sd-0.036218979692355525, 32'sd0.0078854626333737, 32'sd-0.1256532780699483, 32'sd-0.023609151200352525, 32'sd-0.20106239499352038, 32'sd-0.1940306693346716, 32'sd-0.02760022277886319, 32'sd-0.027622681876760976, 32'sd0.05923548984220343, 32'sd-0.10890947829615136, 32'sd-0.04239771131680675, 32'sd-0.186452355110212, 32'sd-0.08749999407429289, 32'sd-0.014403802080627732, 32'sd-0.02174297757119505, 32'sd-0.07420823125738854, 32'sd-0.07381183397785035, 32'sd-0.17157809024566137, 32'sd0.02369805522636162, 32'sd0.022028896501178487, 32'sd0.08417409588343994, 32'sd0.0894099296369742, 32'sd0.00959061674651013, 32'sd0.003119594866157705, 32'sd0.08765939245730989, 32'sd0.069583804158887, 32'sd-0.037125424492843236, 32'sd-0.025731736773686148, 32'sd-0.03920987538139654, 32'sd-0.049325923443141934, 32'sd-0.08926862736030863, 32'sd-0.18141559927307277, 32'sd-0.11821576371431614, 32'sd-0.1410652001576946, 32'sd-0.054750917553704134, 32'sd-0.06062518569503312, 32'sd-0.018729132111240124, 32'sd-0.0860628182912393, 32'sd-0.13695253051838555, 32'sd0.006254080094807587, 32'sd-0.05219372176199899, 32'sd0.024736971501802544, 32'sd0.043749066638612645, 32'sd0.0010790723797160621, 32'sd-0.05420495437215255, 32'sd0.05092452914140126, 32'sd0.08342456247315998, 32'sd0.02720444471572151, 32'sd0.07450681125961653, 32'sd0.14892231277847992, 32'sd0.05877728125846062, 32'sd0.07591946956344262, 32'sd-0.03003295452629907, 32'sd-0.01921101068346582, 32'sd-0.07380994051166102, 32'sd0.08448127374534967, 32'sd0.034047055503022415, 32'sd-0.011517825415043011, 32'sd-0.07029994844522285, 32'sd-0.042995331077955744, 32'sd-0.10478298882893246, 32'sd-0.00044700372229508666, 32'sd-0.14588184235893717, 32'sd-0.11806480821138328, 32'sd-0.0631400705899451, 32'sd-0.03932516266607539, 32'sd-0.08068986015227543, 32'sd-0.03784242875836799, 32'sd-0.024535431766114345, 32'sd-0.022772081994207723, 32'sd0.08792908409647725, 32'sd-0.008126006350405683, 32'sd0.09917690952900288, 32'sd-0.05663533055859015, 32'sd-0.009598109616274296, 32'sd0.006789275727964241, 32'sd1.046887212859952e-120, 32'sd0.03757387553570777, 32'sd0.07002076430052102, 32'sd0.03161350344933165, 32'sd-0.016954034261699252, 32'sd0.008207843849825999, 32'sd-0.018063461768193657, 32'sd0.08309509683128438, 32'sd0.0003990814029698824, 32'sd-0.0474194924981266, 32'sd-0.040221936776403025, 32'sd-0.06851547191058834, 32'sd0.005994467841538067, 32'sd-0.0541466101957808, 32'sd-0.07678751443894746, 32'sd-0.07496832063061383, 32'sd-0.010481028049097892, 32'sd0.00457540592207297, 32'sd-0.07086257010156594, 32'sd-0.057792576200704174, 32'sd-0.12228749498438597, 32'sd0.026359158847277284, 32'sd-0.014107490097422364, 32'sd-0.04907562467642296, 32'sd-0.07698151805485139, 32'sd-0.15524178795992888, 32'sd-0.049722628676995874, 32'sd-1.2162054752879677e-124, 32'sd7.598629389723853e-122, 32'sd-3.5282889909357644e-127, 32'sd-0.06842823180375289, 32'sd-0.029964060168978252, 32'sd-0.02903106971075665, 32'sd-0.00040881829821032387, 32'sd-0.07743251878038583, 32'sd-0.040507281701968094, 32'sd-0.015555591577037405, 32'sd-0.008254045747727753, 32'sd-0.0900517090435014, 32'sd-0.10484685584187291, 32'sd-0.03726322633094393, 32'sd-0.04303789702565847, 32'sd0.02125545525464858, 32'sd-0.0885385781841125, 32'sd-0.03662866589658926, 32'sd0.014983537819147744, 32'sd-0.030515684363020924, 32'sd-0.0906860566206437, 32'sd-0.06930507167205083, 32'sd-0.0966720936694007, 32'sd-0.03986828668207338, 32'sd0.06890391917833649, 32'sd0.027895050411219056, 32'sd0.010350312414829576, 32'sd0.09652252521640564, 32'sd1.70064340601612e-123, 32'sd-1.18126236750769e-128, 32'sd1.3410884954835864e-122, 32'sd0.009052938593035041, 32'sd0.003964706402954109, 32'sd-0.0669993686011989, 32'sd-0.08334951748080378, 32'sd0.03442345018810349, 32'sd-0.12443702628765581, 32'sd-0.004793154939946944, 32'sd-0.05041094771072188, 32'sd-0.09932848684584679, 32'sd0.03078013193867639, 32'sd0.04125471188714634, 32'sd-0.052876476456181626, 32'sd-0.07029474766349852, 32'sd0.060951657783241533, 32'sd-0.015666214187065867, 32'sd-0.024805810440972773, 32'sd-0.032017270952266266, 32'sd0.022005313675829925, 32'sd0.07349840054210763, 32'sd-0.09300937738112974, 32'sd-0.11459389210106101, 32'sd-0.009080642863348606, 32'sd0.01973764849249092, 32'sd0.07240383237272469, 32'sd0.037235548196983735, 32'sd-3.389206290506163e-120, 32'sd1.554671947718119e-120, 32'sd-4.2173540485609715e-125, 32'sd2.4729072995002547e-119, 32'sd0.10189536954359191, 32'sd0.00562994389790382, 32'sd-0.01776895634523558, 32'sd-0.13508645899544824, 32'sd-0.0496568266982428, 32'sd-0.11871442054209695, 32'sd-0.1125679460158748, 32'sd-0.154228097544314, 32'sd-0.09518659999502162, 32'sd-0.1749954875942171, 32'sd-0.17361634767156794, 32'sd-0.030548663187540515, 32'sd-0.11128847016027495, 32'sd-0.16286585019860683, 32'sd-0.07165617688269474, 32'sd-0.04111489138825797, 32'sd0.054827682145881435, 32'sd0.03435584038640538, 32'sd-0.11994543438400553, 32'sd-0.02085985688028347, 32'sd-0.1077406664168198, 32'sd0.03633120257209454, 32'sd0.08031800987917023, 32'sd-2.407921931620743e-116, 32'sd-6.234255409243419e-121, 32'sd2.093409820941179e-117, 32'sd2.8248108805466853e-122, 32'sd-5.981365328197572e-119, 32'sd3.480472837697327e-122, 32'sd0.05181486945146587, 32'sd0.018089728567696507, 32'sd0.047464707014424394, 32'sd0.029590924180004658, 32'sd0.04923566545769165, 32'sd-0.0685409370786091, 32'sd-0.0698597993724197, 32'sd-0.08359638580491428, 32'sd0.003961197529204327, 32'sd-0.11519441483961981, 32'sd-0.01436297520440813, 32'sd-0.05022252161809395, 32'sd-0.010376084833652684, 32'sd-0.032398818845765086, 32'sd0.03947893194239731, 32'sd0.04140963991270229, 32'sd0.06044263963340006, 32'sd0.0326037928336899, 32'sd-0.016980104723289792, 32'sd0.0031012876357081752, 32'sd-1.8034909245832905e-117, 32'sd-6.621347357342172e-121, 32'sd-4.2897529255721296e-126, 32'sd2.9978626645087005e-122},
        '{32'sd-3.1804873170708634e-114, 32'sd2.2405272007364397e-125, 32'sd2.5515468083133454e-124, 32'sd8.125184212801267e-122, 32'sd-2.241439296491641e-122, 32'sd-2.6157992969167356e-120, 32'sd-3.5399511305591215e-116, 32'sd5.624398590687645e-121, 32'sd-1.551559539557525e-125, 32'sd-3.957477813123101e-119, 32'sd1.0650940843606647e-118, 32'sd-9.805562910419157e-119, 32'sd0.008223019546494128, 32'sd-0.07533946159184998, 32'sd-0.033774958237443024, 32'sd-0.06449497430238953, 32'sd3.6762213725986333e-122, 32'sd-2.8737839476526088e-117, 32'sd-1.120259287791777e-125, 32'sd-2.0992101998592497e-118, 32'sd-1.0776507456003186e-124, 32'sd-1.529432730976883e-123, 32'sd1.8386663040478484e-116, 32'sd-3.5885106743651857e-129, 32'sd-1.7185992045765045e-116, 32'sd2.7312440909636517e-127, 32'sd-1.0116640082684257e-121, 32'sd4.009051074203197e-125, 32'sd2.0252105058485418e-122, 32'sd6.524785456027559e-122, 32'sd-1.4398481976001457e-125, 32'sd-3.241828560134513e-122, 32'sd-0.056961811616581974, 32'sd-0.055026155435547695, 32'sd-0.033063436797184, 32'sd0.0029019329715796248, 32'sd0.026515145182914864, 32'sd-0.040582930939350476, 32'sd0.04651385716380158, 32'sd0.029432727262780532, 32'sd-0.016697954034833918, 32'sd0.029648131349333258, 32'sd-0.0465566908912386, 32'sd-0.05702669734046427, 32'sd-0.091793929116402, 32'sd-0.04764022531570441, 32'sd-0.11405304999514883, 32'sd-0.012535989962413821, 32'sd-0.005951124064204391, 32'sd-0.0011866816640293733, 32'sd0.008656454168778974, 32'sd-0.05142897760215898, 32'sd1.1304420643134237e-124, 32'sd2.2723755742387235e-121, 32'sd-1.6005573859057763e-127, 32'sd-4.952845194768802e-124, 32'sd-8.904216983960219e-127, 32'sd1.0607042550342694e-124, 32'sd0.005421587215688785, 32'sd-0.06357952530559965, 32'sd-0.07986525893386974, 32'sd-0.059534550809819835, 32'sd-0.045488450569039475, 32'sd0.0827503293073234, 32'sd-0.0421489299432393, 32'sd-0.01235228282823357, 32'sd0.004790864978332621, 32'sd-0.08046375259226328, 32'sd-0.023131505203176955, 32'sd-0.06819329666746515, 32'sd0.03104518054520759, 32'sd-0.0872820514600363, 32'sd-0.08882421988052405, 32'sd0.011992446918156149, 32'sd0.01873490602991518, 32'sd-0.06707628049735576, 32'sd-0.12936081459290563, 32'sd-0.07009367238019255, 32'sd-0.09265030846179151, 32'sd-0.017430604630517665, 32'sd0.0578832880607133, 32'sd-0.012156543584445147, 32'sd3.171071144036578e-116, 32'sd8.71903989805905e-126, 32'sd4.015909761867547e-126, 32'sd7.509830901823924e-121, 32'sd-0.07660609127989168, 32'sd-0.06836965227690278, 32'sd-0.026018919822436037, 32'sd-0.01054389769649978, 32'sd0.039045511716906664, 32'sd0.01887180476421972, 32'sd-0.011248358327618415, 32'sd-0.008218717492057038, 32'sd0.04195135968297575, 32'sd-0.1277822646732438, 32'sd-0.07386610151655781, 32'sd-0.15239453406626693, 32'sd-0.03037900465544309, 32'sd-0.09746030122481122, 32'sd0.04301446852779109, 32'sd-0.03852126607796774, 32'sd0.09829240790337151, 32'sd-0.05328926573463417, 32'sd-0.011559733277650797, 32'sd0.05698564978626432, 32'sd-0.10617494722991065, 32'sd0.009634721382471184, 32'sd0.025643772470316212, 32'sd-0.06707202685134177, 32'sd-0.05689473567729398, 32'sd-1.614769303659877e-128, 32'sd-1.934134742057496e-118, 32'sd-0.042787735857078124, 32'sd-0.06843492881205178, 32'sd-0.06722811228954119, 32'sd-0.11441079267297655, 32'sd0.08298782469244315, 32'sd0.006522231247931432, 32'sd-0.0013122121796473164, 32'sd-0.07360189110457664, 32'sd-0.14007896874373787, 32'sd-0.17416952099509259, 32'sd-0.1716929510809351, 32'sd-0.009902565594551938, 32'sd0.017442748452740603, 32'sd-0.011500925959074475, 32'sd-0.0224669350455132, 32'sd0.0374510768940217, 32'sd0.16766575119020136, 32'sd0.12229628103870732, 32'sd-0.060267572880648726, 32'sd-0.03565714350619478, 32'sd-0.041684296857529994, 32'sd-0.03987083889403547, 32'sd0.11510006993635308, 32'sd0.025965846757990057, 32'sd0.03864973188317801, 32'sd-0.057534641758677285, 32'sd0.04104497815288337, 32'sd-7.693078986354805e-125, 32'sd-0.06968330245385242, 32'sd-0.059756558938000456, 32'sd-0.11655665756936262, 32'sd-0.11171263832724816, 32'sd0.041448376734535254, 32'sd0.0007785149965338779, 32'sd-0.015282793631782463, 32'sd-0.11850839918731261, 32'sd-0.13036853963120365, 32'sd-0.08630105272340939, 32'sd-0.030814351645677085, 32'sd-0.04446714800932869, 32'sd-0.01691757990834818, 32'sd-0.00056474272188472, 32'sd0.0270884587090005, 32'sd0.029399575084459853, 32'sd0.13464971887798446, 32'sd0.04353861855696829, 32'sd0.10196854017180448, 32'sd-0.05972262642648667, 32'sd-0.10581934489947604, 32'sd-0.13566916139642599, 32'sd-0.15275058155255047, 32'sd-0.03064891254680533, 32'sd0.09621099718112648, 32'sd-0.04689900458402296, 32'sd-0.04224529888857821, 32'sd-1.7951290972845832e-118, 32'sd-0.0322383672341605, 32'sd-0.09938887211254037, 32'sd0.011548857599795419, 32'sd-0.05480076916300981, 32'sd-0.0741717301379026, 32'sd-0.10403735490504143, 32'sd-0.09668953855377002, 32'sd-0.1958006143917137, 32'sd-0.11950856775876036, 32'sd-0.09325238529800847, 32'sd-0.02687736840972247, 32'sd0.02282872467325161, 32'sd0.008515816692057332, 32'sd0.068159375577409, 32'sd0.10053319557391831, 32'sd-0.008609346902441122, 32'sd0.07478443126602007, 32'sd0.11978624463413318, 32'sd0.013530570927793636, 32'sd0.024406860020613933, 32'sd0.06132264521673857, 32'sd0.020618588279856603, 32'sd0.11376885495262375, 32'sd0.14097805556144835, 32'sd-0.004535211018069407, 32'sd0.0463585018773851, 32'sd-0.049230677313510836, 32'sd-0.06827990744976936, 32'sd0.03573020123014676, 32'sd0.033102405121956266, 32'sd-0.02069463657913133, 32'sd0.09258940492201105, 32'sd-0.1426680902104765, 32'sd-0.12347427103842352, 32'sd-0.11970677158523096, 32'sd-0.13856695637305363, 32'sd-0.09608358927627193, 32'sd0.12581515331687612, 32'sd0.1322504091696623, 32'sd0.23264466235120154, 32'sd0.14545657341824306, 32'sd-0.008533762850956405, 32'sd0.07693742497623414, 32'sd0.011657430108875502, 32'sd-0.02717449850212996, 32'sd0.17170618164089205, 32'sd0.05291875880492966, 32'sd-0.07720547626256292, 32'sd-0.06778089113039357, 32'sd-0.03980858202757377, 32'sd-0.0551093798446467, 32'sd0.12419955912631887, 32'sd-0.009406284909445652, 32'sd-0.04759422584087798, 32'sd0.0028061794741707164, 32'sd0.05383190040391361, 32'sd-0.05870463070327407, 32'sd-0.08119401227908968, 32'sd-0.011102177302106922, 32'sd-0.09527948716694123, 32'sd-0.08013365089476328, 32'sd-0.12404693017410744, 32'sd-0.12219660420466655, 32'sd-0.05248188770904332, 32'sd0.018528185215876486, 32'sd0.15384012169053626, 32'sd0.25765488052549823, 32'sd0.175020083667198, 32'sd0.048130374283014914, 32'sd0.07538401908641923, 32'sd-0.027423383727701107, 32'sd0.04125812886017763, 32'sd0.03570777535808606, 32'sd0.046335553509849775, 32'sd0.10493990521025451, 32'sd0.10155058919335118, 32'sd0.028575656500876713, 32'sd0.014962037507815827, 32'sd-0.005451727453468077, 32'sd0.00957560333630556, 32'sd-0.0464536468470322, 32'sd0.0382708898318063, 32'sd0.03154355270969166, 32'sd-0.037052022852533305, 32'sd-0.08266747490801288, 32'sd-0.08229525339121897, 32'sd-0.058206090834159875, 32'sd0.12639707220616278, 32'sd0.060202721470118285, 32'sd-0.10512207420052773, 32'sd-0.03131682532100459, 32'sd0.05360363924176464, 32'sd0.07466188413856156, 32'sd0.07814057111855995, 32'sd0.08043861615189198, 32'sd0.11384422771310747, 32'sd0.12143591543386345, 32'sd-0.020066404378304415, 32'sd0.0059027603344282455, 32'sd-0.026678277612602087, 32'sd0.040112651492067546, 32'sd0.051517866498456376, 32'sd0.05257033766737139, 32'sd0.21763631511574133, 32'sd0.0947488097009443, 32'sd-0.05759473805861015, 32'sd0.06696300230770358, 32'sd0.016761027315719247, 32'sd0.12866227567902608, 32'sd0.010217206194114325, 32'sd-0.04058026050085536, 32'sd-0.09568111098923232, 32'sd0.0008581873631231974, 32'sd0.06274931558401532, 32'sd-0.006514989996567631, 32'sd0.029080195170436064, 32'sd0.0840128138387322, 32'sd0.03652908863740886, 32'sd0.09552494411648199, 32'sd-0.03578198952007949, 32'sd-0.023647863823216052, 32'sd0.02860927442566427, 32'sd0.0853874182366389, 32'sd0.07327483014678086, 32'sd-0.0026539890247634914, 32'sd0.009210945747078984, 32'sd-0.12483060992828869, 32'sd-0.09024733202758874, 32'sd0.05218294419200067, 32'sd0.10762475684979919, 32'sd0.040430597727611886, 32'sd0.05711716729305041, 32'sd0.15076798358658014, 32'sd0.010571063044664554, 32'sd0.0393923237621885, 32'sd0.07514391192080642, 32'sd0.07298954682818418, 32'sd-0.0669713164163342, 32'sd0.018550573370005072, 32'sd-0.07970642784761096, 32'sd0.11596621308084609, 32'sd0.04129295111546809, 32'sd-0.07913037821783624, 32'sd-0.10882991046775602, 32'sd-0.06627225008112123, 32'sd-0.046045291277835375, 32'sd0.09685175463718068, 32'sd-0.09440780313660485, 32'sd-0.02506042652986765, 32'sd0.08137291263102046, 32'sd0.07024001144367857, 32'sd0.17511878050035545, 32'sd0.09809296259212436, 32'sd0.004611519212435279, 32'sd-0.043732809130829366, 32'sd-0.020907084660447727, 32'sd0.10532689990073495, 32'sd0.023197894327693952, 32'sd-0.005332755591614972, 32'sd0.02794364005578511, 32'sd0.011725772765562179, 32'sd0.024934474000757382, 32'sd0.12110151569923037, 32'sd-0.020342523338050485, 32'sd0.026091659986387572, 32'sd0.05099069550460099, 32'sd-0.13030677359964907, 32'sd-0.0466248417535305, 32'sd0.00499822326581275, 32'sd-0.06986693616998536, 32'sd-0.10343343302078876, 32'sd0.005051892918413838, 32'sd-0.06358977888430743, 32'sd0.04699003216924084, 32'sd-0.0826465318753247, 32'sd0.021647402781652628, 32'sd-0.05176876323313483, 32'sd0.02602626228692521, 32'sd0.056463034618102426, 32'sd0.04108664288783139, 32'sd0.04948789538567077, 32'sd-0.005008711869328053, 32'sd-0.17294045349170295, 32'sd-0.004616337659512262, 32'sd0.12406477282271877, 32'sd0.011777403353907409, 32'sd0.08737862090052777, 32'sd0.010282566573721681, 32'sd0.02766047806596068, 32'sd0.10691857743887533, 32'sd-0.022128558917411795, 32'sd0.040648617482031586, 32'sd-0.04875199962258549, 32'sd0.01583928994599264, 32'sd-0.09783343368114297, 32'sd0.04835612362710686, 32'sd-0.051089022397146265, 32'sd0.019907439575627354, 32'sd-0.03442204124187317, 32'sd0.06645246037308666, 32'sd-0.05545268166337905, 32'sd-0.11813421990392295, 32'sd-0.0811101003031755, 32'sd0.005065077875506945, 32'sd0.018670181535104077, 32'sd0.0038465244811298396, 32'sd-0.08094459334723825, 32'sd0.012027143658224396, 32'sd-0.041565208232081374, 32'sd-0.10866331486830216, 32'sd-0.12193863376391305, 32'sd-0.11845304891301588, 32'sd-0.015673615655133224, 32'sd-0.12300157403585932, 32'sd0.03855524331259701, 32'sd-0.03562424003095533, 32'sd0.017483437239252286, 32'sd0.008196777406906695, 32'sd0.09183565206992828, 32'sd0.06292363888199787, 32'sd0.04080568363987872, 32'sd-0.061643661711112165, 32'sd-0.03336286108378528, 32'sd-0.03772072539968945, 32'sd0.005170604195546823, 32'sd0.06938201462143133, 32'sd-0.034311734743000956, 32'sd0.12177534498114694, 32'sd0.07722454850255756, 32'sd-0.06769584420276901, 32'sd-0.12755545819060468, 32'sd-0.17218047229090314, 32'sd-0.16828248467395016, 32'sd0.007441229823005398, 32'sd-0.12743804751470503, 32'sd0.10076078070480407, 32'sd0.022523178615232755, 32'sd0.03800360367960978, 32'sd0.05692739459010377, 32'sd-0.05621029606942325, 32'sd-0.051614732358346245, 32'sd-0.10068465567866204, 32'sd-0.05962087311836989, 32'sd-0.029730447577675012, 32'sd-0.0016254086984891808, 32'sd-0.0004254318954940048, 32'sd0.08460081335550183, 32'sd0.08826512086800664, 32'sd-0.1397677317840875, 32'sd0.009355258547639222, 32'sd-0.007477669850604462, 32'sd-0.019559084099448145, 32'sd-0.03823282733459277, 32'sd0.027987604270384495, 32'sd-0.00551798689885642, 32'sd0.07078098288600233, 32'sd0.024812272600634212, 32'sd-0.19370570503364812, 32'sd-0.1454545184503975, 32'sd-0.0841301622277525, 32'sd0.07855615265988758, 32'sd-0.0032327784200638604, 32'sd-0.13724319713771646, 32'sd-0.004190667670413578, 32'sd0.02810501339313938, 32'sd0.06826098448954748, 32'sd0.087374856056014, 32'sd0.06229228173882003, 32'sd-0.07326977797981915, 32'sd-0.17396682799489865, 32'sd-0.1665295139194582, 32'sd-0.16598350568157835, 32'sd-0.004170617641147711, 32'sd0.14041249575839557, 32'sd0.07885333945536857, 32'sd0.13693846537796353, 32'sd-0.05035207725001152, 32'sd-0.02140823802362066, 32'sd-0.09966763867581885, 32'sd0.04000639622757615, 32'sd-0.07659145173790924, 32'sd0.009285425532663571, 32'sd-0.0044289318553969725, 32'sd0.0487511710698867, 32'sd-0.020934951856955545, 32'sd-0.1132874690729231, 32'sd-0.16756686887063002, 32'sd0.03162071813965054, 32'sd0.06422741240232213, 32'sd0.14308445523907642, 32'sd-0.058509168658377755, 32'sd0.04302875889352042, 32'sd-0.15449764819527936, 32'sd0.035307101595091935, 32'sd-0.03943945162598378, 32'sd-0.13218397945765067, 32'sd-0.051179902101200096, 32'sd-0.2412241291442364, 32'sd-0.17285819631347726, 32'sd-0.1479617853307533, 32'sd-0.017099350166525067, 32'sd0.02192895028644326, 32'sd-0.04567564991604464, 32'sd-0.035103429264168436, 32'sd-0.075234340459549, 32'sd0.021392985680275603, 32'sd-0.05963836940220747, 32'sd-9.559694243403683e-121, 32'sd0.029189338423988107, 32'sd-0.04840946349813315, 32'sd0.09838026095194262, 32'sd0.07121631781977976, 32'sd-0.0682425067396432, 32'sd-0.012515527114893423, 32'sd0.024274348616732746, 32'sd0.002038895735152091, 32'sd0.024384601843428548, 32'sd-0.020526244618481515, 32'sd0.03968389476265922, 32'sd-0.10522494908944957, 32'sd-0.11984569666892665, 32'sd-0.15776341319465004, 32'sd-0.0059707201376806894, 32'sd-0.16299145361475056, 32'sd0.00797807900928526, 32'sd-0.027227508435809938, 32'sd-0.1326939142959995, 32'sd-0.10523756085870642, 32'sd0.05004005053333737, 32'sd-0.026927198402583237, 32'sd-0.03833351268066062, 32'sd0.07627938953974946, 32'sd0.0520413688535965, 32'sd-0.0032642954201552955, 32'sd-0.06301467718981829, 32'sd-0.06569698310854925, 32'sd-0.0683453808827452, 32'sd0.06332447276059683, 32'sd-0.03916546982597137, 32'sd-0.06030664369979934, 32'sd0.010210664315375935, 32'sd-0.0865332471019796, 32'sd-0.031363756854941076, 32'sd-0.003217120336012605, 32'sd0.02204086461317065, 32'sd0.05126014178894796, 32'sd-0.04218043456203954, 32'sd-0.11659481492508365, 32'sd-0.10936483001789689, 32'sd-0.06087285855953302, 32'sd0.001107072991797601, 32'sd-0.015712694838889332, 32'sd-0.002202289637411828, 32'sd0.0708539499468257, 32'sd-0.09949962389929855, 32'sd-0.07325627988438824, 32'sd0.05558288401089113, 32'sd0.04253747183129651, 32'sd0.05431699008310907, 32'sd0.0634818992718554, 32'sd-0.09628275502139967, 32'sd-0.04631483797668264, 32'sd-0.09702891538619318, 32'sd-0.035232152689866215, 32'sd0.013429355892641395, 32'sd0.013270583167984185, 32'sd-0.052583128447642895, 32'sd-0.01773444807724757, 32'sd0.10864936812487072, 32'sd-0.08467146505016808, 32'sd0.018533888644202124, 32'sd0.00012674227261259653, 32'sd0.031306765772626255, 32'sd0.15734857004582514, 32'sd-0.013017460267727673, 32'sd-0.04140584264614635, 32'sd-0.07011876300128625, 32'sd0.0242511391116603, 32'sd-0.0030911945556490444, 32'sd0.08649345444312613, 32'sd0.1190721119707497, 32'sd-0.0063728825904779875, 32'sd0.03155897970402238, 32'sd-0.047724851139399206, 32'sd0.011758812912287985, 32'sd0.05853051712638161, 32'sd-0.08054295661974546, 32'sd-0.00436659152427751, 32'sd-0.02321761288968633, 32'sd-0.002692525159820374, 32'sd-0.06585127744565615, 32'sd-1.0570458885901404e-124, 32'sd-0.08111316260639656, 32'sd-0.08332725323912064, 32'sd0.014663740496330853, 32'sd0.019894883581029945, 32'sd0.053298384643170535, 32'sd-0.07370086270627521, 32'sd-0.06252693171772997, 32'sd0.1784825446775578, 32'sd0.1178381076922565, 32'sd0.0945128823579022, 32'sd-0.06334333544080163, 32'sd-0.06886537294681572, 32'sd0.02345876836900365, 32'sd-0.13730905881207234, 32'sd-0.12631605602243007, 32'sd-0.06598230586781494, 32'sd-0.006842809156255787, 32'sd-0.017084153648255513, 32'sd-0.020122761833662444, 32'sd-0.12925274244248788, 32'sd-0.1331820256536211, 32'sd-0.013555806200749436, 32'sd0.041078837434469676, 32'sd-0.0026259252923565707, 32'sd0.06317763990157936, 32'sd-0.053372814496766535, 32'sd-0.01094096859353884, 32'sd-0.0348224293615272, 32'sd-0.0737814332073646, 32'sd-0.08924614525762324, 32'sd-0.0514616152214171, 32'sd0.10742180952689492, 32'sd0.11154087084991422, 32'sd0.06878783465707697, 32'sd0.06035833842888535, 32'sd0.13757159689412965, 32'sd0.11229324743191127, 32'sd0.04201411318227669, 32'sd0.07676847025382831, 32'sd-0.09622887958854462, 32'sd0.06628074124774684, 32'sd-0.019083825770718304, 32'sd-0.045919967544391795, 32'sd-0.13581960582628277, 32'sd-0.0396172929801887, 32'sd-0.05731850153719533, 32'sd-0.02474234127894753, 32'sd-0.14785725204493294, 32'sd-0.12228662984506775, 32'sd0.06528121472620042, 32'sd-0.04313778732094086, 32'sd-0.11606728044819149, 32'sd-0.02604392392189518, 32'sd0.1459277035352008, 32'sd0.0076423728870005335, 32'sd-0.042690216421459426, 32'sd-0.08810475735824971, 32'sd0.04387567876854444, 32'sd0.02217193033493629, 32'sd0.09969658121537599, 32'sd0.042250871214294224, 32'sd0.01754964208677321, 32'sd0.09238404975579807, 32'sd0.05631433991723292, 32'sd-0.00048335096102820885, 32'sd0.13393685377172007, 32'sd0.09426992920998471, 32'sd0.035073201132698954, 32'sd0.1544762037147378, 32'sd0.05784476324258017, 32'sd-0.03105297080196578, 32'sd-0.03656836442361695, 32'sd-0.04058947277775399, 32'sd-0.034553068801807585, 32'sd-0.10361991731227228, 32'sd-0.14006559543666294, 32'sd-0.14432328590496046, 32'sd-0.11494769176041474, 32'sd-0.06664710672164488, 32'sd0.03786985469370538, 32'sd0.07464593142774714, 32'sd0.06292043215975782, 32'sd0.042019879506292504, 32'sd-1.7280299950196674e-117, 32'sd-0.02318794946088284, 32'sd0.020615254199615872, 32'sd-0.03935067411669348, 32'sd-0.012652738050727775, 32'sd0.07521692886306246, 32'sd0.0027854495461130066, 32'sd0.05025329468904218, 32'sd0.1655962156133067, 32'sd-0.058692348910150516, 32'sd-0.07759403357572446, 32'sd0.09283209543008708, 32'sd0.0021241642003439606, 32'sd-0.050364937858894565, 32'sd0.08319675421228183, 32'sd-0.02486112927540122, 32'sd0.0678549705660107, 32'sd-0.002445028506487522, 32'sd-0.06964271470011282, 32'sd-0.04506071703654212, 32'sd-0.17096502998189916, 32'sd-0.06915261971026572, 32'sd-0.03694086691938504, 32'sd0.010797709250835298, 32'sd0.060624503331951636, 32'sd0.07672421719684805, 32'sd-0.04976356626967489, 32'sd-1.389027684420969e-126, 32'sd-8.299497508811522e-123, 32'sd1.357733763935336e-115, 32'sd0.02206044353787575, 32'sd0.02366971518720236, 32'sd0.004450493634824555, 32'sd0.07046417132187792, 32'sd0.005992941939074019, 32'sd-0.042246384124837284, 32'sd0.08954541522668891, 32'sd-0.03410593613935731, 32'sd-0.07797650804001037, 32'sd-0.0179048841837472, 32'sd-0.033811659952550574, 32'sd0.01759070818879421, 32'sd-0.046563033325417585, 32'sd0.02109222344507677, 32'sd-0.0527556411780585, 32'sd-0.2160691816454498, 32'sd-0.16073469011455419, 32'sd-0.08169296839902108, 32'sd-0.03129120634137495, 32'sd-0.024900513933804894, 32'sd0.04800307879911911, 32'sd-0.010197211857417583, 32'sd0.051689999232486745, 32'sd-0.03932249353859073, 32'sd-0.04421724553326613, 32'sd2.3609597862370944e-114, 32'sd3.776968257200385e-115, 32'sd-4.704587049226724e-126, 32'sd0.01783437437516339, 32'sd-0.05857297281910527, 32'sd-0.07979791654475807, 32'sd-0.014120618182871202, 32'sd0.02722143697760675, 32'sd-0.02518287647708035, 32'sd0.034004190590855944, 32'sd-0.08464709322287806, 32'sd0.07184453400909317, 32'sd0.027378520136851752, 32'sd-0.015817000477970872, 32'sd-0.1338680509367708, 32'sd-0.08285985356838625, 32'sd-0.00777330616099218, 32'sd-0.06445444698450975, 32'sd-0.03331698454418441, 32'sd0.01727687724316165, 32'sd-0.08619186933149636, 32'sd-0.09059325863467659, 32'sd-0.11383323615187248, 32'sd-0.02848537421101515, 32'sd-0.12432235215822217, 32'sd-0.08103073086104236, 32'sd-0.06891761014179996, 32'sd-0.052984304191549404, 32'sd1.6318871287287622e-115, 32'sd1.0621712553482772e-119, 32'sd1.6816080152083816e-128, 32'sd-2.3985973506319753e-119, 32'sd-0.029029054323559247, 32'sd0.018736061530886944, 32'sd-0.017227999228184358, 32'sd-0.03399060974686827, 32'sd-0.02091942580152406, 32'sd0.11256255074466053, 32'sd0.05856402821711964, 32'sd0.06854280978917072, 32'sd0.10585653856087125, 32'sd0.03984953101145895, 32'sd0.05958859607228717, 32'sd0.004673878005024351, 32'sd-0.03420874181489591, 32'sd-0.008829658504148859, 32'sd-0.028167042649506438, 32'sd-0.12906320154406953, 32'sd0.0008342733819781765, 32'sd-0.10051810316018193, 32'sd-0.07733877187340422, 32'sd0.08407468901518629, 32'sd-0.018244354877306714, 32'sd0.02909755924352922, 32'sd0.018996934426268132, 32'sd-3.48852315619757e-114, 32'sd2.344183894960258e-123, 32'sd-2.13968324241031e-116, 32'sd-1.9715583814987443e-122, 32'sd-2.3554099361244685e-125, 32'sd1.0233187894930553e-122, 32'sd-0.05741607301377898, 32'sd-0.048164036838980684, 32'sd0.007240538401163737, 32'sd0.010895118174739156, 32'sd0.06305589361865065, 32'sd-0.07357938513136116, 32'sd-0.003566762704913977, 32'sd-0.005547179730446774, 32'sd0.013606009166780664, 32'sd0.037527230737264855, 32'sd0.062024447194153336, 32'sd-0.09195464081721764, 32'sd0.05458063983272703, 32'sd0.043456212977804574, 32'sd-0.10989668993141519, 32'sd0.001160607718019869, 32'sd-0.061046308792807334, 32'sd-0.04824400528991385, 32'sd0.028574821286521862, 32'sd0.0018766570383119718, 32'sd2.028971942982214e-121, 32'sd-2.2657625322449532e-122, 32'sd8.387968867695934e-117, 32'sd7.539230687522783e-119},
        '{32'sd7.956911643420058e-120, 32'sd-6.595840769246719e-126, 32'sd-2.1290331776155188e-114, 32'sd-1.4447205801750522e-124, 32'sd-5.6699677858517104e-120, 32'sd-1.964917699817407e-127, 32'sd1.1785155431838853e-122, 32'sd1.630397285586774e-115, 32'sd3.939266321243402e-124, 32'sd1.0876151710506796e-121, 32'sd2.3209815143198e-121, 32'sd3.44560595915516e-116, 32'sd-0.07898092709972393, 32'sd0.024192268021244374, 32'sd0.009952126339669033, 32'sd-0.08051300046242427, 32'sd-1.5907295083830632e-126, 32'sd1.0088034613319927e-117, 32'sd3.9626744029373137e-119, 32'sd8.63363738559585e-127, 32'sd-8.704245412453816e-121, 32'sd-4.5417926330638005e-116, 32'sd-4.0263429340540245e-120, 32'sd-6.507147569420044e-125, 32'sd5.878512799731871e-127, 32'sd-1.3451062983113544e-125, 32'sd-2.3423622434580955e-122, 32'sd-1.331732454919781e-122, 32'sd3.0079158689558335e-117, 32'sd-1.385243489906485e-118, 32'sd-8.014410360044079e-121, 32'sd5.29537951214097e-118, 32'sd-0.03579927596548162, 32'sd-0.0765694832143005, 32'sd0.06361753334596981, 32'sd0.12892058591769984, 32'sd-0.051688668299608824, 32'sd0.02216235296353618, 32'sd0.001965157935920164, 32'sd0.08044002581219384, 32'sd0.07611051107828176, 32'sd-0.1042916852054667, 32'sd-0.025159826919866995, 32'sd-0.018031751626983224, 32'sd0.02912963806146659, 32'sd0.019156038665880462, 32'sd0.055261318446048244, 32'sd-0.04337889320862092, 32'sd0.02226321861540348, 32'sd-0.05199610250800714, 32'sd0.02847730554858039, 32'sd-0.010217695182697184, 32'sd-1.1580465825472153e-128, 32'sd-1.248526929875723e-125, 32'sd-2.941966786349093e-126, 32'sd1.5441267861274098e-128, 32'sd-2.0795325288962735e-121, 32'sd1.2493534870369123e-122, 32'sd-0.04379311267264248, 32'sd-0.06247678374638399, 32'sd0.06012898968166405, 32'sd-0.05756614475299001, 32'sd-0.02240274690552521, 32'sd0.02190566033115605, 32'sd-0.03546471142888159, 32'sd-0.10089727480686084, 32'sd-0.07424285161307978, 32'sd0.08995928948126336, 32'sd0.012239535664622683, 32'sd0.011017607333443487, 32'sd-0.041964228934812456, 32'sd-0.014549993041639068, 32'sd-0.08236378344206076, 32'sd0.022239216451689626, 32'sd-0.014624406586261782, 32'sd-0.06085443574175712, 32'sd-0.006309446254074743, 32'sd-0.05334335381545766, 32'sd0.034871435862850235, 32'sd0.012345943905142992, 32'sd-0.04442996815835932, 32'sd-0.023394477460509176, 32'sd-5.692701734814072e-123, 32'sd-1.767490332663955e-120, 32'sd-1.0596731313027533e-125, 32'sd1.5167503831249051e-124, 32'sd-0.02788233229420824, 32'sd0.046107464604322405, 32'sd0.0964740569792447, 32'sd0.06611347138257649, 32'sd0.11097460276355037, 32'sd-0.06985635140754591, 32'sd-0.05801942658904468, 32'sd-0.030913784256982907, 32'sd-0.046785119997786284, 32'sd0.0018325099849727114, 32'sd-0.1076214015595564, 32'sd0.04002918872284716, 32'sd-0.010030061828881408, 32'sd-0.0846321632321558, 32'sd0.04028593083681204, 32'sd-0.0058886901155342855, 32'sd0.13947376324928099, 32'sd0.04953830043953986, 32'sd-0.06755192812610582, 32'sd0.07641643102223779, 32'sd-0.03335578914887611, 32'sd-0.007484431280981688, 32'sd-0.05900397461044548, 32'sd-0.09451729769108226, 32'sd0.004890157842510806, 32'sd1.109008324488311e-119, 32'sd8.250360761855689e-117, 32'sd-0.029798728029244038, 32'sd-0.013727729902996342, 32'sd-0.04542683065928913, 32'sd0.05132680336744512, 32'sd0.025384560858181294, 32'sd-0.012613038189675178, 32'sd0.03478763870821145, 32'sd-0.025705920426670525, 32'sd0.07054519794192511, 32'sd-0.08845312752888804, 32'sd-0.029076974396755557, 32'sd-0.048029588432562484, 32'sd0.026873492979737568, 32'sd-0.047606287540172, 32'sd-0.014535590718375452, 32'sd0.07605365374592966, 32'sd-0.06474122061207842, 32'sd0.08387974555371737, 32'sd0.023443936350364986, 32'sd-0.04844359690906459, 32'sd0.09422725569735896, 32'sd0.12699485374592165, 32'sd-0.008051313913116894, 32'sd-0.001954038469143548, 32'sd0.010323063783852776, 32'sd-0.06105078062718772, 32'sd0.0761601961592541, 32'sd-8.09532132168115e-117, 32'sd-0.03060702537669834, 32'sd0.030848851151644992, 32'sd0.044087175052187115, 32'sd-0.0494925290588597, 32'sd-0.07947283021872438, 32'sd0.041970301435973724, 32'sd0.12709210449393935, 32'sd0.09922641765302151, 32'sd0.11072579793608117, 32'sd0.11026579204850491, 32'sd-0.04940607915393343, 32'sd-0.10637109565838057, 32'sd-0.02047502569654905, 32'sd-0.05340047966876576, 32'sd-0.05581570651522466, 32'sd0.1380772573595709, 32'sd0.13744312520512178, 32'sd-0.02656895756546543, 32'sd0.017970990699036113, 32'sd-0.04259949883570405, 32'sd0.13975502692815595, 32'sd0.1628625901810996, 32'sd0.03799515749277671, 32'sd-0.06166104707131162, 32'sd-0.08150612802956285, 32'sd0.007608312694740643, 32'sd-0.07870700556675722, 32'sd1.314202602907481e-118, 32'sd-0.004363332940665506, 32'sd-0.00847796903291138, 32'sd-0.06275891070043332, 32'sd0.05088544766213451, 32'sd0.04017267369064744, 32'sd0.03508933181439315, 32'sd0.1259515014906039, 32'sd0.045413730182431604, 32'sd0.13182752882853618, 32'sd0.07018987112788722, 32'sd-0.00943026236262806, 32'sd-0.0012120424540389297, 32'sd0.06096384595943682, 32'sd0.06496464995827422, 32'sd-0.012445458549515788, 32'sd-0.06987670732222553, 32'sd0.08110787838070001, 32'sd0.10643444482336048, 32'sd0.03957865802088402, 32'sd-0.03342659722164953, 32'sd0.04125355494640726, 32'sd0.11097415884935168, 32'sd0.1132571232434333, 32'sd-0.009839670543340442, 32'sd0.05877262836064531, 32'sd-0.011596921448973197, 32'sd0.04815159004607788, 32'sd0.0327291824508857, 32'sd0.005844614819981312, 32'sd0.010289347955793126, 32'sd0.002252145260233085, 32'sd-0.08729473383000577, 32'sd0.07230117303638128, 32'sd0.02626052950705052, 32'sd0.008142576861916048, 32'sd0.20136925201446457, 32'sd0.0803006032158673, 32'sd0.11293745921152804, 32'sd-0.0075416708060552055, 32'sd0.004449837202173015, 32'sd-0.08953539310422118, 32'sd-0.018471091471476003, 32'sd0.06837832933736511, 32'sd0.021543127558186718, 32'sd0.0681173609902029, 32'sd0.08767665990927809, 32'sd0.018253410731752188, 32'sd-0.043382892542663684, 32'sd0.13727959970580364, 32'sd0.08689546360904796, 32'sd0.09763502946777344, 32'sd-0.02852037372511896, 32'sd-0.04349439547712762, 32'sd-0.05028696173156692, 32'sd-0.049687452273404716, 32'sd-0.034996322407146646, 32'sd-0.022898806732778595, 32'sd0.0191499982395949, 32'sd0.035978009158104785, 32'sd0.003367873037111437, 32'sd0.008242486507268007, 32'sd0.08921288358080809, 32'sd0.011650616634101971, 32'sd0.06981445518825079, 32'sd0.1165506465200196, 32'sd-0.09632548405473802, 32'sd0.017821928052045456, 32'sd0.016315720417847235, 32'sd-0.0008560954214266019, 32'sd-0.028692865184598144, 32'sd-0.04062530101581279, 32'sd-0.0603402851246396, 32'sd0.015366936421438071, 32'sd-0.06595302973032226, 32'sd-0.03171547847238518, 32'sd0.05297105861382338, 32'sd0.010591166584715591, 32'sd0.010419608834120974, 32'sd0.04461421975652981, 32'sd-0.06876606150531477, 32'sd0.053998480473139016, 32'sd-0.11638703736542164, 32'sd0.03678798608057054, 32'sd-0.026546973703051598, 32'sd-0.08220113424847784, 32'sd-0.02711348781312651, 32'sd0.04262597142767818, 32'sd-0.050582167459352415, 32'sd-0.051194546904350005, 32'sd-0.09904566794512723, 32'sd0.09362160720127487, 32'sd0.16332447891967827, 32'sd0.11839506485000761, 32'sd0.11088596186175834, 32'sd0.0017259559098775842, 32'sd0.024644673021032387, 32'sd-0.11613584242128072, 32'sd-0.2343889546017405, 32'sd-0.04839866759179928, 32'sd-0.1092175548997519, 32'sd-0.040303305907888755, 32'sd-0.048816426283066094, 32'sd0.08119910668357522, 32'sd-0.08703941377467682, 32'sd0.03552294881188038, 32'sd0.013509660727298317, 32'sd0.07194947421676343, 32'sd0.04367461303336712, 32'sd-0.02848932949105788, 32'sd0.04142948453082828, 32'sd-0.018528443105412826, 32'sd0.010658371842673868, 32'sd0.03230587941036538, 32'sd-0.009133051608202103, 32'sd-0.05870609797930688, 32'sd0.00909302456025894, 32'sd0.11664919871737824, 32'sd-0.022010170786855715, 32'sd0.046790871589953424, 32'sd-0.007232857377749672, 32'sd0.08645218123544209, 32'sd0.08651973474858171, 32'sd0.029154881889853233, 32'sd-0.07377326259021096, 32'sd-0.11507781623874787, 32'sd-0.13914567931370966, 32'sd-0.11844786056828518, 32'sd-0.1409749647981073, 32'sd-0.1163798642834229, 32'sd0.029824704087110313, 32'sd-0.004017662127236074, 32'sd-0.05725895072503947, 32'sd0.14449829909413398, 32'sd0.12274451761835406, 32'sd0.10721909830094765, 32'sd0.067935878787004, 32'sd0.02275960437535844, 32'sd0.010888563124585693, 32'sd0.05651024080568061, 32'sd-0.016223118524873844, 32'sd-0.05330549198866204, 32'sd-0.013342194647748103, 32'sd-0.08806222159013607, 32'sd0.1001264615516594, 32'sd0.05515118254661422, 32'sd-0.08372098987766056, 32'sd-0.02634133328620043, 32'sd-0.05195461230262112, 32'sd-0.03931580115462239, 32'sd0.09190264642640708, 32'sd0.12473196979937949, 32'sd0.006020325947487497, 32'sd0.057153318920526115, 32'sd-0.004618722445040058, 32'sd-0.1912009182101151, 32'sd-0.20204104416858468, 32'sd-0.10975834555495148, 32'sd-0.24497271974611665, 32'sd0.07126558982142395, 32'sd0.0173855504909438, 32'sd-0.08000968639530018, 32'sd-0.12313123266301101, 32'sd-0.19353570126422565, 32'sd0.02851862398222894, 32'sd-0.051103044637299574, 32'sd0.09475600324455252, 32'sd-0.10227384295117234, 32'sd0.0375411688233817, 32'sd-0.07678682301814471, 32'sd0.019709582144260992, 32'sd-0.02922689695493449, 32'sd-0.035624589236172066, 32'sd0.09513017670072291, 32'sd0.04760414064414967, 32'sd0.03153251855497592, 32'sd0.037211589243752, 32'sd0.07520727097470624, 32'sd0.11698284839778554, 32'sd0.13423252369515512, 32'sd0.13273743659902856, 32'sd-0.05388470468712895, 32'sd-0.0913005514324421, 32'sd-0.3217443626360329, 32'sd-0.13778226169508134, 32'sd-0.16036978645607466, 32'sd-0.03319616768747822, 32'sd-0.03809401502076081, 32'sd-0.09350669005586025, 32'sd0.014968541785263556, 32'sd-0.16139972249287582, 32'sd-0.10527329015513005, 32'sd0.07288782173910832, 32'sd0.041722251120916376, 32'sd0.0914051270214561, 32'sd-0.03939368129747455, 32'sd0.051508953962284235, 32'sd-0.010142811535962377, 32'sd-0.10206959419570001, 32'sd0.012212101309951474, 32'sd-0.04030806420402973, 32'sd0.04992991239614689, 32'sd0.030829505569780535, 32'sd0.018060994273527656, 32'sd0.033722622268138304, 32'sd0.14144866501599415, 32'sd0.008072429992441236, 32'sd0.10820234031594594, 32'sd0.08478401779320037, 32'sd0.021710152625833028, 32'sd-0.2266332411885391, 32'sd-0.19946864783088702, 32'sd-0.13413198003525903, 32'sd-0.12124783204332493, 32'sd0.03600300494882191, 32'sd-0.040912089790170386, 32'sd-0.07807084202184571, 32'sd-0.0883400530066564, 32'sd-0.04809336415246404, 32'sd0.04063068963139013, 32'sd-0.012753280120335816, 32'sd0.04808763682444031, 32'sd0.024396442274939426, 32'sd0.033083259200067494, 32'sd0.12112187602924054, 32'sd0.027804949746890014, 32'sd-0.0038439653351310474, 32'sd0.04845746628453988, 32'sd0.04802880816302957, 32'sd-0.08039535659270838, 32'sd0.011438214906790846, 32'sd-0.010750766146780224, 32'sd-0.008473993955900132, 32'sd-0.018834130604424373, 32'sd0.053668204831815045, 32'sd0.13603712291357592, 32'sd0.10184235883305642, 32'sd0.0680820908355002, 32'sd-0.16019463418887855, 32'sd-0.20665583208866825, 32'sd0.01989458163815459, 32'sd-0.05540729418673343, 32'sd-0.011419271964380783, 32'sd-0.15355762769611242, 32'sd-0.10724373311115508, 32'sd-0.0018231300042441379, 32'sd0.008246881235627373, 32'sd0.07310693385429025, 32'sd-0.03280910124473916, 32'sd0.012129953556107746, 32'sd0.03452574981254896, 32'sd0.04462448953837841, 32'sd-0.026699372683909425, 32'sd0.02046295402648755, 32'sd0.04197517195485763, 32'sd-0.09156646948313957, 32'sd-0.031118075770718318, 32'sd-0.016974319211070794, 32'sd-0.008293941480716605, 32'sd0.045811986256349545, 32'sd-0.005575730039005643, 32'sd0.026446166988775697, 32'sd-0.051014580533256006, 32'sd0.090098117752639, 32'sd0.1980711615495655, 32'sd0.11958853269051331, 32'sd0.06315323213860657, 32'sd0.06912298916930293, 32'sd0.005278771696241008, 32'sd-0.061854957865337956, 32'sd-0.10537728269457626, 32'sd-0.1966656778611749, 32'sd-0.19453420191155646, 32'sd-0.09036301869983734, 32'sd-0.11743205121325197, 32'sd-0.006284563575595789, 32'sd-0.009178068448177304, 32'sd0.0020270822853949762, 32'sd-0.008505778411456081, 32'sd0.06235291021666413, 32'sd0.03587028856178332, 32'sd-0.04953090069354394, 32'sd0.11185986269661019, 32'sd-0.056246798757640305, 32'sd-0.058403789996360166, 32'sd-0.06875940599205986, 32'sd-0.04465018204324331, 32'sd-0.15964226361306358, 32'sd-0.1428340818461921, 32'sd-0.030131630613534875, 32'sd0.016578731427375308, 32'sd0.0032104871506440946, 32'sd0.04674381701962088, 32'sd0.13591060568764352, 32'sd0.08097590023278967, 32'sd-0.03239521913366543, 32'sd-0.09126936252231857, 32'sd-0.049373863008491364, 32'sd-0.15440550901267325, 32'sd0.009953410025605637, 32'sd-0.12790645284472907, 32'sd-0.06565759840784396, 32'sd-0.04724023537595767, 32'sd0.0384567621798579, 32'sd0.0058520569687383305, 32'sd0.05227297845220095, 32'sd-0.062081148357311315, 32'sd-0.04196088175505578, 32'sd1.2582617203110214e-115, 32'sd-0.006776975707248803, 32'sd0.04185641568955263, 32'sd-0.08127768742995745, 32'sd-0.03686726295605555, 32'sd-0.06470996209720127, 32'sd-0.03959532387541583, 32'sd-0.19205802959711984, 32'sd-0.1186158083496259, 32'sd-0.0834438955576332, 32'sd0.04672415822194621, 32'sd0.03750741779004929, 32'sd0.22041813286173376, 32'sd0.1952948991327719, 32'sd0.08795679612993493, 32'sd0.0005111487211531683, 32'sd-0.032032237465094586, 32'sd-0.20786379039389233, 32'sd-0.1097638914286889, 32'sd-0.0422806133194355, 32'sd-0.04350576539331243, 32'sd0.0487206170150648, 32'sd0.17668217872858724, 32'sd0.10248488666296003, 32'sd-0.0015897214305791443, 32'sd-0.10207930996500904, 32'sd-0.07263521350057127, 32'sd0.0061196493259551765, 32'sd-0.030199002225319436, 32'sd-0.011593341939750942, 32'sd0.019913652868298142, 32'sd-0.0519974960576089, 32'sd0.015513963337903587, 32'sd-0.08043793958356948, 32'sd-0.0332443020846655, 32'sd-0.17349573983851885, 32'sd-0.11742107564198234, 32'sd-0.060057198622490676, 32'sd-0.061443377267066404, 32'sd-0.07684529380162229, 32'sd0.16540864542563877, 32'sd0.033713041897942025, 32'sd-0.035055646003394336, 32'sd0.008389654562595612, 32'sd-0.14581966251251693, 32'sd-0.17863457859612678, 32'sd-0.13668148360648816, 32'sd-0.0406143998408626, 32'sd0.05134328050325794, 32'sd0.024905055434421033, 32'sd0.07411106656779796, 32'sd-0.017279135498748675, 32'sd0.051320979885955034, 32'sd0.03050232761224155, 32'sd-0.07450793366610986, 32'sd-0.02781766335205377, 32'sd-0.0392183248904462, 32'sd0.008316174029712221, 32'sd0.01082616448054176, 32'sd0.08001742199289377, 32'sd-0.0850963017971517, 32'sd-0.00982589084459442, 32'sd-0.0970165006497301, 32'sd0.034124215869513724, 32'sd-0.10680268107729841, 32'sd-0.15100858740818202, 32'sd-0.059366796295896286, 32'sd-0.12183210735323403, 32'sd0.18363822508539288, 32'sd-0.0899870342519044, 32'sd-0.2182481619189695, 32'sd-0.16175087424965232, 32'sd-0.05478016915013197, 32'sd0.09076049620935396, 32'sd0.046956024446574984, 32'sd0.017714637445339496, 32'sd0.07051820314413762, 32'sd0.12796473904054856, 32'sd-0.019424488731551847, 32'sd-0.005121944911815674, 32'sd0.08839755809534668, 32'sd0.005751767553046695, 32'sd-0.05383279076114165, 32'sd0.0031278021338657447, 32'sd-1.4226719504704986e-118, 32'sd0.09268061051276846, 32'sd0.050638410005708345, 32'sd0.039998544490379914, 32'sd0.006477763961727738, 32'sd-0.05332286963705516, 32'sd0.05609069154713753, 32'sd0.0014924888156899589, 32'sd0.018869851325926695, 32'sd-0.07795059438092573, 32'sd0.07622888676981787, 32'sd0.04519124634589624, 32'sd0.06483929418915241, 32'sd-0.1306598167639222, 32'sd-0.13186936514785733, 32'sd0.057738448992937244, 32'sd0.04373488295232983, 32'sd0.10722737491712137, 32'sd0.1328481414078918, 32'sd0.06769613510127871, 32'sd0.12388493081099292, 32'sd0.008006033093732615, 32'sd-0.0688096366236844, 32'sd0.01717014658579997, 32'sd0.07877707467320581, 32'sd0.022192422180331524, 32'sd-0.015358998233811417, 32'sd0.005087901815992493, 32'sd-0.02482646987611031, 32'sd0.05373514984389989, 32'sd0.01350135196068744, 32'sd-0.03549690977166866, 32'sd0.04831887191607537, 32'sd-0.029816609897109648, 32'sd-0.016559241118535534, 32'sd0.04891483022748273, 32'sd0.022842405121332794, 32'sd0.016514972893219796, 32'sd0.10150468022301082, 32'sd-0.03547904991563744, 32'sd-0.06256850061642215, 32'sd-0.058152794033773055, 32'sd-0.016963625702380313, 32'sd0.051467211951274655, 32'sd0.018845558138977866, 32'sd0.1284503453160053, 32'sd0.08981246313392094, 32'sd0.13159970360788495, 32'sd0.13916612236708156, 32'sd0.11248247749387448, 32'sd0.05767208043417523, 32'sd0.017079407576664006, 32'sd-0.032125071529427576, 32'sd-0.012093737786378404, 32'sd0.051939160877432, 32'sd-0.03922508088719163, 32'sd0.00044568531122440933, 32'sd-0.054594383177302586, 32'sd0.047635900483998336, 32'sd0.08135122772123941, 32'sd0.028037971760096828, 32'sd-0.04018545712510407, 32'sd0.0017334391085350837, 32'sd0.026896105813655355, 32'sd0.004508045081548711, 32'sd0.03582568837107499, 32'sd-0.07702554008345665, 32'sd0.10585754332961379, 32'sd0.054512359830602514, 32'sd0.04189664533457268, 32'sd0.024472003985655702, 32'sd0.13136321841707838, 32'sd0.11085837242041201, 32'sd0.2278336064777484, 32'sd0.1690982563770175, 32'sd0.03313787512535816, 32'sd0.07359080909587355, 32'sd0.04176842342659196, 32'sd0.05214548822131643, 32'sd0.007695776786444667, 32'sd0.0080760751853259, 32'sd0.025251522109381568, 32'sd0.01002485127077231, 32'sd0.04210307869879778, 32'sd-1.834146041228116e-123, 32'sd0.04651708324372418, 32'sd-0.014999375008429376, 32'sd0.1322391006727333, 32'sd0.014245736351932712, 32'sd-0.03918424028578888, 32'sd-0.03903965236190409, 32'sd0.03129152775495993, 32'sd0.02192119809828099, 32'sd-0.05901013679994921, 32'sd-0.030958621430765585, 32'sd-0.007361940945723332, 32'sd0.14842446956892846, 32'sd0.10277764562390758, 32'sd0.054406714307888765, 32'sd0.1930202409322209, 32'sd0.20992455381274563, 32'sd0.13506627747646696, 32'sd0.14045248666707402, 32'sd0.04715888608426747, 32'sd0.08373324244633286, 32'sd0.037525517935562185, 32'sd0.08340186954145203, 32'sd0.05050659471461861, 32'sd-0.031037269687764504, 32'sd0.09475120655803712, 32'sd0.0721208172900591, 32'sd-4.4018661606425747e-122, 32'sd-3.2676203117921696e-121, 32'sd2.466865043528654e-120, 32'sd-0.019967347226287194, 32'sd0.07485625238712225, 32'sd0.0012884804382443536, 32'sd-0.04558869390484455, 32'sd-0.1396811497298128, 32'sd-0.05493322123238028, 32'sd0.08737912278968271, 32'sd0.09354554994139024, 32'sd0.0818286733316744, 32'sd0.15426281449600082, 32'sd0.17684272299007772, 32'sd0.20049606758142113, 32'sd0.19455405828309996, 32'sd0.23947471575458018, 32'sd0.1389164779790135, 32'sd0.10828264192262155, 32'sd0.09130874448947139, 32'sd0.09952111635899963, 32'sd0.06457949839927553, 32'sd0.06697045683061015, 32'sd0.006933440601067088, 32'sd-0.08289418339608096, 32'sd-0.11549840945336218, 32'sd-0.10627340790561669, 32'sd-0.018085713565122834, 32'sd1.5177099433451146e-115, 32'sd-7.041702119828858e-117, 32'sd3.213762972144636e-124, 32'sd0.004326812886017693, 32'sd0.01296679204068734, 32'sd-0.04668387848411941, 32'sd-0.07544320523768304, 32'sd0.02583624528360803, 32'sd0.022441918500144296, 32'sd0.12238873471783306, 32'sd0.028001400872045137, 32'sd-0.02182698537576116, 32'sd0.10588566908628014, 32'sd0.07386378915993755, 32'sd0.0925488957548917, 32'sd0.09208282750940534, 32'sd0.0720912191816172, 32'sd0.06041240991924711, 32'sd0.07225914741475996, 32'sd0.013372300675798065, 32'sd-0.06246213323898211, 32'sd-0.012588204689199937, 32'sd-0.020323479177405686, 32'sd0.0660631257868719, 32'sd-0.06217964207431256, 32'sd-0.06819806074474942, 32'sd0.02072595462205333, 32'sd-0.03534155484242456, 32'sd-2.4538928238210506e-126, 32'sd-1.0602954333220917e-127, 32'sd-6.65571441992575e-126, 32'sd4.1898083736864103e-125, 32'sd-0.014044092888181042, 32'sd0.01933274413707329, 32'sd-0.0719828872862894, 32'sd-0.06903256226997333, 32'sd0.0032874905465628997, 32'sd-0.03953328506674447, 32'sd0.01681731162803591, 32'sd-0.015552697528599436, 32'sd-0.0008524089407557698, 32'sd0.07443703777807338, 32'sd0.0988895554689115, 32'sd-0.07223092225078431, 32'sd0.047404771458684596, 32'sd0.015266863409145454, 32'sd-0.011436374336461549, 32'sd-0.008219533483489461, 32'sd-0.06246147051930873, 32'sd0.06374630771491349, 32'sd-0.008415563231781597, 32'sd-0.023161889095266765, 32'sd-0.018480943077889993, 32'sd-0.0023605387877858094, 32'sd-0.03857457420227266, 32'sd-2.116107760681473e-117, 32'sd4.392550980742641e-126, 32'sd-4.140205290289721e-117, 32'sd-1.0774153975547105e-125, 32'sd-6.388691031043862e-119, 32'sd2.533256043516194e-126, 32'sd0.025100763976502207, 32'sd0.0029237210807736046, 32'sd-0.04565437503362735, 32'sd0.08050492103201909, 32'sd0.024917142143254446, 32'sd0.0645956959440237, 32'sd-0.0054791300348257755, 32'sd-0.025353178207857176, 32'sd0.03974749609321751, 32'sd0.02324676368463316, 32'sd-0.011831870868295237, 32'sd-0.043553626077677536, 32'sd-0.031134379556624694, 32'sd0.031868404753482106, 32'sd0.03861141974601928, 32'sd-0.028854768814252578, 32'sd-0.019049979252498017, 32'sd-0.0244463339759657, 32'sd-0.05292952507531527, 32'sd0.0017539754803343117, 32'sd2.939077010782581e-116, 32'sd1.5903282710685132e-127, 32'sd3.8369501877420013e-119, 32'sd2.884683398838237e-116},
        '{32'sd-5.157293655288435e-119, 32'sd9.916271153144517e-121, 32'sd-2.5140579120046628e-126, 32'sd2.5139995544897284e-116, 32'sd-1.5204885689284832e-124, 32'sd6.178680750348032e-119, 32'sd1.7160984183262052e-123, 32'sd2.975345377601722e-124, 32'sd-1.143488856427244e-116, 32'sd6.128336888707011e-126, 32'sd-1.818759038456638e-123, 32'sd8.6793750463479e-118, 32'sd0.004746853889246333, 32'sd0.08300865513536959, 32'sd0.05298436529982529, 32'sd0.08101889824436932, 32'sd3.376310211802032e-123, 32'sd-2.519162461249735e-125, 32'sd8.67978972009326e-121, 32'sd1.0097413016972184e-120, 32'sd-2.1535479160105312e-127, 32'sd3.960071045228798e-119, 32'sd-1.2198620333555577e-122, 32'sd3.057253851817317e-125, 32'sd-6.4204685781490805e-124, 32'sd-3.235926778045225e-122, 32'sd-4.8615080511629585e-117, 32'sd-6.845945684738761e-115, 32'sd-3.138454000015314e-119, 32'sd-1.8090062114795018e-117, 32'sd7.528348462868912e-118, 32'sd-2.0673716870611397e-129, 32'sd-0.05632275921383646, 32'sd0.027621093341412696, 32'sd0.07576151775488058, 32'sd0.09595686270074864, 32'sd0.058103724113618055, 32'sd0.08268808104814114, 32'sd0.018842257730703377, 32'sd-0.05304200990656846, 32'sd0.06358658116815934, 32'sd0.09363190749424995, 32'sd0.009458252700806889, 32'sd0.056672440183882476, 32'sd-0.07489087833786671, 32'sd0.05745567719320671, 32'sd0.0025686881462520113, 32'sd-0.020368346045866733, 32'sd0.013924441253868401, 32'sd0.016841910220205064, 32'sd-0.036054337761554325, 32'sd0.0031504581778766037, 32'sd-3.7642024404929516e-122, 32'sd-2.5863068289492494e-125, 32'sd3.611171210237963e-119, 32'sd1.9113447682492764e-114, 32'sd4.1146473439104104e-121, 32'sd-9.480542160035956e-123, 32'sd0.013431779027507515, 32'sd-0.03909082588699758, 32'sd0.01048754499027999, 32'sd-0.024339890196030327, 32'sd0.045923063627940006, 32'sd0.11611385910804255, 32'sd0.08464582118934057, 32'sd0.13412638802350452, 32'sd0.05111125050670305, 32'sd-0.020591220117705932, 32'sd-0.07219206257246137, 32'sd-0.07350624924903688, 32'sd0.0958826437556774, 32'sd-0.011975350278187382, 32'sd-0.06245207501709325, 32'sd0.03259788513149184, 32'sd-0.11048604806030775, 32'sd-0.09248364865900846, 32'sd-0.0005132153991580704, 32'sd0.017906315774739286, 32'sd0.009773418397401862, 32'sd0.11429866319494615, 32'sd0.022828598233202, 32'sd0.050289889594894124, 32'sd9.268440247820917e-125, 32'sd1.5669446753625302e-121, 32'sd-1.3947982529984633e-127, 32'sd2.5409308633692914e-120, 32'sd0.016259671764812147, 32'sd0.0046815959440476285, 32'sd-0.03382044631008816, 32'sd0.06338691095732787, 32'sd0.04515437683197708, 32'sd0.007610066895960023, 32'sd-0.05062894776864608, 32'sd-0.00895325457172144, 32'sd0.043274356354151014, 32'sd-0.01635853104934425, 32'sd0.05959325631902697, 32'sd-0.12588828971605517, 32'sd0.06562353745710227, 32'sd0.004851329175521719, 32'sd0.12663530910430285, 32'sd0.028177968668886916, 32'sd-0.10807256453393843, 32'sd0.024999030800360738, 32'sd0.03201220478746805, 32'sd0.10709967691816263, 32'sd-0.010183013599371135, 32'sd-0.052398715186788965, 32'sd-0.07968253486373357, 32'sd0.09084821662250725, 32'sd0.006145314575929346, 32'sd-1.360351222374455e-118, 32'sd1.681727581059299e-122, 32'sd0.04211836917873234, 32'sd-0.03589976582489864, 32'sd0.011429749513184867, 32'sd-0.005919165715619852, 32'sd-0.009327696691914904, 32'sd-0.03324176817230624, 32'sd-0.04500427721092858, 32'sd-0.12989650569953648, 32'sd-0.18047797620876896, 32'sd-0.13480152338735027, 32'sd-0.11931499193550908, 32'sd-0.11171099757629008, 32'sd0.005095826968571172, 32'sd0.0968870767998335, 32'sd0.09292070735662494, 32'sd0.09658805763755333, 32'sd0.07883256401010635, 32'sd-0.03809973105067377, 32'sd-0.08093587942692494, 32'sd0.12165896497709308, 32'sd0.07338325506863376, 32'sd-0.008775757191802484, 32'sd-0.03710591937848533, 32'sd-0.09644950083290003, 32'sd-5.878879347224479e-05, 32'sd0.015585086119461551, 32'sd-0.009416917250685474, 32'sd-1.3803739975366327e-125, 32'sd-0.0030496062310515133, 32'sd0.032060188307782546, 32'sd-0.06029484151203943, 32'sd0.05389869158498978, 32'sd0.03252487662563725, 32'sd0.07017180182691575, 32'sd-0.17253541089771152, 32'sd-0.13640621061021854, 32'sd-0.20472945675273777, 32'sd-0.08546539683606959, 32'sd-0.052060578273275745, 32'sd-0.050383899998717604, 32'sd0.05972990947781621, 32'sd0.07453438844487467, 32'sd0.030148075210400086, 32'sd0.1270430822593419, 32'sd0.15536080302373123, 32'sd0.046909190218913294, 32'sd0.06893495954243807, 32'sd0.015429751101453289, 32'sd-0.10317282052763758, 32'sd-0.06998431440007484, 32'sd-0.1230232730716536, 32'sd-0.09423406785206523, 32'sd0.028983233183064668, 32'sd0.013497737665621273, 32'sd-0.0384241255215276, 32'sd6.591979576198536e-124, 32'sd0.019060634205196787, 32'sd0.036906992409115935, 32'sd-0.08149203953736392, 32'sd-0.04751875249063364, 32'sd0.005561734042460748, 32'sd-0.051560264870149496, 32'sd-0.07515621002228147, 32'sd-0.1442727313894161, 32'sd-0.15541309453051413, 32'sd-0.08757479589252637, 32'sd-0.09429258144487956, 32'sd-0.040746043329211265, 32'sd-0.022650257853137658, 32'sd0.010788589998932006, 32'sd-0.05214281298824099, 32'sd-0.07674773068424087, 32'sd0.02700043008486763, 32'sd-0.13248997480539249, 32'sd0.004540400379594792, 32'sd-0.032492987954365345, 32'sd-0.11744033353916629, 32'sd0.011940324518624017, 32'sd0.07379268947739523, 32'sd0.05514819432181609, 32'sd-0.010322255398386649, 32'sd-0.00874151229075574, 32'sd-0.05459262879146759, 32'sd0.03602774580093371, 32'sd0.030415935930000738, 32'sd0.07197870233211447, 32'sd-0.03553772150367064, 32'sd0.020282673735702725, 32'sd-0.051365599223237315, 32'sd-0.08414914032138754, 32'sd-0.0953827668475112, 32'sd-0.045967688279239735, 32'sd-0.17296681224664529, 32'sd-0.05432770883080943, 32'sd0.005208646841490312, 32'sd-0.03836904673740063, 32'sd-0.03584985554703082, 32'sd0.03585470493557845, 32'sd-0.11123932567634688, 32'sd-0.11365233473360531, 32'sd-0.008091019083239696, 32'sd-0.14895802044778794, 32'sd-0.050449074551419844, 32'sd-0.05416651107751817, 32'sd-0.03871522167817937, 32'sd0.04496243144982514, 32'sd-0.034961248947794156, 32'sd0.050523440224556904, 32'sd-0.011047772427450394, 32'sd0.02318939594969527, 32'sd-0.06729641853107231, 32'sd0.012883948439925519, 32'sd0.023370987374149027, 32'sd0.05813263548277211, 32'sd-0.2090092050111403, 32'sd-0.06057860029363814, 32'sd-0.054911427608702594, 32'sd0.002181166246914267, 32'sd-0.0958315516592934, 32'sd-0.02002721666029509, 32'sd-0.06560811451053328, 32'sd-0.18411064224557688, 32'sd-0.0027739081519167004, 32'sd0.08093761547517915, 32'sd0.087901931429995, 32'sd0.03867399076615216, 32'sd0.018213595525445308, 32'sd-0.02375670317190229, 32'sd-0.13693247462028085, 32'sd-0.12067599685261174, 32'sd-0.11415431545647751, 32'sd-0.029890353240257454, 32'sd-0.02039283635988437, 32'sd-0.14133757501343913, 32'sd-0.03446138558199865, 32'sd-0.05479916125434881, 32'sd0.11070463542362118, 32'sd0.10981285505581287, 32'sd0.042167194567502134, 32'sd0.05074769926916587, 32'sd-0.009336305325970653, 32'sd-0.04264662625017002, 32'sd-0.08654346299254137, 32'sd-0.024851052186078845, 32'sd0.051362993476478845, 32'sd-0.057863941460374047, 32'sd0.01691775878488382, 32'sd-0.08212843050218817, 32'sd0.03947082256845058, 32'sd-0.1650388176521438, 32'sd-0.09913714261493581, 32'sd0.0873897556398726, 32'sd0.0014965314723924955, 32'sd-0.03931615936019704, 32'sd-0.001179648677310157, 32'sd-0.015188796897799174, 32'sd-0.09850403297954441, 32'sd-0.12156298725552789, 32'sd-0.07124773484942908, 32'sd-0.07686028328214198, 32'sd-0.060364084850322054, 32'sd-0.1286809799744428, 32'sd-0.14165505642055282, 32'sd-0.11007145925121002, 32'sd-0.08463043968884477, 32'sd0.032272889713436705, 32'sd-0.04951286682924544, 32'sd-0.030262763533891887, 32'sd-0.06889567269282224, 32'sd-0.06443234945985818, 32'sd-0.06859587117415462, 32'sd-0.0044867045540139885, 32'sd0.0576252317108493, 32'sd-0.016724111156286563, 32'sd0.10016559950101875, 32'sd0.07024192536887287, 32'sd-0.03904937625673222, 32'sd-0.04435284206017132, 32'sd-0.08262936554684319, 32'sd-0.08841170643788342, 32'sd-0.09411575332562021, 32'sd-0.08946346373364217, 32'sd-0.10350475277977646, 32'sd-0.03574501225991484, 32'sd-0.05513016521651629, 32'sd-0.004891946493693619, 32'sd-0.007705358705921043, 32'sd-0.09969456082766631, 32'sd-0.14037314214731533, 32'sd-0.07375598771253841, 32'sd-0.20257858069690313, 32'sd0.03481902134656224, 32'sd0.05968373518655309, 32'sd0.12941675894277246, 32'sd-0.027615883279887947, 32'sd-0.013789520256231829, 32'sd0.05654798501440152, 32'sd-0.02798929383755225, 32'sd-0.059839440846342226, 32'sd-0.021089669766127663, 32'sd-0.0316486220800896, 32'sd0.15721822235910557, 32'sd-0.004603042505043898, 32'sd0.1264636260238548, 32'sd-0.0471239899201313, 32'sd-0.046839771032600924, 32'sd-0.07851054545566465, 32'sd0.031463869914683605, 32'sd-0.11182878903638051, 32'sd-0.081580800568974, 32'sd-0.05282087626004399, 32'sd-0.04002520499114163, 32'sd0.00333099189260656, 32'sd0.10238042736072998, 32'sd0.10578521288564448, 32'sd-0.06835179587760697, 32'sd-0.03274975121794253, 32'sd-0.15423571429995028, 32'sd0.002218736811700651, 32'sd0.01987190427770558, 32'sd0.07041678005145768, 32'sd-0.028235433677435473, 32'sd-0.06669384207615846, 32'sd-0.007407638016839174, 32'sd-0.056507039948130264, 32'sd-0.11937554233024775, 32'sd-0.01604930130843251, 32'sd-0.009619744472537651, 32'sd0.004496782224943858, 32'sd0.07611245934544376, 32'sd0.05560373428578256, 32'sd0.029653909540279598, 32'sd-0.08992981162491266, 32'sd-0.09951921902720764, 32'sd0.009473117335254475, 32'sd0.1279844902305383, 32'sd-0.08361375363639856, 32'sd-0.1086569242976662, 32'sd-0.08292999330394699, 32'sd0.06970751136150317, 32'sd-0.008951084454748409, 32'sd-0.0051457065180525495, 32'sd0.08908610894244044, 32'sd0.04817718266854948, 32'sd-0.0427571815043901, 32'sd0.032323924995940674, 32'sd-0.11187160466856476, 32'sd0.010185945937584429, 32'sd-0.015115351668037822, 32'sd0.027223799032908193, 32'sd-0.02493336404875123, 32'sd0.03244983459540413, 32'sd-0.036814111213774946, 32'sd-0.1656357165735542, 32'sd0.01804340569972603, 32'sd-0.023127769403981698, 32'sd0.10680956700024571, 32'sd0.09718842872349331, 32'sd0.1904896045543564, 32'sd0.097092874843325, 32'sd0.12706636162345275, 32'sd0.1299367228202502, 32'sd0.10896529771845392, 32'sd0.1650812661604044, 32'sd0.005984038900435398, 32'sd-0.026412189364026863, 32'sd-0.021486758320937858, 32'sd0.02705390223203296, 32'sd-0.11780808342693003, 32'sd0.06896693480664276, 32'sd0.019866898637007233, 32'sd-0.08497686986642386, 32'sd-0.041476539927449325, 32'sd-0.12507994126726124, 32'sd0.007303328532756729, 32'sd0.09609932687560457, 32'sd0.052374052696034505, 32'sd-0.012141653317389447, 32'sd-0.008976667628871367, 32'sd-0.023926541264847088, 32'sd0.04110542923528104, 32'sd-0.050074930458348134, 32'sd-0.08151889273284842, 32'sd-0.059397637016226495, 32'sd0.0760251186231477, 32'sd0.03200636699454223, 32'sd0.2200445515194834, 32'sd0.08915620076337782, 32'sd0.12442606972865736, 32'sd0.12129210226050963, 32'sd-0.006768003520582663, 32'sd0.08747889491363132, 32'sd-0.06915058762868356, 32'sd-0.039367344230590295, 32'sd0.10860534713683753, 32'sd0.12459465745049476, 32'sd0.008121752882236618, 32'sd0.04951158142621487, 32'sd0.017359224468303583, 32'sd-0.13862413908319354, 32'sd0.05116093325523968, 32'sd0.003741821476070519, 32'sd0.024910178325482788, 32'sd0.039857298203864064, 32'sd0.09656058113652781, 32'sd-0.012872986338933683, 32'sd0.0623107226345251, 32'sd-0.02390174811509832, 32'sd-0.008236401497793939, 32'sd0.09472886709549774, 32'sd-0.06996009939398529, 32'sd0.06211374536932481, 32'sd0.0666186554333277, 32'sd0.17866328968536954, 32'sd0.12211744249220126, 32'sd0.17828263745030212, 32'sd0.1158587234300048, 32'sd0.14284586367077007, 32'sd0.014531343217497902, 32'sd0.11751941537081682, 32'sd-0.025572776976197555, 32'sd0.006785950713892051, 32'sd0.07515941104198387, 32'sd0.11175993527006373, 32'sd0.17554953119441438, 32'sd0.17705888824246604, 32'sd0.13650012839103098, 32'sd0.023423627993339406, 32'sd0.027085131206968014, 32'sd0.026604292736938828, 32'sd-0.00839396672622936, 32'sd0.025409622646994656, 32'sd0.1412000271598886, 32'sd0.022110865066904503, 32'sd0.09732524895140952, 32'sd-0.02979687128655932, 32'sd-0.03330490109187831, 32'sd0.002305014634661595, 32'sd0.09549276251496955, 32'sd-0.017664854566793873, 32'sd-0.10356186571679951, 32'sd0.021199784421480253, 32'sd0.029513935258357406, 32'sd0.14848802672543812, 32'sd0.01688887022107178, 32'sd-0.010110104245393799, 32'sd0.06889808556591397, 32'sd0.10580353310411716, 32'sd-0.006745055454090973, 32'sd0.06704110894352536, 32'sd0.24855572713688348, 32'sd0.24873948172079957, 32'sd0.17300996591721693, 32'sd0.05344157598960836, 32'sd0.1422041420512886, 32'sd0.10800493250216543, 32'sd0.05600051709128595, 32'sd0.1250171363004398, 32'sd-0.012584217887074714, 32'sd-0.03000664066552564, 32'sd0.06057383226421702, 32'sd0.05140518541955187, 32'sd0.021231980509149137, 32'sd-9.385349569559551e-126, 32'sd-0.02036949934983427, 32'sd0.08807813576006938, 32'sd-0.0005349958323213171, 32'sd0.011689075054693979, 32'sd0.11979375930735905, 32'sd0.025653110432552813, 32'sd0.0038539760337305065, 32'sd-0.0074769432885053375, 32'sd0.047024192740915856, 32'sd0.12755100269482544, 32'sd0.24872300027178854, 32'sd0.12407545217789431, 32'sd0.15875478438710922, 32'sd0.12751392807447445, 32'sd0.2378271970318997, 32'sd0.10759802423846672, 32'sd-0.02944117445346014, 32'sd0.04128514491304113, 32'sd-0.05358735069550673, 32'sd0.14892658026555855, 32'sd0.14708491632832718, 32'sd0.17013198859866396, 32'sd0.021154194872284007, 32'sd-0.07198802869186045, 32'sd0.04806194534426588, 32'sd0.04712061800807052, 32'sd-0.014814464140369767, 32'sd-0.009475418339402504, 32'sd-0.021103434920992214, 32'sd-0.04982429396157402, 32'sd0.1151008210816697, 32'sd0.07471554923086507, 32'sd0.028782130270184513, 32'sd-0.02248319173043363, 32'sd0.04705903946124826, 32'sd0.046836343957569096, 32'sd0.07151224530062399, 32'sd-0.007654992034593955, 32'sd0.19695442069451255, 32'sd0.28469573524746467, 32'sd0.1165123538913789, 32'sd0.06300386048273364, 32'sd0.07826082968238211, 32'sd0.11082421999877168, 32'sd0.0635777125575715, 32'sd-0.0431778746485818, 32'sd0.05805571818040209, 32'sd0.15817649897844607, 32'sd0.17818768521741876, 32'sd0.06007270268961508, 32'sd0.08265166045822572, 32'sd0.05574233080011169, 32'sd0.07047561393631742, 32'sd-0.030749605846220298, 32'sd0.021704838790140502, 32'sd-0.014915609793980052, 32'sd-0.07999272789771322, 32'sd0.006019598964371507, 32'sd0.08936471655069665, 32'sd0.17609348988955492, 32'sd0.04741345075804168, 32'sd0.05614404491239928, 32'sd0.028311076072547316, 32'sd-0.05041661058735072, 32'sd0.014275693317685982, 32'sd0.004305673882246369, 32'sd0.049541298725045264, 32'sd0.15938951952615643, 32'sd-0.009651973039882201, 32'sd0.01205045266091479, 32'sd0.05306299894045264, 32'sd0.12739467731409526, 32'sd0.03986912890905662, 32'sd0.0753274395433932, 32'sd0.04370405239363972, 32'sd0.10938712772965807, 32'sd0.14995328827303, 32'sd0.09267721485725859, 32'sd0.16641449717583778, 32'sd0.15882002392040412, 32'sd0.06761858802775429, 32'sd0.08554129906448418, 32'sd-0.0026447438723746328, 32'sd7.442000441026734e-120, 32'sd0.04488239983015212, 32'sd0.06459451346734199, 32'sd0.07642704764376516, 32'sd0.031126103958976872, 32'sd0.02352910263174459, 32'sd-0.04002675370264625, 32'sd-0.028541027955619518, 32'sd-0.08101265269220408, 32'sd-0.038843724889121786, 32'sd-0.08465003621534663, 32'sd0.01965735626892018, 32'sd-0.013456210328654093, 32'sd0.02610082999592378, 32'sd-0.09636047315152249, 32'sd-0.07349278061216466, 32'sd-0.02283684696379816, 32'sd0.06340196070507577, 32'sd0.029581229267982, 32'sd-0.004180125219415051, 32'sd0.1121425326584697, 32'sd0.1461557432767449, 32'sd0.05905558493586361, 32'sd0.09686798473199015, 32'sd0.07248545036734289, 32'sd0.034680313831183425, 32'sd0.03776538902975128, 32'sd0.01055293534656376, 32'sd0.00874706583102543, 32'sd0.03425955344113774, 32'sd-0.10168119223030812, 32'sd-0.11693935723826818, 32'sd0.06373809334259951, 32'sd-0.013589870837847549, 32'sd-0.0039057731163224373, 32'sd0.02857863297905565, 32'sd0.016593546733719364, 32'sd-0.01676384621805603, 32'sd-0.06632724598999645, 32'sd-0.10750679991700075, 32'sd-0.04363901857985267, 32'sd-0.08597956437230307, 32'sd-0.09492251472181407, 32'sd-0.12202137391331325, 32'sd0.04243002653069355, 32'sd-0.057915704829149296, 32'sd-0.10399387440555691, 32'sd-0.06836233079873338, 32'sd0.026989250384368228, 32'sd-0.0405121603419363, 32'sd0.15413898250151542, 32'sd0.10298528795360247, 32'sd0.07264837628951844, 32'sd0.06998126584516094, 32'sd-0.05953591263189475, 32'sd0.0010194192585629032, 32'sd-0.037217634395523835, 32'sd-0.08391918234433463, 32'sd0.046881335838970195, 32'sd-0.12750423840783107, 32'sd0.03668025174616242, 32'sd-0.08126807375704799, 32'sd-0.009756185261919122, 32'sd0.004075509578560254, 32'sd-0.021104782420428292, 32'sd-0.07804136769453407, 32'sd-0.11160150418489609, 32'sd-0.01606431918958792, 32'sd-0.09299512145925587, 32'sd-0.11482810140113592, 32'sd-0.09216509524279795, 32'sd-0.05309637004844691, 32'sd0.011171756654049042, 32'sd-0.044315922714467104, 32'sd-0.049126742553399085, 32'sd-0.04159935175984354, 32'sd0.058997967406754816, 32'sd-0.07691618763300144, 32'sd0.033962490545365584, 32'sd0.004380898857346151, 32'sd0.08904637771723972, 32'sd-0.029994262725083223, 32'sd0.07570212486089066, 32'sd-0.02284867719323977, 32'sd-6.541109918762312e-118, 32'sd-0.016161897575039566, 32'sd-0.005447673810715371, 32'sd0.10501558703120098, 32'sd0.11922860656612166, 32'sd-0.1446690848203544, 32'sd-0.09820228725760596, 32'sd-0.09822252994095068, 32'sd-0.1611521231482897, 32'sd-0.1858868896491393, 32'sd-0.15456893080666834, 32'sd-0.10586735211414025, 32'sd-0.16096461554822583, 32'sd-0.024942638055408514, 32'sd-0.05146162037349845, 32'sd-0.1421701064892276, 32'sd-0.09339505877739696, 32'sd-0.06279717826386935, 32'sd-0.04762557517427654, 32'sd-0.05696287063015866, 32'sd0.005915638740167596, 32'sd-0.05044364964430971, 32'sd-0.020552616454650355, 32'sd-0.04744755159882381, 32'sd-0.01533291193796267, 32'sd-0.019011852405118636, 32'sd0.0210047807291681, 32'sd-5.860479062037891e-115, 32'sd-1.4712622022238289e-126, 32'sd-7.756031592137034e-124, 32'sd0.004225452518948916, 32'sd0.020790265382714748, 32'sd0.150043289668982, 32'sd0.08219220756845431, 32'sd-0.009289394969713857, 32'sd-0.041577018606283773, 32'sd-0.08980781132998979, 32'sd-0.025402648901288467, 32'sd-0.07189410364938975, 32'sd0.024083986865426812, 32'sd-0.0665811050568391, 32'sd-0.010414518145602385, 32'sd-0.006909418101437301, 32'sd-0.04595849704476767, 32'sd-0.015107295194203028, 32'sd-0.0887008936817814, 32'sd0.02686815927627048, 32'sd0.007873278785543746, 32'sd-0.017640415180661173, 32'sd0.03785476962608727, 32'sd-0.04412416090335139, 32'sd0.06547410656631629, 32'sd-0.048053187183641405, 32'sd0.010694976681407535, 32'sd-0.026475829672015637, 32'sd-2.25391286301784e-118, 32'sd-3.902371549931205e-119, 32'sd-1.8253276883396562e-117, 32'sd0.014790035926718698, 32'sd-0.0237466263163601, 32'sd-0.07639398107902692, 32'sd-0.043653603105825486, 32'sd0.01524692794866728, 32'sd0.015308319241825328, 32'sd-0.01693616411946513, 32'sd0.032312054881033815, 32'sd0.03990069333722838, 32'sd0.03301123942500421, 32'sd-0.060744205279508696, 32'sd-0.11530843260325623, 32'sd-0.036774228662539564, 32'sd-0.06049465928003954, 32'sd0.04011675976929184, 32'sd-0.06653407137494656, 32'sd0.0307585128826292, 32'sd-0.03936341419200208, 32'sd-0.05392836582876066, 32'sd-0.06858229501393591, 32'sd-0.04866672988784245, 32'sd0.08527024369375552, 32'sd-0.02161650662500952, 32'sd-0.0016488154115581275, 32'sd0.05302824981503886, 32'sd1.0844976971422828e-123, 32'sd-1.0580815629015581e-115, 32'sd-2.860269306741146e-118, 32'sd-3.745157446717952e-125, 32'sd-0.01962369143570047, 32'sd0.010796801277421546, 32'sd-0.03536056939509567, 32'sd-0.08307088454841467, 32'sd-0.0695697157357401, 32'sd0.03910875585243824, 32'sd-0.08380481633768883, 32'sd-0.06915438881330845, 32'sd-0.017629475302351122, 32'sd0.007826123257352692, 32'sd-0.04490131878881252, 32'sd-0.014356757193023715, 32'sd0.04654012657964138, 32'sd-0.07293543849811666, 32'sd0.08063868404355268, 32'sd0.032721609900473854, 32'sd0.016960987319668958, 32'sd-0.03554622148756686, 32'sd0.016245940324766086, 32'sd-0.12602443595071558, 32'sd-0.045991063080793856, 32'sd0.00024097838483718654, 32'sd0.022171693695551057, 32'sd1.2375083118502952e-121, 32'sd3.5733035430462046e-114, 32'sd5.896063972571847e-127, 32'sd-2.324548639878692e-120, 32'sd-1.817594256564321e-117, 32'sd5.517777068293862e-124, 32'sd-0.0010515375451273098, 32'sd0.03920781906977539, 32'sd0.07368256425241905, 32'sd0.02111006256687729, 32'sd-0.012596285761632886, 32'sd0.022545712782161897, 32'sd0.0007640652046520837, 32'sd0.061959895422333953, 32'sd-0.049692363135021615, 32'sd0.04639154397214353, 32'sd-0.02858472105933874, 32'sd0.04473604703910531, 32'sd0.010203944209872275, 32'sd0.013417555857908709, 32'sd-0.015642362454383805, 32'sd0.05410121001248414, 32'sd0.07236914228230425, 32'sd0.07102349372092, 32'sd-0.02205454369755428, 32'sd0.008567683443659121, 32'sd-1.312193527370669e-115, 32'sd-1.5040502321935456e-115, 32'sd-6.479794585039244e-124, 32'sd-2.025719864438709e-127},
        '{32'sd2.7604103918684044e-116, 32'sd3.991064281917732e-123, 32'sd6.551264945670975e-127, 32'sd3.6640013454777645e-116, 32'sd-1.4691262384565545e-121, 32'sd1.0725862111596379e-116, 32'sd7.00925945489747e-125, 32'sd1.0354872468537485e-115, 32'sd3.332444089573529e-115, 32'sd2.5112425933471157e-121, 32'sd-3.0910602056418186e-120, 32'sd-8.715419392869727e-123, 32'sd-0.004690549344790203, 32'sd0.019572520568328717, 32'sd0.05457001118160732, 32'sd0.07757308571944967, 32'sd-9.840991988428419e-120, 32'sd8.548436243860593e-117, 32'sd-3.356913859545579e-121, 32'sd-6.036205629776601e-120, 32'sd8.845835235129169e-127, 32'sd7.346681712169826e-117, 32'sd2.0868612157220146e-114, 32'sd9.560007797618902e-119, 32'sd-1.0299374109396178e-124, 32'sd-2.2749081868729616e-127, 32'sd5.27467068854936e-118, 32'sd-1.0279824690810015e-121, 32'sd-2.7246411505209834e-116, 32'sd-2.8602607156862173e-122, 32'sd-3.4830043353132066e-116, 32'sd7.976667365831411e-120, 32'sd-0.01670867115748237, 32'sd-0.029193487313006854, 32'sd-0.08472123930971855, 32'sd0.014975057550348536, 32'sd0.011656914005492326, 32'sd-0.013606150423673927, 32'sd0.002616925122394205, 32'sd0.0407852153195104, 32'sd-0.07748266547218723, 32'sd-0.0020008448680403834, 32'sd0.03113420984717467, 32'sd0.04362172182814591, 32'sd0.03253548476944127, 32'sd-0.07901944286274036, 32'sd0.005175531535389818, 32'sd-0.04245918394534456, 32'sd-0.019270192291068477, 32'sd0.029100225819519047, 32'sd-0.015030534809700383, 32'sd0.06240240796995625, 32'sd3.539728279783314e-125, 32'sd-3.9671920316056483e-119, 32'sd2.715989360514161e-124, 32'sd-5.988252347892566e-126, 32'sd2.0532101992835853e-126, 32'sd-6.03722065819514e-121, 32'sd0.03873189312494699, 32'sd0.04797778726291348, 32'sd0.0317008127808214, 32'sd0.08544491899247196, 32'sd0.031560353924501475, 32'sd0.01152972258693213, 32'sd-0.08204932451015114, 32'sd-0.07016488198161647, 32'sd0.04720954436673524, 32'sd-0.10289917240383414, 32'sd0.023449132012385868, 32'sd0.02487230334221363, 32'sd-0.07536848885101599, 32'sd0.014742821615287933, 32'sd-0.006023505768225852, 32'sd0.07117012566322732, 32'sd0.04180420684889836, 32'sd0.07920864840316456, 32'sd-0.051818855130861055, 32'sd0.05131753025021014, 32'sd-0.03588419682447816, 32'sd-0.06954766901790195, 32'sd0.044414236977196396, 32'sd0.014100256662482524, 32'sd6.468886127322614e-127, 32'sd1.966008462160546e-123, 32'sd6.887930147199955e-127, 32'sd-1.6256356034314838e-126, 32'sd0.03935599496152746, 32'sd-0.05088733698474664, 32'sd-0.01178963946719901, 32'sd-0.0983448592342785, 32'sd0.02928802533587259, 32'sd0.04224790163511154, 32'sd-0.023242333403894862, 32'sd0.007057397587137963, 32'sd0.03415878942889862, 32'sd-0.05374624966371631, 32'sd-0.1517808864731953, 32'sd-0.09285939997647426, 32'sd0.030163233004367712, 32'sd0.02930622288627159, 32'sd0.03374711954604529, 32'sd0.06088078435153755, 32'sd-0.005204359958417482, 32'sd-0.033971991973447004, 32'sd-0.03555214796679199, 32'sd-0.057932291382459956, 32'sd-0.02800283784088793, 32'sd-0.010931158142174878, 32'sd0.04296288134639926, 32'sd0.026020063115082568, 32'sd-0.15846917040458722, 32'sd3.125410495895047e-123, 32'sd-1.1327627487643289e-126, 32'sd0.0011352045265339303, 32'sd0.034695112176854614, 32'sd0.04369501080227438, 32'sd0.10970277845585077, 32'sd-0.010283878237318482, 32'sd-0.04596572995542938, 32'sd-0.08715713143916383, 32'sd-0.008055761064324683, 32'sd0.07520019978388844, 32'sd0.13474514020218584, 32'sd0.001302453811268115, 32'sd0.051389505770765585, 32'sd0.037758487174621894, 32'sd-0.05285199002897382, 32'sd-0.022709452857415713, 32'sd-0.028311762341707583, 32'sd-0.04632068092999656, 32'sd0.012970686191473613, 32'sd0.09390262883194396, 32'sd0.13326531861081792, 32'sd-0.004012118209696566, 32'sd0.1113032741041339, 32'sd0.02581401362205995, 32'sd0.05061523079579428, 32'sd-0.00904289816906405, 32'sd-0.027876836162737978, 32'sd-0.038806411602107765, 32'sd4.738343659642926e-125, 32'sd0.050338061557877414, 32'sd-0.0013953474928140898, 32'sd-0.04799257126563223, 32'sd-0.017431491242370395, 32'sd0.012271304998571576, 32'sd0.08141485340164131, 32'sd0.00337844478457582, 32'sd-0.022933170984525297, 32'sd0.0645636602497568, 32'sd0.09302703122346029, 32'sd0.050011179129730146, 32'sd-0.02337054713175402, 32'sd-0.19441833950303242, 32'sd-0.05617941141656937, 32'sd-0.06193414430469172, 32'sd-0.09777236597816778, 32'sd-0.06709585429741456, 32'sd0.019634691440975776, 32'sd0.08233035992871851, 32'sd0.04577607402221286, 32'sd0.02868470681496019, 32'sd0.15659318893970126, 32'sd0.028869841957427568, 32'sd0.07143627395736475, 32'sd0.12394062609929965, 32'sd0.0076982914081691525, 32'sd0.04316974780688214, 32'sd-3.6422717847352354e-123, 32'sd0.045783435874787066, 32'sd-0.023819501964961524, 32'sd-0.027281039494791742, 32'sd0.026274486163371257, 32'sd0.009663991387352062, 32'sd0.06513331938145522, 32'sd-0.03764711119477878, 32'sd-0.03309857759958823, 32'sd-0.07091011479685118, 32'sd-0.07356445730320911, 32'sd0.008714699403445126, 32'sd0.04366454403466712, 32'sd-0.04922104585555778, 32'sd-0.03547412955054416, 32'sd-0.224148454171237, 32'sd-0.30699053787911995, 32'sd-0.06418085464001456, 32'sd-0.016677152609187233, 32'sd-0.013233184725825723, 32'sd0.024200609411190156, 32'sd-0.035108237555438536, 32'sd0.041516975283921245, 32'sd0.12541747414218055, 32'sd0.1471449185533728, 32'sd-0.06243289430231265, 32'sd-0.02617783854987878, 32'sd-0.006845224109662947, 32'sd0.010633054406226226, 32'sd-0.013491772979362231, 32'sd0.05158296906961183, 32'sd0.017802468411033993, 32'sd0.1853672181795916, 32'sd0.12560490550893316, 32'sd0.05161740201924672, 32'sd-0.03757277974528009, 32'sd-0.14854056448956768, 32'sd0.0768528471021121, 32'sd-0.030535308409567925, 32'sd0.11973096922623283, 32'sd0.19142963500200993, 32'sd0.21692243751996076, 32'sd-0.03505838112665013, 32'sd-0.2526810807393269, 32'sd-0.19862968861542168, 32'sd0.035357445469172966, 32'sd0.13919791882557175, 32'sd0.05643115407627347, 32'sd-0.060132675111838084, 32'sd0.059928296905782795, 32'sd0.06313969408766426, 32'sd0.17206444850588085, 32'sd0.12795396967271938, 32'sd-0.060916433610031066, 32'sd-0.006115930404857743, 32'sd-0.16516452660453512, 32'sd0.023740061701563994, 32'sd-0.0003992251496012768, 32'sd0.0663241685922064, 32'sd0.029987155653324663, 32'sd0.024794641912184393, 32'sd-0.13148557324496124, 32'sd0.02335377515735377, 32'sd0.10267016878705343, 32'sd-0.1170524176462143, 32'sd-0.07764894607325323, 32'sd0.028031278067062484, 32'sd0.009620047810520801, 32'sd0.12319509448488204, 32'sd0.1820952682832238, 32'sd-0.14004335476444688, 32'sd-0.23166869472442428, 32'sd-0.16412925628868835, 32'sd0.017084725465166567, 32'sd0.07901780778640428, 32'sd-0.03878824873183955, 32'sd0.01851452908937528, 32'sd0.07231430211156072, 32'sd-0.015754702514844128, 32'sd-0.03516562421742521, 32'sd0.024880553297392943, 32'sd-0.01802531908290987, 32'sd-0.10795227977212442, 32'sd-0.012114535456125113, 32'sd0.11436050915052218, 32'sd-0.011051927522093042, 32'sd0.03879755050123514, 32'sd0.04464490517954095, 32'sd-0.08716522499225372, 32'sd0.024605389782161237, 32'sd-0.05833882348598383, 32'sd0.0468138240248354, 32'sd-0.08884668328299988, 32'sd-0.010449650500777693, 32'sd-0.041327526843112465, 32'sd0.09373834493981935, 32'sd0.09187079406227679, 32'sd0.015929241775525495, 32'sd-0.04947539422754137, 32'sd-0.3057417984619185, 32'sd-0.2460194090800234, 32'sd-0.057771907334997576, 32'sd0.19380558293943886, 32'sd0.13737803569313692, 32'sd0.079556011213883, 32'sd0.1863417784999145, 32'sd-0.08851346149893499, 32'sd-0.04954596809155648, 32'sd0.028681607642514026, 32'sd-0.08958706429917437, 32'sd0.005167154395788273, 32'sd0.0033010588134041664, 32'sd-0.02114596397654383, 32'sd0.018585437273304143, 32'sd-0.13375418350280502, 32'sd0.027904540502301043, 32'sd-0.020108312093797737, 32'sd-0.018024769123775698, 32'sd0.0004383099550093595, 32'sd-0.03708046110839354, 32'sd-0.08485963099924258, 32'sd-0.011375361204175708, 32'sd-0.000738608695432344, 32'sd0.10463707507377897, 32'sd0.12895341700467064, 32'sd0.012362881345245725, 32'sd-0.2696415690317154, 32'sd-0.45057726304440515, 32'sd-0.1917224068944652, 32'sd0.0895174772382873, 32'sd0.1433135676976798, 32'sd0.07622388550009412, 32'sd-0.02508166901402488, 32'sd0.10006675395267974, 32'sd-0.014072316850306564, 32'sd0.024108699689980098, 32'sd0.01543211261161444, 32'sd-0.05765048542907405, 32'sd-0.09481535779510046, 32'sd-0.1094058665007115, 32'sd0.015939647371116666, 32'sd-0.007334852184193388, 32'sd-0.0390254758638069, 32'sd-0.015502863600767958, 32'sd0.036006342141931415, 32'sd0.011695081537778632, 32'sd-0.017713517052306286, 32'sd0.053398376228304234, 32'sd-0.018673880388969152, 32'sd-0.023661720870969502, 32'sd0.03286941459862412, 32'sd-0.030229545727911974, 32'sd0.07139573098787284, 32'sd-0.10209718391734657, 32'sd-0.227890762539877, 32'sd-0.4027579617347347, 32'sd-0.055763853782269175, 32'sd0.12987980321201167, 32'sd0.12891841137812712, 32'sd0.06427589765565483, 32'sd0.0539036583853566, 32'sd0.052143531292965124, 32'sd0.021038023907263104, 32'sd-0.10072940162789328, 32'sd-0.03988337193002216, 32'sd-0.13633867336309502, 32'sd0.014707362548538393, 32'sd0.01670328812974445, 32'sd0.030159795062223375, 32'sd0.0015427787589028968, 32'sd-0.01898995226665387, 32'sd-0.0017888335655764061, 32'sd-0.07225080454585009, 32'sd-0.05125495653099162, 32'sd-0.04460941929448356, 32'sd-0.09857781845428672, 32'sd-0.018017461629144988, 32'sd0.08858252061862867, 32'sd-0.0009009561931614122, 32'sd0.01373262897446112, 32'sd0.04542202960835377, 32'sd-0.014049681425239192, 32'sd-0.1296485106163065, 32'sd-0.29150706834131024, 32'sd-0.02925857987055191, 32'sd0.14021716830456835, 32'sd0.028170235793321792, 32'sd0.03933903225883354, 32'sd0.021711732891890947, 32'sd0.07370889058192105, 32'sd0.15223410426593442, 32'sd-0.11611193437129362, 32'sd-0.004907425678055212, 32'sd0.015972373844973988, 32'sd0.034088519559273806, 32'sd-0.04700483169181956, 32'sd-0.0034269424837733847, 32'sd0.028837539196788903, 32'sd-0.07226326080445945, 32'sd-0.03335608380400932, 32'sd0.05598231163033635, 32'sd-0.025155151464462365, 32'sd0.01392380083502094, 32'sd-0.04736996741827843, 32'sd0.030512491183862837, 32'sd0.1440065592586242, 32'sd-0.028053455299628584, 32'sd0.09231129447454231, 32'sd0.08101217301407222, 32'sd-0.1182981275450529, 32'sd-0.18323643414976862, 32'sd-0.19698031968814125, 32'sd0.034380719381519306, 32'sd0.1465583954284121, 32'sd0.10997595643268317, 32'sd0.08479452153208841, 32'sd-0.034651648280051635, 32'sd0.1261205863503332, 32'sd0.04094487066385231, 32'sd-0.014222095438139747, 32'sd-0.023850671243596452, 32'sd-0.13376283182896923, 32'sd-0.03501784631488758, 32'sd0.07281518346905133, 32'sd-0.0018074079215998173, 32'sd0.02659042447008962, 32'sd-0.012361287665666432, 32'sd-0.05187388915933712, 32'sd-0.05494942718027587, 32'sd0.05127777763925935, 32'sd-0.00039641305765135556, 32'sd0.14812168238631662, 32'sd0.03367825187787112, 32'sd0.10210321097949202, 32'sd0.03273890256859964, 32'sd0.027271572469970744, 32'sd0.007522945540601436, 32'sd-0.14080613234589828, 32'sd-0.12069023572772411, 32'sd-0.2007799936026945, 32'sd-0.0005146135675505574, 32'sd0.17205886027281778, 32'sd-0.0873653846381319, 32'sd0.03734949453497092, 32'sd-0.009436706112584313, 32'sd0.12286413798464611, 32'sd-0.007692945151476341, 32'sd-0.02367143639569565, 32'sd0.00859677714891652, 32'sd0.04119267297203028, 32'sd-0.12388363369976299, 32'sd0.06169128952944574, 32'sd-0.015401963758779025, 32'sd0.1393793574918949, 32'sd0.11754192168428818, 32'sd-0.0549244809740607, 32'sd0.018188423073636162, 32'sd-0.05771753289280716, 32'sd-0.042544727952156136, 32'sd0.16185357716251647, 32'sd0.09539671861130795, 32'sd0.0021667671337464163, 32'sd0.030495925514182846, 32'sd0.12706449920374066, 32'sd0.0872619642823265, 32'sd-0.07483905048639325, 32'sd-0.039488308196107665, 32'sd-0.03950912473321824, 32'sd0.04778966527499725, 32'sd0.1010198325588613, 32'sd-0.018459015927790354, 32'sd0.04043612345511026, 32'sd-0.018378638014229415, 32'sd-0.12255815704758487, 32'sd-0.003568589846697168, 32'sd-0.11824222661978175, 32'sd0.030035311328028544, 32'sd0.04486479361154082, 32'sd-0.01534560630325365, 32'sd0.0616966085635834, 32'sd0.048437955468127195, 32'sd-0.023441775161209898, 32'sd0.028223239819167103, 32'sd0.033754246426092434, 32'sd0.04905940169013584, 32'sd-0.09693474231816712, 32'sd0.026430023033693704, 32'sd-0.041667291601671416, 32'sd-0.00637005521261496, 32'sd-0.03352364235774693, 32'sd-0.021820790925706768, 32'sd-0.10086384494542162, 32'sd-0.07495072640306705, 32'sd-0.005164509929802598, 32'sd-0.009016063564008149, 32'sd0.024859068869499498, 32'sd-0.06423032184149918, 32'sd0.052807339669284865, 32'sd0.008455035089727975, 32'sd-0.012662428368938232, 32'sd-0.08246277983777266, 32'sd-0.03888110400922639, 32'sd-0.03256255820872247, 32'sd-0.13370018548274842, 32'sd-0.07318746174442642, 32'sd-0.004310595602662091, 32'sd-0.011628912267128096, 32'sd-0.015761063133260967, 32'sd-2.6308446330589834e-114, 32'sd-0.023176578359078433, 32'sd-0.04462443020022007, 32'sd0.047721718452694364, 32'sd0.10460830727815724, 32'sd-0.03760432127076465, 32'sd0.0044329193488078095, 32'sd0.01897333317123289, 32'sd0.03847257890791026, 32'sd-0.09001882785604533, 32'sd-0.0504007917744555, 32'sd0.006278584914829292, 32'sd0.04038205570084362, 32'sd0.19130015436263387, 32'sd-0.022427460294389027, 32'sd0.017527106970848205, 32'sd-0.03463543144805029, 32'sd0.07764929145177284, 32'sd0.0077592277334183135, 32'sd0.09126134314662648, 32'sd-0.03453033468119889, 32'sd-0.011510889028521492, 32'sd0.08560636026765313, 32'sd-0.03928794104859989, 32'sd-0.16986316506991322, 32'sd0.04851570143278727, 32'sd0.018662839795818134, 32'sd0.016943733314837946, 32'sd-0.01105357946436385, 32'sd-0.039123646150564004, 32'sd-0.07182322520538197, 32'sd0.02114722522703916, 32'sd-0.006632480586689822, 32'sd0.008128224653614012, 32'sd-0.014707893558652561, 32'sd0.025039490300033055, 32'sd-0.01852350859470428, 32'sd0.07088127525871205, 32'sd0.004390840492756595, 32'sd0.0020430590243422733, 32'sd0.13129855922544206, 32'sd0.04398576528102205, 32'sd0.07049198082397296, 32'sd-0.013703395068646885, 32'sd0.04019910934843802, 32'sd-0.02116646476754495, 32'sd0.053641406390904534, 32'sd0.09013282730949451, 32'sd0.0020108635508298794, 32'sd-0.03183440478107291, 32'sd-0.07577875541207771, 32'sd-0.10424266308762019, 32'sd-0.048138803655473746, 32'sd-0.006429174386933481, 32'sd0.08251851228421439, 32'sd0.05095349226519012, 32'sd0.02077387648547296, 32'sd0.032061701019393464, 32'sd0.011917750287222735, 32'sd0.00435017084432544, 32'sd0.021479110177144645, 32'sd0.02151820845983356, 32'sd-0.05972088082480302, 32'sd0.013312303450704183, 32'sd0.048388236022341116, 32'sd-0.0007071754671515942, 32'sd-0.037563136370358984, 32'sd0.01464503948891033, 32'sd0.0871935483265059, 32'sd0.05175325037745046, 32'sd0.0038438889019962075, 32'sd0.0342320052414681, 32'sd0.031128092536612317, 32'sd0.022785818303047805, 32'sd0.04828180878936564, 32'sd-0.04098053831643844, 32'sd0.0032244996281722478, 32'sd0.1379758152017521, 32'sd0.014626020626357396, 32'sd0.015196407466950548, 32'sd0.022566408435147855, 32'sd0.010895675906200889, 32'sd0.0016027975373004177, 32'sd0.12538503402830747, 32'sd8.485842474443568e-122, 32'sd0.028170570742661914, 32'sd-0.032364360688034256, 32'sd-0.07297150207632777, 32'sd-0.10367574241416448, 32'sd0.01094954996207686, 32'sd-0.011884809321432929, 32'sd0.011064100733050905, 32'sd-0.0819214114590567, 32'sd-0.038815821303185616, 32'sd0.022540514812856, 32'sd0.10627300820196652, 32'sd0.01669967371487459, 32'sd0.08914984499379715, 32'sd0.014053178765543035, 32'sd-0.0732594694964056, 32'sd0.11331037464375109, 32'sd0.037691101022115, 32'sd0.032772509653099954, 32'sd0.13220376860794614, 32'sd0.015285183864204127, 32'sd0.13279080727424908, 32'sd0.08789103169889222, 32'sd0.053064209060156665, 32'sd-0.05792419667045586, 32'sd-0.013055589411641304, 32'sd-0.023344809488049352, 32'sd-0.023178383681063265, 32'sd-0.020185697637252985, 32'sd-0.007574158324102241, 32'sd0.08868387162611055, 32'sd-0.001894178533011763, 32'sd-0.12552010943910197, 32'sd-0.025044451253550967, 32'sd-0.031108532840963724, 32'sd-0.04999230333476879, 32'sd-0.018353800162944547, 32'sd-0.03506640304603434, 32'sd-0.032021907742721394, 32'sd0.0686902923403117, 32'sd0.03180636883442473, 32'sd0.054138069009663815, 32'sd-0.07304628937084588, 32'sd-0.06829882598214443, 32'sd0.03428237211496884, 32'sd0.038991182605814856, 32'sd0.036644457528569555, 32'sd0.0836287532508967, 32'sd0.12536141664041855, 32'sd-0.08205673637393512, 32'sd-0.03011086726827662, 32'sd0.0284752971552018, 32'sd0.02605365637648222, 32'sd-0.05610209203864915, 32'sd-0.013749289149312864, 32'sd0.08182971555670708, 32'sd0.019108716335752292, 32'sd0.07451207475979733, 32'sd-0.0049639640047733375, 32'sd0.06874235345864091, 32'sd-0.0031198033190232544, 32'sd-0.0430361301378147, 32'sd-0.0021965467388703297, 32'sd-0.04355859255417674, 32'sd0.002818091860713866, 32'sd-0.08905692005202541, 32'sd-0.09356914612516923, 32'sd0.04107121018979666, 32'sd0.1124678656023374, 32'sd0.011831757247319153, 32'sd0.012436367448382663, 32'sd-0.0444893973449762, 32'sd0.03825199983091002, 32'sd-0.11052088047750874, 32'sd-0.11230209217273589, 32'sd0.05371714506483527, 32'sd0.08740274303063017, 32'sd0.10462587585491831, 32'sd-0.032275718906436345, 32'sd0.1172332208220609, 32'sd0.09164578336541472, 32'sd0.022321059239538994, 32'sd0.05773369354623826, 32'sd0.02785263435896592, 32'sd-4.1046663250256626e-120, 32'sd-0.0012635693711811383, 32'sd-0.04330633781045698, 32'sd-0.007134016577458461, 32'sd-0.02418931967420342, 32'sd-0.14042799827313898, 32'sd0.010462906641421356, 32'sd0.11194261851731385, 32'sd-0.000102992236630512, 32'sd-0.047687390597655005, 32'sd-0.041046000765090455, 32'sd0.08098665954351245, 32'sd0.09173548960435737, 32'sd0.060269384545643255, 32'sd0.05351418690221116, 32'sd0.07101619811382459, 32'sd0.05338984038761699, 32'sd-0.06297078470724318, 32'sd-0.12890836550844376, 32'sd-0.13460422576777759, 32'sd-0.0014833577660468347, 32'sd-0.0169233847755794, 32'sd-0.010593581851129729, 32'sd0.06042434684251901, 32'sd0.112051274627668, 32'sd0.07898581711241034, 32'sd-0.03900836493126912, 32'sd-2.12857700283652e-124, 32'sd-2.7670525976957805e-114, 32'sd-7.759354772406389e-117, 32'sd-0.006992539859317579, 32'sd-1.1953124139250761e-05, 32'sd-0.05465961416650539, 32'sd-0.0315178306736076, 32'sd-0.058532842847934356, 32'sd0.06220463762238276, 32'sd0.07974062969025832, 32'sd-0.053288993430414405, 32'sd-0.010271945013900547, 32'sd0.049071274743326385, 32'sd0.16565166338629506, 32'sd0.05607221288743807, 32'sd0.08841479302126108, 32'sd-0.033636818702808345, 32'sd0.10554587931024116, 32'sd-0.07045037690744414, 32'sd-0.11633900303708236, 32'sd-0.0737875487604125, 32'sd-0.0743534307056024, 32'sd-0.053998930903784145, 32'sd0.02936838287874721, 32'sd-0.02646085635073382, 32'sd0.028719854796235164, 32'sd0.007272976022986162, 32'sd-0.022538674742549666, 32'sd9.105650827647206e-125, 32'sd3.62755732418259e-122, 32'sd-2.4161650625567848e-114, 32'sd-0.024005561082109276, 32'sd-0.04026283326211619, 32'sd0.004961755698754259, 32'sd-0.11254438517943897, 32'sd0.1315848335022591, 32'sd-0.044407500900844034, 32'sd0.02814286735645689, 32'sd-0.03611624622340477, 32'sd0.07929606188441271, 32'sd0.0015541033097133093, 32'sd0.08065116015384934, 32'sd-0.10076998837922599, 32'sd-0.0010270632200207015, 32'sd0.00217348779190653, 32'sd0.05119617727644804, 32'sd-0.04666312592197582, 32'sd-0.09332741217768038, 32'sd-0.011401843984403144, 32'sd-0.018895699420345965, 32'sd-0.047755564841948775, 32'sd-0.0221351166862154, 32'sd0.05987379387199164, 32'sd-0.11579986488653228, 32'sd0.033529426419638665, 32'sd0.08573009604514595, 32'sd9.494236965128082e-126, 32'sd-2.969827903223168e-121, 32'sd2.4047618282346158e-116, 32'sd-1.1857485455174213e-126, 32'sd0.03809326891690466, 32'sd-0.019801124682013893, 32'sd-0.07102131652960028, 32'sd-0.015704263934448816, 32'sd-0.05977202458874218, 32'sd0.018678382040435437, 32'sd-0.08371855599203494, 32'sd-0.08724778435254209, 32'sd-0.07428661402637714, 32'sd-0.059613642455900596, 32'sd0.008297868439603041, 32'sd-0.09331003432706497, 32'sd0.03997966404076983, 32'sd-0.08125511795524355, 32'sd0.06955185118487145, 32'sd0.05480679426806934, 32'sd-0.11590344633478362, 32'sd-0.09148387920580003, 32'sd-0.028356628416486344, 32'sd0.03797843063111681, 32'sd0.007459511470504579, 32'sd0.09414029267481279, 32'sd0.04730179989282916, 32'sd2.4263064781705124e-120, 32'sd3.8592787099528734e-120, 32'sd-8.2607412179027e-121, 32'sd8.841529729617866e-119, 32'sd1.1683956464508045e-117, 32'sd-3.882981995191178e-116, 32'sd0.021433368362029193, 32'sd0.040845379267463296, 32'sd0.02450956630235675, 32'sd0.03906575250533854, 32'sd-0.06805287061221911, 32'sd0.06020126049798806, 32'sd0.01718132778255911, 32'sd0.013774638181616252, 32'sd-0.013366907239838183, 32'sd0.02065145027515521, 32'sd0.009378719778949109, 32'sd-0.031186547022657832, 32'sd-0.10318419871318983, 32'sd-0.0166961882621348, 32'sd0.013914267083397104, 32'sd0.05232959321938282, 32'sd-0.02372987586746414, 32'sd0.05152541620886105, 32'sd-0.057995824763349815, 32'sd0.013545979402362913, 32'sd4.853889657518533e-123, 32'sd-1.81737641107417e-120, 32'sd-6.633537712988243e-122, 32'sd-2.1702950752958647e-121},
        '{32'sd1.7937832525550188e-123, 32'sd1.7607808963440817e-117, 32'sd1.2650380859092057e-119, 32'sd-4.617324578611032e-120, 32'sd5.736331483041447e-121, 32'sd2.104689265954844e-117, 32'sd-6.360483338232933e-120, 32'sd-2.03399900877873e-123, 32'sd-9.894766077661026e-122, 32'sd-3.0090273086470426e-125, 32'sd-9.53844120142783e-124, 32'sd-3.663992501385753e-116, 32'sd-0.024574886777604107, 32'sd-0.05040130265795263, 32'sd-0.03118729631783589, 32'sd-0.004817814680072434, 32'sd-3.677817066817497e-116, 32'sd-1.5951075323989315e-119, 32'sd-7.203446615983731e-119, 32'sd4.3319895994836605e-119, 32'sd-1.6814197260029726e-123, 32'sd2.835733198379295e-125, 32'sd-5.107426330302359e-126, 32'sd3.6627443835903634e-122, 32'sd8.777224628690707e-120, 32'sd-3.106809629753331e-125, 32'sd-1.1359636882401965e-119, 32'sd1.6308206887891688e-115, 32'sd-6.745537617397135e-126, 32'sd6.445268556581211e-127, 32'sd6.835598614305548e-124, 32'sd1.2109600075583842e-124, 32'sd-0.07674201785229941, 32'sd-0.083709649024501, 32'sd-0.0470140737666392, 32'sd0.03252906644436456, 32'sd0.01979006606706713, 32'sd-0.007215418475521896, 32'sd-0.033423851869028014, 32'sd-0.024632502849910847, 32'sd-0.10338085682049804, 32'sd0.0265117857279413, 32'sd-0.018899449206695985, 32'sd-0.14091486319390462, 32'sd-0.07097390658211702, 32'sd0.10326847737754791, 32'sd0.10221896218601917, 32'sd0.06364033000618038, 32'sd0.02900092080460337, 32'sd-0.03849213270950506, 32'sd-0.08347259786461718, 32'sd-0.009703563883010753, 32'sd-3.804627440632947e-119, 32'sd-1.6791198883849158e-116, 32'sd4.75810942597572e-124, 32'sd-1.0285630420515787e-120, 32'sd9.050794247774749e-125, 32'sd-4.147611528945907e-126, 32'sd-0.06742082386457983, 32'sd-0.027358448360638412, 32'sd0.06166073561090444, 32'sd-0.026882896128928746, 32'sd0.05537267044994496, 32'sd0.0067216379288874955, 32'sd0.021079851037701644, 32'sd0.07452793942637746, 32'sd0.042487526451254795, 32'sd-0.12997073877107898, 32'sd-0.011898163654947941, 32'sd0.04658044864514535, 32'sd-0.12035981465237026, 32'sd-0.007845273742200313, 32'sd-0.026565893022068365, 32'sd-0.07616365227919572, 32'sd0.0023116539073484714, 32'sd0.017654192905333956, 32'sd-0.006490326154703772, 32'sd0.02271155076085114, 32'sd0.07019925211499167, 32'sd0.07110379477014768, 32'sd-0.060134005010521824, 32'sd-0.07037286075010726, 32'sd9.813648984029276e-121, 32'sd2.5347881841510693e-118, 32'sd6.405925308435033e-122, 32'sd-3.8447981579056066e-123, 32'sd-0.07713908774866615, 32'sd-0.04825476852079323, 32'sd0.08738073325982303, 32'sd-0.04051007548781684, 32'sd0.010855426411468793, 32'sd0.06126965155310798, 32'sd-0.0772658208487311, 32'sd0.009322120158636957, 32'sd0.07117928429379941, 32'sd-0.020892283054893906, 32'sd-0.046090056275233604, 32'sd0.07470165709661486, 32'sd0.00025193121273246646, 32'sd-0.03659924340629733, 32'sd0.001106561347709039, 32'sd-0.007563944743309427, 32'sd0.13430123617513146, 32'sd0.027288752310471953, 32'sd-0.12807333870312615, 32'sd0.09972052838537902, 32'sd0.047785430386741545, 32'sd-0.033910269959691756, 32'sd-0.05570799960663669, 32'sd-0.03598734469411976, 32'sd-0.05128068911403847, 32'sd2.413178849917287e-126, 32'sd-3.631611093713778e-116, 32'sd-0.036889985800327894, 32'sd-0.058009461448656874, 32'sd-0.07854933131989911, 32'sd0.03854140845893546, 32'sd-0.08808343676073137, 32'sd0.03390170764432448, 32'sd0.06318533275490575, 32'sd-0.06953941807260954, 32'sd-0.04411678953185375, 32'sd-0.059792614623067834, 32'sd-0.06428697512777522, 32'sd0.05483138896066703, 32'sd0.013012624539249043, 32'sd0.048290176027651725, 32'sd0.10986296574138542, 32'sd-0.023822953241324503, 32'sd-0.07822545994281199, 32'sd0.0837680014441148, 32'sd0.06918078092607345, 32'sd0.07075461218480424, 32'sd0.11108845491458776, 32'sd-0.031055037193781186, 32'sd-0.08726561329809022, 32'sd-0.14429271451588066, 32'sd-0.062420644547765095, 32'sd-0.00428495386881889, 32'sd-0.047734162000930204, 32'sd-1.6119921662427589e-115, 32'sd-0.05201753111190538, 32'sd-0.0605604199006108, 32'sd0.004346207324023904, 32'sd0.0448804059296093, 32'sd-0.023957559267913466, 32'sd-0.00437996413240291, 32'sd0.005619590472203197, 32'sd0.005354581634281398, 32'sd0.0037197681300687835, 32'sd0.0032301696246155682, 32'sd0.04286116970522855, 32'sd-0.043684463759350416, 32'sd0.15259551765121043, 32'sd0.08146321365993707, 32'sd0.11736314252272002, 32'sd0.01735650720860058, 32'sd-0.009686769169881359, 32'sd-0.029599597725573745, 32'sd0.08667683960502914, 32'sd0.07775556310917034, 32'sd0.010431415237809867, 32'sd-0.0463144510136923, 32'sd-0.15520865813440612, 32'sd-0.07752250593472478, 32'sd-0.09292715236929497, 32'sd-0.026879474674008683, 32'sd-0.08729213630048266, 32'sd1.1646218778421347e-126, 32'sd0.05431948334880265, 32'sd-0.051339341722200595, 32'sd-0.023951316836175407, 32'sd0.0045781147409687944, 32'sd-0.05608109344598525, 32'sd-0.09809755010333567, 32'sd0.09241399407802325, 32'sd0.034607507543774625, 32'sd-0.0830173638656609, 32'sd-0.04572382337338536, 32'sd-0.01719563619321074, 32'sd-0.06275465880861768, 32'sd-0.02940662884091875, 32'sd-0.004895285554622919, 32'sd-0.045041283986871856, 32'sd0.008695745109874139, 32'sd0.03853730947188689, 32'sd0.10423128453803004, 32'sd0.07037170297571062, 32'sd0.07886293107266265, 32'sd-0.02940215535984124, 32'sd0.09284211294530759, 32'sd-0.02331310539222161, 32'sd-0.02745449729655767, 32'sd-0.0030144426501038327, 32'sd-0.0076571996074637156, 32'sd0.006718123536010567, 32'sd-0.033545384984684, 32'sd-0.05604562233012897, 32'sd-0.019721658914485022, 32'sd-0.06259256750741271, 32'sd0.059660521066018275, 32'sd-0.08979044276753767, 32'sd-0.09152340370837767, 32'sd-0.17299214292560153, 32'sd0.014813661759133123, 32'sd-0.021485498566787945, 32'sd-0.0427635125176746, 32'sd-0.049289017919133704, 32'sd-0.14886834167827634, 32'sd-0.13911425637603664, 32'sd-0.09582100736281565, 32'sd0.06372387841213842, 32'sd0.0024765022854416016, 32'sd0.1425798403990677, 32'sd0.12591095683722445, 32'sd0.028752330493134175, 32'sd0.07280846709624807, 32'sd0.01064988498124976, 32'sd0.07819151001995957, 32'sd-0.00839075339243223, 32'sd-0.09735295048773888, 32'sd0.005558815112768533, 32'sd-0.03262773499605717, 32'sd-0.030755016160487213, 32'sd0.08389243213812453, 32'sd-0.09679849311469574, 32'sd-0.07791731348370773, 32'sd-0.04658454055554871, 32'sd-0.032348826056314076, 32'sd-0.12553821083121314, 32'sd0.007187851731022351, 32'sd-0.06430688618738722, 32'sd-0.062128213065583755, 32'sd-0.10519652921726914, 32'sd-0.04270483232593188, 32'sd0.08042391506465667, 32'sd0.026884088876371275, 32'sd-0.016381463219370427, 32'sd0.07327512172973841, 32'sd-0.05495376306528663, 32'sd0.06758637749272353, 32'sd0.12381198703919946, 32'sd0.04865605084686392, 32'sd0.12801113948369267, 32'sd0.0777251778374697, 32'sd0.008441896027153466, 32'sd-0.02426568984567757, 32'sd0.06463711398343822, 32'sd0.03805862885822396, 32'sd0.05970369435694634, 32'sd0.018998740302625657, 32'sd0.02367896989198951, 32'sd-0.00028295594419477336, 32'sd-0.030095934924752116, 32'sd0.045818092218938664, 32'sd0.015148415861012746, 32'sd-0.04031802340641031, 32'sd-0.1363174191701158, 32'sd-0.062451711247774516, 32'sd-0.031182197370813153, 32'sd-0.09533344087436271, 32'sd-0.04561360924022387, 32'sd0.028236511706281903, 32'sd0.16600598057372792, 32'sd0.11349970367746576, 32'sd0.14970219207664434, 32'sd0.10825465520098916, 32'sd-0.01021180930852919, 32'sd-0.13111452856234476, 32'sd-0.10695423805125391, 32'sd-0.16281953615202602, 32'sd0.018607903379575054, 32'sd0.12879492512905844, 32'sd0.11313168910329412, 32'sd-0.03225275843401337, 32'sd0.017926828651660412, 32'sd0.03286913807949443, 32'sd0.12620400898079598, 32'sd0.053922162435454335, 32'sd-0.09456826013795729, 32'sd0.010324847979633227, 32'sd0.0017944090620902456, 32'sd0.006777935602757702, 32'sd-0.049759884225309546, 32'sd0.024319436771702826, 32'sd-0.035600569892108073, 32'sd-0.08205590133810985, 32'sd-0.11774551442252915, 32'sd-0.12631684699642287, 32'sd0.12420696895670975, 32'sd0.1229188900949635, 32'sd-0.02870742251422915, 32'sd0.007603078508743056, 32'sd0.16613849119292645, 32'sd0.15959996473707122, 32'sd-0.025797248581231655, 32'sd-0.03238348520955561, 32'sd-0.011897498647115756, 32'sd-0.009933701636850107, 32'sd-0.04861833549622203, 32'sd0.08199279999265574, 32'sd0.024205049058516698, 32'sd0.043094993411265665, 32'sd0.00135342603738153, 32'sd0.060538747349050126, 32'sd0.053746587593459454, 32'sd0.056657327030239624, 32'sd-0.02955904462700175, 32'sd0.044763405719249985, 32'sd0.024179910311835365, 32'sd0.08991571856264904, 32'sd-0.008479548799147736, 32'sd-0.030241729065571793, 32'sd0.011410431490672992, 32'sd-0.007938633459911313, 32'sd0.09462102471847435, 32'sd0.01846342549383302, 32'sd0.05350026523733001, 32'sd0.1448618404963379, 32'sd0.11907815840434557, 32'sd0.06397934080670527, 32'sd0.09310528686906931, 32'sd0.15956540235245562, 32'sd0.0659644463426044, 32'sd0.07812641712969146, 32'sd-0.043907690787763756, 32'sd-0.13920536909090522, 32'sd-0.041314015420710636, 32'sd0.08557221515934664, 32'sd0.1749574165148764, 32'sd0.08268907184910984, 32'sd0.06758049885830877, 32'sd0.0006921600470375717, 32'sd0.0910521143665151, 32'sd-0.06384015656630605, 32'sd-0.07532754917245328, 32'sd0.010886315423032537, 32'sd-0.08498332727277405, 32'sd-0.06305318260033797, 32'sd0.005982220344164997, 32'sd0.006790893917638737, 32'sd-0.06719264782413494, 32'sd0.07556467261261463, 32'sd0.08124919045759657, 32'sd0.03528365472157137, 32'sd0.14157092835406454, 32'sd0.08551453559830914, 32'sd0.10009682399059766, 32'sd0.05170653661902051, 32'sd0.2206804467003461, 32'sd0.1103672959591857, 32'sd0.0692978108671421, 32'sd0.12078131867544604, 32'sd0.0716258210626226, 32'sd0.0005947450640909563, 32'sd0.0405918426974476, 32'sd0.038069555366090094, 32'sd0.06675016430688759, 32'sd0.01489252660163982, 32'sd0.10347688126715135, 32'sd-0.04673653695811063, 32'sd0.01029004229085705, 32'sd-0.010332112908717196, 32'sd0.03974896658884224, 32'sd0.05160446134875102, 32'sd-0.08890428265042094, 32'sd-0.11083594911463876, 32'sd-0.045784282888748896, 32'sd-0.1640122305972848, 32'sd-0.016134437511518156, 32'sd0.06215046245021288, 32'sd0.10430831209288528, 32'sd0.050815498761916544, 32'sd0.1326955343654945, 32'sd-0.021387353274014982, 32'sd0.07752703813808175, 32'sd0.07507545369130092, 32'sd0.10142290421338204, 32'sd0.059206642561893785, 32'sd0.07364033305897756, 32'sd0.14618113163369628, 32'sd0.03724182535954925, 32'sd0.03024968542009406, 32'sd-0.04223351482153481, 32'sd-0.024768285386456736, 32'sd-0.026922089551257102, 32'sd-0.02104095432984336, 32'sd-0.06776781640019248, 32'sd-0.0572941375763308, 32'sd0.06251284352012165, 32'sd-0.05711420711564224, 32'sd-0.027816558907499657, 32'sd-0.059288887852652225, 32'sd-0.08109115240119873, 32'sd-0.055440215255882955, 32'sd0.0379234969526629, 32'sd0.01858253817915656, 32'sd-0.010355303682371824, 32'sd-0.03126388519636588, 32'sd0.09418910796889599, 32'sd0.13355118374513403, 32'sd-0.01656526396696306, 32'sd0.04721798007205885, 32'sd0.08684575845278195, 32'sd0.03751762605913042, 32'sd0.05365083005029169, 32'sd0.00374104913271637, 32'sd0.029544923284075205, 32'sd0.03919113156686277, 32'sd0.11757535117328914, 32'sd0.03164673341518106, 32'sd-0.09361774950681304, 32'sd-0.11814907252636442, 32'sd-0.05319229371915907, 32'sd-0.031268738854951905, 32'sd0.016923012561311773, 32'sd-0.12292635494345597, 32'sd-0.07046386128650697, 32'sd0.04134874688717489, 32'sd0.007749551788919699, 32'sd-0.0840139584705146, 32'sd-0.05369112718728957, 32'sd-0.07140110512088704, 32'sd-0.05101018641752919, 32'sd0.013889656596956727, 32'sd0.022968044596012798, 32'sd-0.0035828962683217814, 32'sd0.12961423539777434, 32'sd0.02456089620584289, 32'sd0.11119739950057769, 32'sd-0.03170236075449356, 32'sd0.08048582192230558, 32'sd0.12927902500641364, 32'sd0.07307606513851306, 32'sd-0.06049738250294121, 32'sd-0.06869142681106878, 32'sd-0.029776213047825576, 32'sd-0.04132058071648517, 32'sd-0.1078818089729023, 32'sd-0.08222390943734986, 32'sd-0.10682108818285298, 32'sd-0.03182041286095892, 32'sd-0.06922643112108817, 32'sd0.004368067799060373, 32'sd-0.08399669076216262, 32'sd-0.03447056794673023, 32'sd-0.02720957327947438, 32'sd-0.0029796380843794923, 32'sd0.053898973968680625, 32'sd-0.0934470373497868, 32'sd-0.01977964092202378, 32'sd-0.1338547306621466, 32'sd-0.15351943038933707, 32'sd0.017162251565218913, 32'sd0.02801135305541403, 32'sd0.16268139101210816, 32'sd0.1592345907918448, 32'sd0.21402125239397368, 32'sd0.19388962558257075, 32'sd0.142966340679494, 32'sd0.0341517077430397, 32'sd-0.0709118138903978, 32'sd-0.24814140093941778, 32'sd-0.17883561134651174, 32'sd-0.11958556575471516, 32'sd-0.04320345443281973, 32'sd-0.1834568572236694, 32'sd-0.08575030398867917, 32'sd-0.04923966906404076, 32'sd-0.05937186298764445, 32'sd0.01726940275351931, 32'sd-0.020464707772943812, 32'sd0.006350125373239087, 32'sd-0.03415748937849107, 32'sd-0.052052485823789886, 32'sd-0.037242446771820495, 32'sd1.732435704979729e-125, 32'sd0.047280665400710103, 32'sd-0.014880571531857782, 32'sd-0.15245281274539388, 32'sd-0.020998448745801198, 32'sd-0.06466343932813562, 32'sd-0.01615845582368678, 32'sd0.12229772350360542, 32'sd0.12057130991214751, 32'sd0.16865612342183825, 32'sd0.2966723794604098, 32'sd0.03291625679406171, 32'sd-0.08457050993493526, 32'sd-0.27943623960130076, 32'sd-0.22729368117716292, 32'sd-0.1619125603151277, 32'sd-0.033662486283261836, 32'sd-0.1399017859843097, 32'sd-0.10667118088857222, 32'sd-0.02704244481258898, 32'sd0.057472001568598274, 32'sd-0.06017944520327409, 32'sd0.00615500281210537, 32'sd0.0038840736469989445, 32'sd-0.009681626887280755, 32'sd-0.1456845329329316, 32'sd-0.10821031065568042, 32'sd-0.07901214771919933, 32'sd-0.044476019210594894, 32'sd-0.06667313164359571, 32'sd0.03872475029211452, 32'sd-0.08232414432937162, 32'sd0.024782831509874967, 32'sd-0.038055460118002656, 32'sd0.005079886198752959, 32'sd0.11934055699118395, 32'sd0.036841737363706106, 32'sd0.1799775823635961, 32'sd0.1727003563978449, 32'sd0.006501528466938504, 32'sd-0.20038090136628148, 32'sd-0.1807095979615709, 32'sd-0.13351928349990932, 32'sd-0.04231452348500074, 32'sd-0.03612582845258006, 32'sd-0.11103793485005338, 32'sd-0.10127225119430944, 32'sd0.0027325360473503977, 32'sd-0.07253503272601945, 32'sd-0.036366331140542586, 32'sd-0.1387985268532916, 32'sd-0.0905244681134845, 32'sd-0.021214552748306532, 32'sd-0.07850202413348596, 32'sd-0.04623103732585647, 32'sd-0.09423487350161282, 32'sd-0.03220996171014231, 32'sd-0.062235040396261126, 32'sd-0.0018121578943045284, 32'sd0.004497103483714596, 32'sd-0.04333167154134936, 32'sd0.07182986116690672, 32'sd-0.07329821614868902, 32'sd0.06290692032732058, 32'sd0.08856457239493813, 32'sd0.07196503392880402, 32'sd0.1344108671311125, 32'sd0.035718835925698425, 32'sd-0.2648568104316301, 32'sd-0.20084425721960525, 32'sd-0.11850442921115524, 32'sd0.050579682777761904, 32'sd-0.0006453305495202755, 32'sd-0.08564423843457371, 32'sd-0.08573815902908577, 32'sd-0.07615136095767429, 32'sd-0.052485577130218314, 32'sd0.08693885793869045, 32'sd0.05541429950089924, 32'sd0.005017840145744503, 32'sd0.012939010380467316, 32'sd-0.050217817938005296, 32'sd-0.12202498233077215, 32'sd-0.0787919196181697, 32'sd-7.747421847490907e-126, 32'sd0.04269480156504889, 32'sd-0.06196331557273683, 32'sd0.03552428491649458, 32'sd-0.018924432324111992, 32'sd0.13599493396838178, 32'sd0.021577923120197687, 32'sd0.04445311581381494, 32'sd0.08349998195817825, 32'sd0.08749487043107022, 32'sd0.038232672338053095, 32'sd0.07185581826602411, 32'sd-0.18282589192165508, 32'sd-0.16215156495637584, 32'sd-0.03682734738832135, 32'sd-0.06506909692213811, 32'sd-0.08888893087546801, 32'sd-0.15744290599595331, 32'sd-0.04832790422875332, 32'sd0.027602801685520248, 32'sd0.04583721640146427, 32'sd0.01074374980557452, 32'sd-0.050662337334472535, 32'sd-0.10582631888567574, 32'sd-0.02728412723610144, 32'sd-0.0123539968066233, 32'sd-0.10263795523102871, 32'sd-0.056995123282714416, 32'sd-0.0194277785666498, 32'sd0.021206997949056318, 32'sd-0.08670477164678227, 32'sd0.07865589006382484, 32'sd-0.051320648998943605, 32'sd-0.029868726505414972, 32'sd0.14018165482472486, 32'sd0.12201013831111392, 32'sd0.044021735689885724, 32'sd0.0758035491197619, 32'sd0.1417204836702847, 32'sd0.03860858222849449, 32'sd-0.044120946320387655, 32'sd-0.10340431733645816, 32'sd-0.009746541674832972, 32'sd-0.006653875513142912, 32'sd-0.022653054841472453, 32'sd0.025657412464295735, 32'sd-0.003925069344806339, 32'sd0.027135158299629536, 32'sd0.09201999162727709, 32'sd-0.003470957554380235, 32'sd0.060046501459589806, 32'sd-0.09880834958173246, 32'sd0.01565219070697496, 32'sd0.02703802219288423, 32'sd0.008883671546774198, 32'sd0.041353805602139485, 32'sd-0.05956314539817678, 32'sd-0.07542181251396651, 32'sd-0.10078500435587893, 32'sd0.06040126942206177, 32'sd-0.033887065800214014, 32'sd0.015678580203169135, 32'sd0.03713236989331986, 32'sd0.037723627152641055, 32'sd0.09296941928976017, 32'sd-0.005994695630481482, 32'sd0.10728660189437804, 32'sd0.1623855931391038, 32'sd0.09861844248108352, 32'sd0.02570462715487156, 32'sd0.040168831219326226, 32'sd0.052518599661473854, 32'sd-0.07717136156016055, 32'sd0.008785831360930018, 32'sd-0.03525821945572896, 32'sd-0.05554149699754286, 32'sd0.01691883003949053, 32'sd0.03529335807003249, 32'sd0.07693251244785504, 32'sd-0.05371509159356663, 32'sd-0.13940113183863712, 32'sd-0.017127927090999025, 32'sd-0.06736401661587077, 32'sd0.04706583533502201, 32'sd-3.2162627756209417e-125, 32'sd-0.06587150828854049, 32'sd-0.0004992776003914042, 32'sd-0.02904175516306446, 32'sd-0.0358776146932115, 32'sd-0.043767818094581884, 32'sd0.0028677724494728415, 32'sd0.06745568790260605, 32'sd0.030982957954986096, 32'sd0.09913589187245245, 32'sd-0.05984394025121033, 32'sd-0.016770284733863404, 32'sd0.11370096001789112, 32'sd0.07485781308843018, 32'sd0.0824652251617563, 32'sd0.040107379553799505, 32'sd-0.10102880443179207, 32'sd0.0509313785339003, 32'sd-0.05577127234628183, 32'sd0.019712776953147472, 32'sd-0.1352883453402542, 32'sd-0.059177455425376176, 32'sd0.07503321584956725, 32'sd-0.11956291665304536, 32'sd-0.06604467723462709, 32'sd-0.0493537893570793, 32'sd-0.09134831165676353, 32'sd-2.6030086470193165e-126, 32'sd-1.849453231804414e-124, 32'sd-2.137865838269837e-122, 32'sd-0.009258015879794813, 32'sd-0.023198757331033642, 32'sd-0.11489228361610274, 32'sd-0.03330528230818615, 32'sd0.015173168315783732, 32'sd0.004332201294652969, 32'sd-0.0300485368596228, 32'sd-0.010687034366064573, 32'sd0.051040584025647755, 32'sd0.1552637746985823, 32'sd0.23470587241392535, 32'sd0.08678288591251318, 32'sd-0.04830417692396373, 32'sd-0.04018544530876669, 32'sd-0.024820269269888368, 32'sd0.060179348578783896, 32'sd-0.03338929502797525, 32'sd-0.0943346470646554, 32'sd-0.14541493249299425, 32'sd-0.0668973093360618, 32'sd0.02272053376316938, 32'sd-0.05207767514727585, 32'sd-0.06414839361837706, 32'sd-0.08516225909360495, 32'sd-0.07440950925116947, 32'sd-2.7406509524837175e-123, 32'sd-1.0453821281830589e-125, 32'sd1.876683991712574e-126, 32'sd0.016545363322629104, 32'sd0.002160694080659545, 32'sd-0.04087046880354733, 32'sd-0.03570470933852461, 32'sd0.1106908351804991, 32'sd-0.048735084771882, 32'sd0.06713907690657234, 32'sd0.055536261151973805, 32'sd0.07641375668181917, 32'sd0.09029135881449711, 32'sd0.0656030589417411, 32'sd0.06786641144775298, 32'sd0.021090387191484303, 32'sd-0.07352190243812377, 32'sd0.0515727020281583, 32'sd-0.01906921936157498, 32'sd-0.03613451152524805, 32'sd0.021783707462216244, 32'sd0.03600725427275676, 32'sd-0.0549173952615143, 32'sd-0.063359636390718, 32'sd-0.07958547403277177, 32'sd-0.11034021391054201, 32'sd-0.0846407548125143, 32'sd-0.06999716840140954, 32'sd5.387183066965334e-125, 32'sd7.962159252445419e-117, 32'sd6.271921013205145e-116, 32'sd-1.8881055332745734e-125, 32'sd-0.048050594079435176, 32'sd-0.07447325397408636, 32'sd-0.01511253552779658, 32'sd-0.06770872016711592, 32'sd-0.041638303051540176, 32'sd0.0021284638377185613, 32'sd0.03158980573112148, 32'sd-0.005777146352175058, 32'sd0.050635260562622623, 32'sd0.025166314280488416, 32'sd0.06447518582509189, 32'sd0.10509535764877356, 32'sd-0.1383200998885735, 32'sd-0.11371187637251041, 32'sd-0.017992159631901344, 32'sd-0.011938048704570386, 32'sd0.013354190640341575, 32'sd-0.08191072688540632, 32'sd-0.0882446506961793, 32'sd-0.010916034122289319, 32'sd-0.09760738295864914, 32'sd-0.06942490279910793, 32'sd-0.07725913288207178, 32'sd7.761733075056758e-129, 32'sd1.0270037743604062e-121, 32'sd-1.636378404465493e-126, 32'sd-5.9390519185834304e-124, 32'sd2.7704668197473047e-117, 32'sd1.8873097750868623e-117, 32'sd-0.008052596245396833, 32'sd-0.07671013749149722, 32'sd-0.03918675932891396, 32'sd-0.06179720727621401, 32'sd-0.07754854484890003, 32'sd-0.03750779890969645, 32'sd0.04140698299122228, 32'sd0.061140444620929234, 32'sd0.04653150097639899, 32'sd0.09299462000239411, 32'sd-0.015134890503184796, 32'sd0.0819560055487033, 32'sd0.05989903892907359, 32'sd0.04529561183208615, 32'sd-0.08511958774788526, 32'sd0.011667441561046116, 32'sd-0.07697403286243536, 32'sd-0.06744754384871927, 32'sd-0.020632151872670645, 32'sd-0.06123367639284619, 32'sd1.9562022675944195e-118, 32'sd1.4729841692142964e-125, 32'sd-4.821871460069672e-118, 32'sd-2.9517132813488945e-114},
        '{32'sd-3.178232165667208e-116, 32'sd-1.273640224845973e-125, 32'sd1.8622428955808866e-124, 32'sd-7.063815806151492e-117, 32'sd4.184881345889048e-125, 32'sd1.0560575418881105e-127, 32'sd7.844506635652054e-122, 32'sd1.8190188135206717e-123, 32'sd-2.026504304704816e-121, 32'sd2.061046232822533e-124, 32'sd3.5660820129187014e-123, 32'sd7.247996942725282e-119, 32'sd-0.05190818333941244, 32'sd-0.03131381617412387, 32'sd-0.01197436177826024, 32'sd-0.01844646910143864, 32'sd6.10783849531861e-125, 32'sd-4.978784195575481e-127, 32'sd-2.58664056589471e-122, 32'sd-7.303086338151166e-120, 32'sd3.3247504696555998e-118, 32'sd2.2062011327692703e-116, 32'sd7.285516485399792e-121, 32'sd8.793049910621801e-122, 32'sd2.8536115004691265e-121, 32'sd3.65485805687139e-123, 32'sd1.2360661213511948e-118, 32'sd6.528763576847544e-131, 32'sd1.4315336466820435e-116, 32'sd-2.104062208536315e-126, 32'sd3.35919257914906e-120, 32'sd3.919176688064936e-124, 32'sd-0.03335218278098231, 32'sd-0.0028909460876793735, 32'sd-0.036599150141205926, 32'sd-0.02072432931515926, 32'sd0.009023166398651477, 32'sd-0.00468975501429399, 32'sd-0.005218027883353318, 32'sd0.02747508740504216, 32'sd0.008278526553428965, 32'sd0.04570081101193539, 32'sd-0.0042941190183630774, 32'sd-0.04090443735646288, 32'sd0.029309060886523332, 32'sd-0.06417587898721895, 32'sd0.05953811062601043, 32'sd-0.05984075227934625, 32'sd0.007488172162941293, 32'sd0.016115584033340086, 32'sd-0.03784603986207058, 32'sd-0.019511087011685604, 32'sd3.281237403344506e-123, 32'sd-1.248012825820387e-122, 32'sd-2.930469502258637e-123, 32'sd-2.4625502693879934e-121, 32'sd-4.752598060262948e-123, 32'sd3.2869674309694643e-121, 32'sd-0.01934009579368351, 32'sd-0.000868313135548917, 32'sd0.024662100002612188, 32'sd-0.06219414143508273, 32'sd-0.013868872144221413, 32'sd0.025949554701726885, 32'sd0.09837987002906659, 32'sd0.04670533497577504, 32'sd-0.061169249285883485, 32'sd-0.016069664521287674, 32'sd-0.03927341765648583, 32'sd0.026045125172175745, 32'sd-0.014680128602016068, 32'sd-0.022918238360387058, 32'sd-0.03887532089342654, 32'sd0.004223250926216192, 32'sd0.11102399744673153, 32'sd0.09793514562403692, 32'sd0.0704089896187925, 32'sd-0.04644906343941783, 32'sd0.013353509155292676, 32'sd0.03436455123706391, 32'sd0.06201262005600644, 32'sd0.01729528178693254, 32'sd2.5006310908861323e-125, 32'sd4.996022208163588e-124, 32'sd3.815579750391658e-127, 32'sd-7.761519237765785e-123, 32'sd0.05318596242883383, 32'sd0.020073796022396482, 32'sd0.054666866259130226, 32'sd-0.03251372197533772, 32'sd-0.04316856575314836, 32'sd0.06103686575498198, 32'sd-0.014210460783357316, 32'sd-0.06896915578480033, 32'sd-0.0069651847560976265, 32'sd0.14071535204886004, 32'sd0.026248876263944506, 32'sd0.047118487514221735, 32'sd0.013644465408039423, 32'sd-0.04446750242299271, 32'sd-0.09797998417969275, 32'sd0.024844622336954985, 32'sd0.006208522437867849, 32'sd-0.10959224694292365, 32'sd-0.04219902115072249, 32'sd0.023374967578201986, 32'sd-0.0038850565783440905, 32'sd-0.020943460520202413, 32'sd0.06377862812911653, 32'sd0.012565828395929159, 32'sd0.0004916253439044817, 32'sd-3.039127343799257e-125, 32'sd-2.7702418999317e-121, 32'sd-0.0025847720098530307, 32'sd0.001665143199658768, 32'sd-0.07494468638177741, 32'sd-0.06110951713226365, 32'sd-0.00039026421825455275, 32'sd-0.07324612550470601, 32'sd-0.0756642384343242, 32'sd-0.1182670905131931, 32'sd-0.01754403920910837, 32'sd-0.03707852729504809, 32'sd-0.050648984377192084, 32'sd-0.1027229340542722, 32'sd0.06920548650960726, 32'sd-0.0073601274471246396, 32'sd0.06376044747688162, 32'sd-0.05895089072805217, 32'sd0.03174510875217456, 32'sd0.10125903753893371, 32'sd-0.03469297216310144, 32'sd0.00409352149935327, 32'sd0.008274771692274112, 32'sd0.15238111791253345, 32'sd0.08421322414551703, 32'sd-0.06042420327574667, 32'sd-0.08109889318301627, 32'sd-0.05824664674580971, 32'sd-0.01845624387891533, 32'sd-3.38481684078451e-123, 32'sd0.012157519512645413, 32'sd-0.004209715294276402, 32'sd-0.02046664572281472, 32'sd0.06718339149108263, 32'sd0.08957053150860993, 32'sd0.05031958007223054, 32'sd0.0011049823842329395, 32'sd0.04018603073445033, 32'sd-0.011934565129800337, 32'sd-0.046524735256126666, 32'sd0.021098649510803116, 32'sd-0.0075106437859899546, 32'sd0.15679476532168005, 32'sd0.15625714401672247, 32'sd-0.09311715925512429, 32'sd0.005892576800490359, 32'sd0.13124705916170154, 32'sd0.01885762995217652, 32'sd0.009752848926888253, 32'sd0.05625176985231402, 32'sd0.062180786583979616, 32'sd0.03405773965670473, 32'sd0.005797227936450278, 32'sd-0.11800561145927285, 32'sd0.02356282909166497, 32'sd-0.06781032453217595, 32'sd0.057290509357285725, 32'sd-6.882708329277035e-126, 32'sd-0.005578759992207306, 32'sd-0.015368773444169155, 32'sd-0.015710456454390866, 32'sd-0.004489154563675007, 32'sd-0.038739053777731215, 32'sd-0.11105876215103662, 32'sd-0.04365410165936856, 32'sd-0.13724761268298444, 32'sd-0.014715586410384424, 32'sd-0.0031643172488148444, 32'sd-0.006355498686437028, 32'sd0.06889947818187324, 32'sd0.13758762985943368, 32'sd0.08146189772294118, 32'sd0.18624936413842477, 32'sd0.12478658158203507, 32'sd0.24586928790050505, 32'sd0.1616710563350522, 32'sd0.07878861634081485, 32'sd-0.005349034010319099, 32'sd-0.03398108640545081, 32'sd-0.037779529442539046, 32'sd-0.13035205279349818, 32'sd-0.09031424563278864, 32'sd-0.11751114022515471, 32'sd-0.06791276197645546, 32'sd0.06411929147424816, 32'sd0.0022082488248147485, 32'sd-0.04806499580991054, 32'sd-0.0016693268914674186, 32'sd-0.034537666165751366, 32'sd0.06178408590298507, 32'sd-0.07170006696364627, 32'sd0.03502329674383055, 32'sd0.07124385234888318, 32'sd0.09137671328993438, 32'sd0.11103487656581933, 32'sd0.03200877031216616, 32'sd0.026757771581467023, 32'sd0.10102332226698794, 32'sd0.06064192525128094, 32'sd0.04401291470078637, 32'sd0.07947397155135467, 32'sd0.161982719913171, 32'sd0.04812389116081901, 32'sd0.1329921193010915, 32'sd0.11140854568958057, 32'sd0.10223383945211219, 32'sd-0.03756536904029196, 32'sd-0.07355691779538234, 32'sd-0.03829998211417069, 32'sd0.006624034547672947, 32'sd-0.011275371125940138, 32'sd0.03202320728158183, 32'sd0.10496153596634672, 32'sd-0.003541845163643695, 32'sd0.020865067559647784, 32'sd0.02189629581262146, 32'sd0.026209341157562283, 32'sd-0.053107374110911286, 32'sd0.036200673995672075, 32'sd-0.010471796355986643, 32'sd0.014349434141736126, 32'sd-0.02865113124772408, 32'sd0.03241579834901474, 32'sd0.06619368147710815, 32'sd0.07363786271378979, 32'sd0.04053017482334515, 32'sd0.019342207722192733, 32'sd-0.005391458174947399, 32'sd-0.007468594494914334, 32'sd-0.04308175550895223, 32'sd-0.056957976584813, 32'sd0.004324264698365665, 32'sd-0.058969886063419526, 32'sd0.030616265145913833, 32'sd-0.00705276161912784, 32'sd-0.10935916568262263, 32'sd-0.11791139522131684, 32'sd-0.1395256255610832, 32'sd-0.03401406812594518, 32'sd0.014517357000761509, 32'sd-0.03639920356167913, 32'sd-0.003559293214172193, 32'sd-0.04043139852075997, 32'sd0.05027167247207373, 32'sd-0.0546461612023083, 32'sd0.028459552079276692, 32'sd-0.009714358111329894, 32'sd-0.0648710912281709, 32'sd-0.03999320044746711, 32'sd-0.06623435775625008, 32'sd-0.04839643273911534, 32'sd0.06712503140408221, 32'sd-0.04817867579616003, 32'sd-0.09778319651383803, 32'sd-0.14113084267255285, 32'sd-0.06616878484282739, 32'sd-0.046666666953757395, 32'sd-0.06774139915568089, 32'sd-0.0447351328305197, 32'sd-0.043685349516207304, 32'sd0.007856929120500502, 32'sd-0.003318284197632085, 32'sd-0.11049326084985776, 32'sd-0.14412820046380487, 32'sd-0.19019300921671303, 32'sd-0.04861167285459425, 32'sd-0.07335185484915657, 32'sd-0.0053314130446538545, 32'sd-0.058998979064125254, 32'sd-0.04125694841734123, 32'sd0.022103577192598194, 32'sd0.07708063079452716, 32'sd-0.12399673914308922, 32'sd-0.027393991295600262, 32'sd-0.0008245047529720297, 32'sd-0.010105909400480735, 32'sd-0.018079478092707938, 32'sd0.04350825716437509, 32'sd-0.07422669949918494, 32'sd0.042824081838927726, 32'sd0.03369728890855424, 32'sd-0.18015261587218553, 32'sd-0.10292784447729127, 32'sd-0.09769505810810147, 32'sd-0.09988502268733662, 32'sd-0.07831806451769437, 32'sd-0.056451968257967486, 32'sd0.11201483467072783, 32'sd0.010728697213473717, 32'sd-0.03521122569483112, 32'sd-0.11284351588434881, 32'sd-0.040547141876974335, 32'sd-0.03916588552602533, 32'sd0.003181805706892734, 32'sd-0.06502523813125458, 32'sd-0.009590253955581711, 32'sd-0.036047270572500074, 32'sd0.04856431286223879, 32'sd-0.057068315812874186, 32'sd-0.12632655353375255, 32'sd0.0016845562849075756, 32'sd-0.07504617947147484, 32'sd-0.03476042008510506, 32'sd0.0009593377499409798, 32'sd0.07292071683377183, 32'sd0.1268699403912292, 32'sd0.03482992587113982, 32'sd-0.06431086819181085, 32'sd0.02633737641815451, 32'sd-0.05591897239729406, 32'sd-0.005019798411278423, 32'sd-0.08025084083408071, 32'sd-0.10645609821427982, 32'sd0.017901565695382197, 32'sd0.03332401133046237, 32'sd0.07317744657781262, 32'sd-0.03281913388706241, 32'sd-0.02181735028364615, 32'sd-0.0624843350719444, 32'sd0.02712886220898102, 32'sd0.08986400257886464, 32'sd0.059704323830740154, 32'sd-0.01699641784540856, 32'sd0.05915654242399865, 32'sd0.06264415755996446, 32'sd-0.030844051348300885, 32'sd0.019050716154256894, 32'sd0.07255238864615485, 32'sd-0.059233323406615725, 32'sd0.05912928471064561, 32'sd0.0040790194121497585, 32'sd-0.0582208278243248, 32'sd0.11250565838540141, 32'sd0.06184341215330573, 32'sd-0.03223808152653059, 32'sd0.09317179567763699, 32'sd0.07949911099120506, 32'sd-0.007013317929030035, 32'sd-0.03539615995189059, 32'sd-0.11189793325635587, 32'sd-0.0665513643076213, 32'sd-0.008818543712293389, 32'sd-0.08891666871583938, 32'sd-0.06583572504896675, 32'sd-0.0789174468525237, 32'sd-0.03218740665997289, 32'sd-0.029840927361876497, 32'sd-0.003329060636126703, 32'sd0.013370551151063625, 32'sd-0.11694739098498962, 32'sd-0.15003952466426346, 32'sd-0.0831393496792669, 32'sd-0.010004086509823465, 32'sd-0.03155461186244603, 32'sd0.0027691265270169923, 32'sd0.08271019710021707, 32'sd0.013990939955274688, 32'sd0.00533863560890758, 32'sd0.14521575089394484, 32'sd-0.012072570994563842, 32'sd0.005492748741985905, 32'sd0.04127311837836846, 32'sd-0.0018248980816459382, 32'sd0.007189208475565518, 32'sd-0.04703457065303873, 32'sd-0.007006567672940935, 32'sd-0.04233831122580119, 32'sd-0.13813067144188887, 32'sd-0.08181655758910013, 32'sd-0.03907754628167524, 32'sd-0.11307527696391001, 32'sd0.014470866680774118, 32'sd0.013889689142575892, 32'sd-0.038459901778172274, 32'sd-0.09191635113554754, 32'sd-0.14522109603572075, 32'sd-0.0643321831520689, 32'sd0.015146631347458608, 32'sd0.025253309833573993, 32'sd-0.08520037969477764, 32'sd0.017231578191593887, 32'sd0.04672076330500069, 32'sd0.0712920235528409, 32'sd-0.02304952415738892, 32'sd-0.08492202491924757, 32'sd0.016000107540340664, 32'sd0.038232903119497216, 32'sd-0.01315360558966858, 32'sd-0.12002225219339144, 32'sd-0.045340022264122606, 32'sd0.03065796752239193, 32'sd0.16527455070841432, 32'sd0.06682789087551044, 32'sd-0.021649956876067987, 32'sd0.07491038946028118, 32'sd0.02331467467453208, 32'sd-0.13194352001165097, 32'sd-0.08968204597225166, 32'sd-0.04155454743836372, 32'sd-0.004671502699629251, 32'sd-0.08777967581648607, 32'sd0.01937310462911387, 32'sd0.047616808971105186, 32'sd0.06413768250824532, 32'sd0.034111155688878424, 32'sd-0.054550221645226556, 32'sd0.08119295149005734, 32'sd-0.06754519308633648, 32'sd-0.07665495747176988, 32'sd0.09298781791549562, 32'sd-0.04809202930673792, 32'sd-0.07046529136101022, 32'sd-0.03534666070851361, 32'sd-0.12397875821859224, 32'sd-0.0750033016317187, 32'sd-0.15850229775049318, 32'sd-0.05963264342606137, 32'sd-0.11322510013674027, 32'sd0.04614293384554138, 32'sd0.050432455977955454, 32'sd0.06226476156825837, 32'sd-0.012101293115312555, 32'sd0.11929933667021649, 32'sd-0.019641095250052188, 32'sd0.10185198175215755, 32'sd0.025464902379208645, 32'sd-0.0329010676277447, 32'sd0.025557443895335798, 32'sd-0.1382380705120047, 32'sd-0.06850089101758473, 32'sd0.11761751887976107, 32'sd0.06644649264838129, 32'sd0.043815565895945104, 32'sd0.004014268341276134, 32'sd0.006362869034999441, 32'sd0.06591565649180922, 32'sd-0.0450197641690726, 32'sd0.00393650578519462, 32'sd-0.001544667909212704, 32'sd-0.1459969918239318, 32'sd-0.07441785755103988, 32'sd-0.058442510486168074, 32'sd-0.09047548955991244, 32'sd-0.07093783963540529, 32'sd-0.14820618751313122, 32'sd-0.024116318178592774, 32'sd0.042018475421341, 32'sd0.033498033386392054, 32'sd0.05667409371105131, 32'sd0.00544116179958723, 32'sd0.04887432276797144, 32'sd0.09452562803335214, 32'sd0.03154328643761688, 32'sd0.03154490522107791, 32'sd-0.020116178157899168, 32'sd-0.1501911340952899, 32'sd-0.12370538583661167, 32'sd0.005947450804310761, 32'sd0.05548729692611853, 32'sd-0.03981407020479431, 32'sd-0.13067480806413734, 32'sd-0.15809279185701833, 32'sd-0.012386652393627927, 32'sd0.02151877071739785, 32'sd-0.024082636105387113, 32'sd2.826270108700147e-118, 32'sd0.005229846101571997, 32'sd-0.0002393468969970106, 32'sd-0.041823564114388055, 32'sd-0.01627027920619437, 32'sd-0.08738062138072673, 32'sd-0.09825920407668857, 32'sd-0.06064560539583798, 32'sd-0.17904157440371682, 32'sd-0.08037261429859384, 32'sd-0.12107146273968325, 32'sd-0.06156540874706638, 32'sd-0.022522571508085322, 32'sd0.11103004456424642, 32'sd0.058432248294926534, 32'sd-0.010241937470423597, 32'sd0.015810076426741926, 32'sd0.04900130105985571, 32'sd0.056792039628626514, 32'sd-0.0896396757603372, 32'sd-0.06133544359655054, 32'sd0.012299377039079521, 32'sd0.013851715198060222, 32'sd-0.09971957487231957, 32'sd0.0469859818778481, 32'sd0.06177484774181271, 32'sd0.03519461836585362, 32'sd-0.04103016482084, 32'sd-0.029942971960081152, 32'sd-0.003510127556276764, 32'sd-0.10212931733661634, 32'sd-0.007801697996064841, 32'sd0.08378944791329948, 32'sd-0.14259636506075535, 32'sd-0.09893430704419831, 32'sd-0.14690068840576792, 32'sd-0.17194821207160224, 32'sd-0.2359067895908219, 32'sd-0.033612886967919184, 32'sd-0.025050927937070026, 32'sd0.10204641972590119, 32'sd-0.038174005374618895, 32'sd0.011243085136882635, 32'sd0.0051962847809400884, 32'sd0.1649024130185118, 32'sd0.10984304450199746, 32'sd0.0333355060733408, 32'sd-0.10622192796319914, 32'sd-0.12568991710708627, 32'sd0.04304191944161877, 32'sd-0.050804442026725675, 32'sd-0.0742163869708692, 32'sd-0.04261511642898719, 32'sd0.037204839176673034, 32'sd0.06672778650265278, 32'sd-0.04675342746744905, 32'sd-0.033056505959935784, 32'sd-0.07053826079688393, 32'sd0.06411435843470102, 32'sd-0.05689194059503459, 32'sd0.05229007364435106, 32'sd-0.07995327264018988, 32'sd-0.10873560708211653, 32'sd-0.17262780306284883, 32'sd-0.17633126686593661, 32'sd-0.19911347589177678, 32'sd-0.23733692527283884, 32'sd-0.11177242895068651, 32'sd0.00044932528862224924, 32'sd-0.07414208640406589, 32'sd0.028223197230534326, 32'sd0.01558069133715965, 32'sd-0.04663329336117122, 32'sd0.07825910864948671, 32'sd-0.020562826902324492, 32'sd-0.009970197820633934, 32'sd-0.10996223507672119, 32'sd0.027662499742835946, 32'sd-0.00013431689496835267, 32'sd-0.03318651250445742, 32'sd0.1011328051019861, 32'sd-0.005868782714315671, 32'sd-0.0333522832880005, 32'sd0.0227150051431339, 32'sd9.99891032091784e-122, 32'sd-0.019637882826934117, 32'sd0.09657190635589104, 32'sd0.1133154149773919, 32'sd-0.003770669748685348, 32'sd-0.10083200594957692, 32'sd-0.051128145701500746, 32'sd-0.03628152818073727, 32'sd-0.01629601737463636, 32'sd-0.25599328784969516, 32'sd-0.15206788544475075, 32'sd-0.09552104358755704, 32'sd-0.013727422016580488, 32'sd-0.10419177035759908, 32'sd-0.09559725657664027, 32'sd-0.06165037142625863, 32'sd-0.0937754204395602, 32'sd-0.03266561764789716, 32'sd-0.13379413457702669, 32'sd-0.11776708253066755, 32'sd0.015000090290736609, 32'sd-0.008943698466122595, 32'sd0.039976029575339016, 32'sd-0.031023772986050562, 32'sd0.03327526512481553, 32'sd-0.041052247581601274, 32'sd-0.029018338288691298, 32'sd-0.01966586811433162, 32'sd-0.022406738211121897, 32'sd-0.015034012067505428, 32'sd0.0020340755589564204, 32'sd0.0920001187838139, 32'sd0.05717478746962896, 32'sd0.00505770623383455, 32'sd-0.057194575260836315, 32'sd0.04660626510625303, 32'sd-0.029331328420259678, 32'sd-0.07391703201659691, 32'sd0.0919793313962873, 32'sd-0.008656992472633704, 32'sd-0.04001637500087818, 32'sd0.005681558462718674, 32'sd-0.024540855327479662, 32'sd0.02327661157794952, 32'sd0.0075564889193923965, 32'sd-0.07282481119611374, 32'sd-0.023248846739111432, 32'sd-0.10251993439439427, 32'sd-0.17764626802573613, 32'sd0.05643868562400882, 32'sd-0.009731688239308622, 32'sd-0.04838857161208222, 32'sd-0.05924513687580056, 32'sd-0.0595464366528179, 32'sd0.06802255699825198, 32'sd0.03668182085823855, 32'sd0.011058882944866233, 32'sd-0.02430765536652892, 32'sd0.041815036772578876, 32'sd0.08953764028624563, 32'sd-0.06970298592105346, 32'sd-0.004603607366017926, 32'sd0.056282844849990216, 32'sd0.03506059238796054, 32'sd0.023301546680460437, 32'sd0.030407178572753272, 32'sd0.0892345531750653, 32'sd0.024297593878908418, 32'sd0.13897968578979814, 32'sd0.032564350235510436, 32'sd0.09132153710420864, 32'sd-0.0327661643603432, 32'sd-0.17644042131090548, 32'sd0.055488280512466986, 32'sd-0.08305581086682783, 32'sd-0.1548287530763054, 32'sd-0.013987138927566815, 32'sd0.010972314205782391, 32'sd-0.048407552861504465, 32'sd-0.1101887710403982, 32'sd-0.04392880000098581, 32'sd-0.04036436792048122, 32'sd-0.05732852705694063, 32'sd0.009815997499048252, 32'sd-4.591843813266732e-122, 32'sd-0.0019762441800180025, 32'sd-0.059219941329673086, 32'sd0.00864138288794722, 32'sd0.016992941574812584, 32'sd0.08337922635384135, 32'sd0.1469488335708825, 32'sd0.03688520802812027, 32'sd0.010375596582591733, 32'sd-0.017092070572671664, 32'sd0.10091466956871341, 32'sd0.13510471126150467, 32'sd0.005610596434500022, 32'sd0.14607765333470343, 32'sd0.06405307277746153, 32'sd-0.0433298286530456, 32'sd-0.17425326537987937, 32'sd-0.1935529680626486, 32'sd-0.07093749396555993, 32'sd-0.14431133270609908, 32'sd-0.08933687077545095, 32'sd-0.03933203622127695, 32'sd0.04422064090369658, 32'sd0.029228313422264417, 32'sd0.020030661639944148, 32'sd0.05033201849468074, 32'sd-0.0458771699213689, 32'sd-3.8243358239749633e-116, 32'sd9.641112070642699e-116, 32'sd2.8013664837285928e-115, 32'sd0.04047712807897053, 32'sd-0.0615066311867657, 32'sd0.029547754723242444, 32'sd-0.021650350294109645, 32'sd0.07442515934429138, 32'sd0.013855162432840157, 32'sd0.061438476568533795, 32'sd0.05749337724690529, 32'sd0.11552333706741343, 32'sd0.016841796307572134, 32'sd0.04286874242030901, 32'sd-0.011168326709738031, 32'sd0.04434820044177109, 32'sd0.047475878929520196, 32'sd-0.20630599183624432, 32'sd-0.23445755641712998, 32'sd-0.16888227675661785, 32'sd-0.1757118120156598, 32'sd-0.005856660850144941, 32'sd-0.01112017677554646, 32'sd-0.04636814679505942, 32'sd-0.011258456977359143, 32'sd-0.021273360146221408, 32'sd-0.12042363813684141, 32'sd-0.014937118237393533, 32'sd-1.3797503082935262e-115, 32'sd6.469327638134299e-124, 32'sd-2.7357489892829676e-121, 32'sd0.05513067969014506, 32'sd-0.0028957583604778477, 32'sd0.030805195489469646, 32'sd-0.029541991038901007, 32'sd-0.1272391085293792, 32'sd0.08857393932287327, 32'sd-0.014194624114189546, 32'sd-0.06282799706812857, 32'sd0.010149645134316276, 32'sd0.09507540945520908, 32'sd0.11271465024890581, 32'sd0.1335547250804177, 32'sd-0.048471327450275443, 32'sd-0.07957077311148829, 32'sd0.02724482901517983, 32'sd-0.050586749125464084, 32'sd0.0531735588913268, 32'sd-0.03888613782641977, 32'sd-0.0379468262970787, 32'sd0.08400753001695048, 32'sd0.049089348384554, 32'sd0.050502140581399, 32'sd-0.055682119671792124, 32'sd-0.0416268503386943, 32'sd-0.023562293690106734, 32'sd2.2546855715570107e-116, 32'sd1.5158221510413924e-124, 32'sd-8.594061901932895e-117, 32'sd-1.3095821642422558e-118, 32'sd-0.027163151320190752, 32'sd-0.010058435652258056, 32'sd-0.00583205423684882, 32'sd0.03802054491111687, 32'sd-0.07824166324927542, 32'sd-4.410696218973898e-05, 32'sd0.1021460272100937, 32'sd0.15000380102587182, 32'sd0.15472997469802774, 32'sd0.04986225897602019, 32'sd0.16681151075402012, 32'sd0.062057189306451675, 32'sd-0.041611251730319675, 32'sd-0.08990540754437691, 32'sd0.067535735785233, 32'sd-0.0010884992698513617, 32'sd-0.030850624257868865, 32'sd0.0046789913373463205, 32'sd0.06389933772379001, 32'sd-0.02099336635951195, 32'sd-0.044152645086253384, 32'sd0.04052590830468415, 32'sd-0.02730406784404743, 32'sd-4.230983818076809e-118, 32'sd-3.823512654592185e-116, 32'sd-3.1057799688467617e-127, 32'sd3.71073829732101e-116, 32'sd2.3712589065048053e-126, 32'sd3.3722524694027756e-120, 32'sd0.020446165368886292, 32'sd0.009323570383887021, 32'sd0.01913808720959935, 32'sd0.03182614219085104, 32'sd0.024589945583762863, 32'sd0.004517798533484597, 32'sd0.057140206203218497, 32'sd0.1013830889321225, 32'sd-0.013893307075876847, 32'sd0.031100895353247577, 32'sd0.10849943460795847, 32'sd0.08778968657758823, 32'sd0.07429292772296642, 32'sd0.033508144291791095, 32'sd0.08362961836237592, 32'sd0.09287956719271542, 32'sd0.12025643229063451, 32'sd-0.054862536834241464, 32'sd-0.08756850801622816, 32'sd0.008149219191820076, 32'sd1.2678939426685674e-115, 32'sd-3.809632605524883e-123, 32'sd-4.50293945068612e-117, 32'sd-8.59473407338148e-122},
        '{32'sd-1.9174416259053567e-121, 32'sd-1.064082883725278e-119, 32'sd-5.258759208192989e-115, 32'sd-3.5981486524287384e-121, 32'sd3.741310886611454e-122, 32'sd1.4352599457525756e-118, 32'sd2.2140089452046894e-125, 32'sd-3.833677855306148e-126, 32'sd-4.609123053047049e-122, 32'sd-1.6780271167396494e-123, 32'sd1.1632017983592289e-116, 32'sd-6.857307517086328e-126, 32'sd0.06430613695141547, 32'sd0.054518630106769765, 32'sd0.034206786278280256, 32'sd0.012300029079406293, 32'sd6.025450816493213e-124, 32'sd-1.5295268128936734e-126, 32'sd-4.756770875055464e-123, 32'sd4.298386733658924e-117, 32'sd1.062016812359005e-124, 32'sd8.922031788051981e-119, 32'sd4.0582155180217025e-125, 32'sd1.6917435678130803e-125, 32'sd-1.0578131848283958e-124, 32'sd3.3572734778059706e-121, 32'sd-3.4266840208967176e-123, 32'sd-5.744427518896481e-115, 32'sd-6.130335473325089e-122, 32'sd9.861064636170924e-121, 32'sd-5.305012420938208e-127, 32'sd8.880227365285885e-123, 32'sd-0.006005539456005898, 32'sd0.047223266785782377, 32'sd-0.003677780976690518, 32'sd0.02782588801124432, 32'sd0.11065920168093812, 32'sd-0.026811164735088697, 32'sd0.07797607458974803, 32'sd0.04925716913132526, 32'sd0.04308382077243413, 32'sd-0.06206757443617972, 32'sd-0.0361257837355485, 32'sd-0.04292155863960705, 32'sd0.017617142931493714, 32'sd0.06386747327260169, 32'sd0.014072155717752, 32'sd0.025561138580216664, 32'sd0.03541200716813443, 32'sd0.0286690816650414, 32'sd0.04008723769521291, 32'sd0.08395770626876536, 32'sd1.8931803728486085e-119, 32'sd1.2127838716572336e-118, 32'sd-3.3098885683020783e-121, 32'sd1.6172430537678277e-122, 32'sd-1.8628221008131332e-123, 32'sd-1.6795274331136705e-126, 32'sd0.10246615868760907, 32'sd0.030128688306659882, 32'sd-0.009802297775459181, 32'sd0.06759924212905516, 32'sd0.08752921843488604, 32'sd0.10161498366173627, 32'sd-0.040990005367447534, 32'sd-0.014269748246377348, 32'sd0.054593739838222334, 32'sd0.03282907806658113, 32'sd0.10572687482133897, 32'sd0.04724414708257162, 32'sd-0.07812166286416557, 32'sd0.0316420248575622, 32'sd-0.051414574284281964, 32'sd0.07012691176518439, 32'sd0.09508017680278143, 32'sd0.014662648674298062, 32'sd0.10258598475435417, 32'sd0.015021748743553725, 32'sd0.1041792293627228, 32'sd-0.002999769560684012, 32'sd0.0026060562006642875, 32'sd0.08588833468939593, 32'sd7.63929346986693e-121, 32'sd-1.3954555786438005e-124, 32'sd1.2068848529349344e-126, 32'sd1.423629621386271e-118, 32'sd0.09857103939830898, 32'sd0.028710224308940203, 32'sd-0.039483138448895234, 32'sd0.13137577460444547, 32'sd0.03024844113329249, 32'sd-0.14197332440778945, 32'sd-0.011747750873271876, 32'sd0.00907695555885663, 32'sd0.07428316812938009, 32'sd-0.03635186560353336, 32'sd0.11910348440626461, 32'sd0.10955977442200728, 32'sd0.0030508042890575976, 32'sd-0.16976170422067857, 32'sd0.03365496723572253, 32'sd0.10142376761439129, 32'sd-0.03022593331250128, 32'sd-0.038893884113042586, 32'sd-0.028869681193023307, 32'sd-0.012441388531525125, 32'sd-0.022906483299236686, 32'sd-0.03556827882048698, 32'sd0.018759017248931427, 32'sd-0.07029462794415316, 32'sd0.019136609569016503, 32'sd4.5319114529681474e-123, 32'sd6.436716580827755e-118, 32'sd0.07412694482732216, 32'sd0.0822466600382327, 32'sd-0.004460466189083929, 32'sd0.08626377712075518, 32'sd-0.045510570839192674, 32'sd-0.004247222539590384, 32'sd0.0355876292561427, 32'sd-0.031625373223446475, 32'sd-0.013995723025107355, 32'sd0.10008425273493146, 32'sd0.004544440224108608, 32'sd0.04282342056211986, 32'sd0.022566930750084018, 32'sd0.10097661645523347, 32'sd0.06048470219270294, 32'sd-0.028510977885640866, 32'sd0.027143660005227742, 32'sd0.031489477414281354, 32'sd0.005617317250708068, 32'sd0.06395201203997021, 32'sd-0.0425224423107929, 32'sd-0.09236916107391095, 32'sd0.04484254902293246, 32'sd-0.0747938813384203, 32'sd0.04626943209698817, 32'sd0.050392011391137394, 32'sd-0.035533875025309185, 32'sd-9.964274599206299e-120, 32'sd0.023650683198573698, 32'sd0.0238058985281599, 32'sd0.05221744705255625, 32'sd0.0476032715864257, 32'sd0.02918724735433062, 32'sd-0.09302882679660494, 32'sd0.010941703430472394, 32'sd0.043168994908430625, 32'sd-0.053651965796896024, 32'sd-0.0022097509977174134, 32'sd-0.0041799982911988436, 32'sd0.0739248399264076, 32'sd0.14554340907421115, 32'sd0.0736368282216288, 32'sd0.00789222821803541, 32'sd0.08007791324218183, 32'sd0.09471670790838595, 32'sd-0.05359789024822531, 32'sd-0.06307223597545898, 32'sd-0.08122331135111907, 32'sd0.04332605367413422, 32'sd0.011730072381004878, 32'sd0.04861553768164083, 32'sd0.03598041561428791, 32'sd0.050827243814500926, 32'sd-0.04583652085568894, 32'sd0.08897401335776434, 32'sd-2.138107015940739e-120, 32'sd0.07064297641022142, 32'sd-0.018930242142231823, 32'sd0.0353073536783477, 32'sd-0.009873814292836227, 32'sd0.06535405972219224, 32'sd-0.046015187034697334, 32'sd-0.14658623175799212, 32'sd0.034329615312817294, 32'sd-0.07487715271128527, 32'sd-0.04863458834580969, 32'sd-0.042619193679355585, 32'sd-0.0240931830306837, 32'sd0.11816576979790876, 32'sd0.03142361898858448, 32'sd-0.005301928918458501, 32'sd-0.01890887389741571, 32'sd-0.10848702460675032, 32'sd-0.050880460347912784, 32'sd-0.07758184809012171, 32'sd-0.02014679810007432, 32'sd0.12912357970773558, 32'sd0.014714117244039347, 32'sd0.0955966729862712, 32'sd0.02836440078716297, 32'sd0.0008054979237550481, 32'sd0.03275280551102962, 32'sd0.0019489064497419943, 32'sd0.08489724999115426, 32'sd0.026975004312084296, 32'sd0.09111644940826923, 32'sd0.013164971836129507, 32'sd0.024050805696117783, 32'sd0.06390450785211049, 32'sd0.04509074289788938, 32'sd0.02591355721929874, 32'sd-0.10382418860878305, 32'sd-0.032638849983670226, 32'sd0.03653563542994144, 32'sd-0.02282733155852384, 32'sd0.056786751956323475, 32'sd-0.030034797246837452, 32'sd0.042295435171867644, 32'sd0.09157203881310604, 32'sd0.10781083824270316, 32'sd0.1021260082300904, 32'sd0.011025569572724773, 32'sd-0.018772951100482146, 32'sd0.11571115000122957, 32'sd0.15133090304505, 32'sd0.04522090232505515, 32'sd-0.019153764558603455, 32'sd0.10473630679165588, 32'sd0.07570457440113869, 32'sd-0.0626972839319223, 32'sd0.05402982696248177, 32'sd0.08653180372761432, 32'sd-0.018382047978417287, 32'sd0.06493210129345517, 32'sd0.06032318875908754, 32'sd0.065734570016936, 32'sd0.08168237777998075, 32'sd0.08251463860406989, 32'sd0.13828112083185687, 32'sd0.05944403586780433, 32'sd0.061350853166594985, 32'sd0.026134216913332446, 32'sd-0.056224125943574704, 32'sd0.0352935365626909, 32'sd-0.0006021763445329485, 32'sd-0.009816400494687415, 32'sd0.1350129128981447, 32'sd0.07789471660750004, 32'sd0.0024558228214368147, 32'sd0.006685717321693392, 32'sd0.0315813906668258, 32'sd0.07361110596192001, 32'sd0.09599359775788832, 32'sd-0.05301099776422412, 32'sd-0.06893852080535273, 32'sd0.022197504709897214, 32'sd0.036308550842473405, 32'sd0.10596465236299753, 32'sd0.08741230490876767, 32'sd0.03166335972949297, 32'sd0.08974217123119177, 32'sd0.08725517588283789, 32'sd0.015560590480670189, 32'sd-0.031382257727682224, 32'sd0.047092579883291345, 32'sd0.01313493096834378, 32'sd0.05622607424312329, 32'sd-0.0992753005798059, 32'sd-0.023533083689183363, 32'sd-0.04240592519106036, 32'sd-0.06342887369479083, 32'sd-0.0010743254211848113, 32'sd0.07754435787425619, 32'sd-0.1418651939430515, 32'sd-0.13530418017299742, 32'sd-0.08546882168425825, 32'sd-0.04933606553624739, 32'sd-0.06482009967923436, 32'sd-0.01787197838062208, 32'sd0.09568372689112173, 32'sd0.020404515928184833, 32'sd-0.033668845589381616, 32'sd-0.021761102161415677, 32'sd0.03549621044227509, 32'sd0.04863880232096154, 32'sd0.005076307433415467, 32'sd-0.10029114567065985, 32'sd-0.003473347161993324, 32'sd0.01916036180903988, 32'sd0.009722692993001441, 32'sd0.13849518735032795, 32'sd-0.032500763354339914, 32'sd-0.007432926866736332, 32'sd-0.011951817272106303, 32'sd-0.11858851518684163, 32'sd-0.09834567849665446, 32'sd-0.05573430596117518, 32'sd0.0203967977030064, 32'sd0.040050171691190434, 32'sd0.0790911172579482, 32'sd-0.059046079675522126, 32'sd-0.07494390696727937, 32'sd-0.20039572373521633, 32'sd-0.15728524094806468, 32'sd-0.15516972516602603, 32'sd-0.07058615858630955, 32'sd-0.1196158202012063, 32'sd0.014484866375644107, 32'sd0.1616382864665262, 32'sd-0.027005533703586077, 32'sd0.03793832181782463, 32'sd0.016148697076220766, 32'sd0.07996482608133332, 32'sd0.1249709512358704, 32'sd0.005119914882446274, 32'sd-0.01226692793488981, 32'sd0.04677595451890445, 32'sd0.03807933352993329, 32'sd0.06462329837875491, 32'sd0.029592993692528113, 32'sd-0.04889357468718473, 32'sd-0.008820290809242876, 32'sd-0.013949430058488095, 32'sd0.04517149736078413, 32'sd0.05923497427620554, 32'sd-0.024384144438576238, 32'sd-0.023329486545326364, 32'sd-0.11412218173487637, 32'sd-0.10576965562596853, 32'sd-0.07024165140286895, 32'sd-0.09703749767450882, 32'sd-0.05541635092704765, 32'sd-0.12141335648356705, 32'sd-0.13863948970370749, 32'sd-0.027360737065328523, 32'sd-0.10307788830633978, 32'sd-0.08679359176917321, 32'sd0.08242663312015946, 32'sd0.22389116678915835, 32'sd0.035980741707215436, 32'sd0.07188001201329806, 32'sd0.019475917952194676, 32'sd-0.0009129844185360346, 32'sd0.03675905947680618, 32'sd-0.03214820886213709, 32'sd-0.05529811733447796, 32'sd0.03167938457839234, 32'sd0.07245514725170944, 32'sd-0.029991637672159316, 32'sd-0.01171477726065126, 32'sd0.058318448571379494, 32'sd0.13316408929759332, 32'sd-0.005462463820832472, 32'sd-0.0016487857792257937, 32'sd0.036576321073289876, 32'sd0.02728067240257589, 32'sd-0.042724638733892026, 32'sd0.035085474643676375, 32'sd-0.08470670684898604, 32'sd0.021182368560940423, 32'sd-0.0010974587087796892, 32'sd-0.022597842691626274, 32'sd-0.13381623188086725, 32'sd-0.1003838226941572, 32'sd-0.07290140510187171, 32'sd0.005908803808749931, 32'sd0.07342989130887821, 32'sd-0.007467637445501802, 32'sd-0.02840526013542934, 32'sd0.04220167529993591, 32'sd-0.03502621160236817, 32'sd0.04605525062841655, 32'sd-0.009447246332370549, 32'sd0.04740042558141101, 32'sd0.011478409488600119, 32'sd-0.04242958759394839, 32'sd0.07575555262890875, 32'sd0.0688068722363832, 32'sd0.10651779178102912, 32'sd0.11058801667141457, 32'sd-0.0038373744197468624, 32'sd0.16427591865002628, 32'sd0.09629058469328429, 32'sd0.10156722938443136, 32'sd0.16161853350554106, 32'sd0.1103406597943042, 32'sd-0.012658767307544162, 32'sd0.04220491758830964, 32'sd-0.10536625770146169, 32'sd0.043020753558521314, 32'sd-0.15041113768380235, 32'sd0.014563892754669724, 32'sd-0.06995709645114268, 32'sd-0.024081598353126107, 32'sd0.06995531111067503, 32'sd-0.026671272686573648, 32'sd-0.012300957428998218, 32'sd0.035021928983548514, 32'sd-0.013673401487575645, 32'sd0.14719319109439474, 32'sd-0.03505288967045727, 32'sd-0.014518464562830641, 32'sd-0.0881848385361464, 32'sd0.017284698221316244, 32'sd0.018124535267599003, 32'sd0.005070816543891885, 32'sd0.13015191968125478, 32'sd0.12707081625675976, 32'sd0.06226368105519063, 32'sd0.1330054771966317, 32'sd0.11800737240083524, 32'sd0.020929139640172987, 32'sd0.21845381900569402, 32'sd0.24528894586554154, 32'sd0.17215011048196072, 32'sd0.05409186417378168, 32'sd-0.06433081459813539, 32'sd0.0003014158561143357, 32'sd-0.029644992641581516, 32'sd0.06408829510125617, 32'sd0.01930227413495414, 32'sd-0.012687673428692573, 32'sd-0.11450152640107815, 32'sd-0.0676382197122539, 32'sd-0.07896753129631214, 32'sd0.07312988954025301, 32'sd0.033084411861392736, 32'sd0.11172362450457111, 32'sd0.03308897846869587, 32'sd-0.05952879787313519, 32'sd-0.09928024694934606, 32'sd-0.048199194399519134, 32'sd0.06115471207192571, 32'sd0.05970744072330671, 32'sd0.019651834992438947, 32'sd-0.0739278265243328, 32'sd0.04710681094269705, 32'sd0.11029963599976086, 32'sd0.22458870802188854, 32'sd0.16573621931835933, 32'sd0.2651147766020162, 32'sd0.22170301028537515, 32'sd0.15073519254991946, 32'sd0.07381566822667429, 32'sd0.035917002226936036, 32'sd0.1012172445659089, 32'sd-0.10381956504275489, 32'sd-0.03347994333533369, 32'sd0.08268806263037873, 32'sd0.13419634065789485, 32'sd-0.10065745227192291, 32'sd-0.1251400948976373, 32'sd-0.017797004847787543, 32'sd0.08863637659413434, 32'sd0.014206568723901266, 32'sd0.05980542916462936, 32'sd0.07338888989348485, 32'sd0.06948468524651574, 32'sd-0.034215979263073834, 32'sd0.028137264498412567, 32'sd-0.015090354401071388, 32'sd-0.04205917628894215, 32'sd-0.1357523628468708, 32'sd-0.3053294994537075, 32'sd-0.13779591756093346, 32'sd-0.05236686595864358, 32'sd0.05043797406470191, 32'sd0.2216876956955188, 32'sd0.048552183401577194, 32'sd0.06676913767951288, 32'sd0.03993513543317658, 32'sd0.06897204363688224, 32'sd0.020710876513967216, 32'sd0.1678681955849158, 32'sd0.027925219735153856, 32'sd0.03114328450785806, 32'sd0.011242840330219031, 32'sd0.06559720000863933, 32'sd-0.12534501119880637, 32'sd-0.06376099991886469, 32'sd0.11128135002453937, 32'sd0.13360792806708938, 32'sd0.08911412074839632, 32'sd-2.4184729767938807e-124, 32'sd0.045865103464842884, 32'sd-0.059371752208178225, 32'sd-0.04781675829322016, 32'sd-0.08354680371796974, 32'sd-0.1194417782092694, 32'sd0.014962603573856035, 32'sd-0.0976697854860151, 32'sd-0.14749521500366788, 32'sd-0.12059596199842053, 32'sd-0.1528506568398438, 32'sd-0.23890431269638177, 32'sd-0.13640571591187853, 32'sd-0.1706946627381161, 32'sd-0.15905922989773255, 32'sd0.10317447484947243, 32'sd0.17401058706262054, 32'sd0.09435682394632447, 32'sd0.06838512325945147, 32'sd0.11014726067571819, 32'sd0.09220343412113334, 32'sd0.12230691144123067, 32'sd0.10667698588462077, 32'sd-0.08725800562968246, 32'sd0.08235515819235031, 32'sd-0.022844070951421342, 32'sd0.05711208749209926, 32'sd0.03264158139974681, 32'sd0.014542628379810749, 32'sd0.08396430013320973, 32'sd0.014486723942079952, 32'sd-0.15063143034406004, 32'sd-0.019504555775958096, 32'sd-0.029119318183439876, 32'sd-0.09389068536952637, 32'sd-0.15511841490934988, 32'sd-0.1610317007099992, 32'sd-0.32172931514805336, 32'sd-0.1887245183403594, 32'sd-0.2403328432602668, 32'sd-0.23335674076262122, 32'sd-0.3603053810043955, 32'sd-0.14288172996502557, 32'sd-0.05208781974235208, 32'sd0.020505847176793983, 32'sd0.12084732388081962, 32'sd-0.014521735407353832, 32'sd0.04206695744068014, 32'sd0.05672900273865121, 32'sd0.0807046822292509, 32'sd-0.01996734828663799, 32'sd-0.08361968338772889, 32'sd0.04658509799345655, 32'sd-0.03204792540006539, 32'sd-0.0029596772881525634, 32'sd-0.06398844156870183, 32'sd0.0440457308391374, 32'sd0.030733942074634157, 32'sd-0.0402718859508028, 32'sd0.028114870510280984, 32'sd0.03910106024556614, 32'sd-0.08573603835581073, 32'sd-0.08590773676165689, 32'sd-0.12909758743644428, 32'sd-0.2749068332126769, 32'sd-0.17732871655142418, 32'sd-0.253109593770419, 32'sd-0.23666927067181925, 32'sd-0.1362867996538002, 32'sd-0.26891197597328675, 32'sd-0.14587144663694462, 32'sd-0.12489565912819109, 32'sd0.01084455921062884, 32'sd0.03211623198379107, 32'sd0.13192975371856536, 32'sd-0.09529551630396071, 32'sd0.0544400741259835, 32'sd0.09863436985671575, 32'sd-0.007535252443135509, 32'sd-0.13091958855815447, 32'sd-0.07106910022363973, 32'sd0.10144982191216445, 32'sd0.10526713236981462, 32'sd-0.033299480657516985, 32'sd4.453307658698796e-126, 32'sd-0.015248889964811855, 32'sd0.07083954044345014, 32'sd0.006678252615907971, 32'sd0.01564654524749239, 32'sd-0.09626029798579731, 32'sd-0.037915700416744996, 32'sd-0.06265173178987149, 32'sd-0.08377863663400859, 32'sd-0.08809663595724099, 32'sd-0.039473571744197695, 32'sd-0.03185324274910651, 32'sd-0.054568001546704076, 32'sd-0.016301534093422523, 32'sd0.05355763043272577, 32'sd-0.0959731078826114, 32'sd0.0746016460220017, 32'sd0.1331647934123552, 32'sd0.18441254570620927, 32'sd0.05330664589974266, 32'sd0.09304869817480917, 32'sd0.0795965131578147, 32'sd0.032180650724100375, 32'sd-0.13280182487343367, 32'sd-0.0013997933947118499, 32'sd-0.025325756061734817, 32'sd-0.021095586411802304, 32'sd0.036033322669214204, 32'sd0.032657330738397876, 32'sd0.03897850888944221, 32'sd0.08860770934342532, 32'sd-0.0224243625760971, 32'sd0.21126147356021632, 32'sd0.04779667035291574, 32'sd0.13730411696295566, 32'sd0.07841768968006439, 32'sd0.06015444958921796, 32'sd-0.08622500167175506, 32'sd0.1152964413091525, 32'sd0.08950528046171352, 32'sd0.08084941435303997, 32'sd0.1363422647998775, 32'sd0.10162193249916913, 32'sd0.01041250642974661, 32'sd0.0388961012816347, 32'sd0.004724454863390431, 32'sd-0.021552323940728462, 32'sd0.03316181096109714, 32'sd0.13095961249194185, 32'sd-0.02501248065667962, 32'sd-0.05179003980630147, 32'sd-0.08235753849461196, 32'sd-0.11569149505893453, 32'sd0.08465271735045685, 32'sd-0.09554747009862433, 32'sd0.07154567766671707, 32'sd0.05265508258915227, 32'sd-0.02887386508114118, 32'sd-0.009736703630324528, 32'sd-0.04846651224877408, 32'sd0.12395581476502843, 32'sd0.13494428970594358, 32'sd0.05464458933775742, 32'sd0.13999927203600265, 32'sd0.06707580628913046, 32'sd-0.05329658383265725, 32'sd0.08335703310629979, 32'sd0.13727582033869448, 32'sd0.13373674579786338, 32'sd0.09938757607485069, 32'sd-0.04899957189724179, 32'sd0.09218962780843155, 32'sd0.014800296306621503, 32'sd-0.03920146877744038, 32'sd-0.10162995648944392, 32'sd0.02941837064324411, 32'sd0.03766320098708986, 32'sd-0.026003887765600357, 32'sd-0.20733968417144139, 32'sd-0.015561943249473954, 32'sd-0.06733047117817097, 32'sd0.003696686293472551, 32'sd0.04906225963491886, 32'sd0.04594187904068353, 32'sd-3.4366477550136424e-116, 32'sd0.07842619027607592, 32'sd0.04747582114915196, 32'sd0.10221775834583645, 32'sd0.03234078125563656, 32'sd0.07337662271517902, 32'sd-0.12600431737362397, 32'sd-0.10783716580436024, 32'sd0.0989236349872547, 32'sd0.061617038328221206, 32'sd0.17940029692368448, 32'sd0.20220733213661046, 32'sd0.12250982773095077, 32'sd0.11914008774958575, 32'sd0.008814095785814676, 32'sd0.008421779544183898, 32'sd-0.011971162329396646, 32'sd-0.07693828599637038, 32'sd-0.040996999049361736, 32'sd0.03968092686498749, 32'sd0.013015775472113059, 32'sd-0.14159393324057762, 32'sd-0.0028241515755700075, 32'sd0.00356848039851032, 32'sd-0.03227795859188163, 32'sd0.031516986447735984, 32'sd0.0039208479175715984, 32'sd3.345972321678406e-119, 32'sd-1.5722541003304484e-123, 32'sd-1.81548320293016e-124, 32'sd0.011000961580702621, 32'sd0.09239297788661982, 32'sd0.008793799851775131, 32'sd-0.008177499437961628, 32'sd0.026245516044524922, 32'sd-0.09427327825637076, 32'sd-0.02387159542794036, 32'sd0.013329017980167918, 32'sd0.07399570799876748, 32'sd0.13176434076904578, 32'sd0.12393793721717117, 32'sd0.05249311255645393, 32'sd0.02384710504362452, 32'sd0.0863952946801561, 32'sd0.041463897947917015, 32'sd0.023269248227799008, 32'sd-0.040942454804672575, 32'sd-0.01606451725726282, 32'sd-0.009040590987071244, 32'sd-0.024110831458601992, 32'sd-0.026081460992125223, 32'sd-0.0893560269130151, 32'sd0.04845268731710806, 32'sd0.03583118143855003, 32'sd-0.018501902449145353, 32'sd3.642180248575903e-119, 32'sd-6.5948076637470426e-127, 32'sd4.327685902862792e-125, 32'sd0.024960660210401997, 32'sd-0.009752316227488506, 32'sd0.027198736950218568, 32'sd0.06640524700581645, 32'sd0.05967031651175352, 32'sd-0.06833692113220496, 32'sd0.00590873844786, 32'sd0.10934190910595852, 32'sd0.1117954308908545, 32'sd0.06130815158169605, 32'sd0.11209838119566272, 32'sd0.028115857730702014, 32'sd0.08598730297973389, 32'sd0.06433243053551536, 32'sd-0.08339795499156426, 32'sd-0.21603054121926413, 32'sd-0.0012671134063322934, 32'sd0.0958654958150794, 32'sd0.026574949881666594, 32'sd0.017000992272668696, 32'sd0.1021456490552595, 32'sd0.08474573302926859, 32'sd0.03221254971098638, 32'sd0.0915806848199479, 32'sd0.03760434194005308, 32'sd7.565160944364499e-115, 32'sd-1.557339789222191e-115, 32'sd1.14547356223976e-126, 32'sd1.0061653846616079e-119, 32'sd0.03647993116001749, 32'sd0.03345626728130296, 32'sd0.0683045430224912, 32'sd0.053468557956850224, 32'sd-0.03098018285877315, 32'sd0.002672759050967197, 32'sd0.05170471572523576, 32'sd0.04241737159122286, 32'sd0.015980285042812563, 32'sd-0.04338793774202503, 32'sd0.026433923161172504, 32'sd0.10270101368713563, 32'sd0.031630681696921084, 32'sd0.05313371210976906, 32'sd-0.06848278799690097, 32'sd-0.04893836379052063, 32'sd0.01207744055442899, 32'sd0.026896439214774453, 32'sd0.06887237892444482, 32'sd0.0720440063183322, 32'sd0.08498256640222647, 32'sd0.1089239622025302, 32'sd0.027830197659521657, 32'sd-8.900282114415893e-127, 32'sd3.33180480746178e-121, 32'sd-5.949918460234008e-124, 32'sd-2.355419856808459e-126, 32'sd1.9252981387390084e-120, 32'sd1.9289084039720212e-125, 32'sd0.10555714677732919, 32'sd0.07257768176887394, 32'sd-0.011906815197827304, 32'sd0.04844771765151092, 32'sd0.01319974605529552, 32'sd0.034143478975418064, 32'sd-0.038593419958411895, 32'sd-0.0027885225209208974, 32'sd0.021953146078764862, 32'sd0.09373159864519327, 32'sd0.056118006678772224, 32'sd-0.008618739874656799, 32'sd-0.06551590561586332, 32'sd0.075802480781159, 32'sd0.06031680011993914, 32'sd-0.029329232987698427, 32'sd-0.03440138573299988, 32'sd-0.041684694605891436, 32'sd-0.10989235736943906, 32'sd-0.011813879038216298, 32'sd2.882302756253856e-120, 32'sd2.1844890177116096e-118, 32'sd-1.0544880405810655e-125, 32'sd5.6616048090378586e-123},
        '{32'sd-1.301234907406941e-121, 32'sd-1.3201892181821705e-121, 32'sd3.6578430435522436e-119, 32'sd6.779453060142047e-117, 32'sd2.1114707395290675e-124, 32'sd1.7236648304089828e-125, 32'sd-2.7590572113939745e-120, 32'sd-8.739242904826143e-122, 32'sd7.319257501489618e-117, 32'sd-2.7327440598036436e-116, 32'sd7.040000956158041e-115, 32'sd-8.556897629023046e-127, 32'sd0.02419654322152389, 32'sd0.11389201061231424, 32'sd-0.025447329684156937, 32'sd0.044660815388230565, 32'sd-2.108380477649051e-117, 32'sd9.024746799255338e-121, 32'sd-3.5908879198404425e-115, 32'sd1.392025429388826e-125, 32'sd-6.040360331073348e-121, 32'sd-2.0996019970949635e-127, 32'sd1.0935048520728235e-122, 32'sd3.5441481525571215e-129, 32'sd-2.3295167580786274e-123, 32'sd2.5396988242135725e-117, 32'sd-3.971347695310552e-121, 32'sd-8.024494755054623e-116, 32'sd4.070307770888721e-118, 32'sd-5.205628003438937e-125, 32'sd3.422186535513359e-117, 32'sd3.289678306060463e-116, 32'sd-0.017937117914582065, 32'sd0.01876544684523127, 32'sd0.06341326716011289, 32'sd0.024936542842119432, 32'sd0.07755777477359896, 32'sd0.02826695087398524, 32'sd0.03416505959826575, 32'sd0.08380303106608235, 32'sd0.09837942384484932, 32'sd0.05660645135981885, 32'sd0.0792889380348198, 32'sd0.006700445550980102, 32'sd0.0645904400475951, 32'sd0.07835985376116818, 32'sd0.02978985733691568, 32'sd-0.002969054884058419, 32'sd0.05640407797965238, 32'sd0.10054295641487447, 32'sd0.010635276696695178, 32'sd0.05724827012822466, 32'sd-2.5957834713187935e-115, 32'sd1.4306181641417238e-115, 32'sd1.9022326770098656e-114, 32'sd3.8816055295537027e-118, 32'sd-1.1392967274529057e-119, 32'sd7.871080516294324e-122, 32'sd-0.01111662442267491, 32'sd-0.04702565696571962, 32'sd0.00424158359918692, 32'sd-0.07805735973496353, 32'sd0.03410965188816732, 32'sd0.08616912634884907, 32'sd-0.09097117021048354, 32'sd-0.09791698402623915, 32'sd0.028301137974220188, 32'sd-0.060759264869248084, 32'sd-0.06083752831105797, 32'sd-0.040568876369975845, 32'sd0.07209592014962471, 32'sd0.04598653134164788, 32'sd0.1174157947728046, 32'sd0.13965702940691607, 32'sd0.008061332989217254, 32'sd0.009349674905588367, 32'sd-0.03271145620723866, 32'sd-0.09706905917793442, 32'sd0.014474890076443392, 32'sd0.0069654047310402836, 32'sd0.01767490934217332, 32'sd0.05649689097293773, 32'sd-7.371094097178309e-115, 32'sd9.874962685280048e-117, 32'sd-1.2754474547556028e-116, 32'sd1.4274934005551051e-119, 32'sd-0.02038337000254969, 32'sd0.0852853835861942, 32'sd0.07547535262943855, 32'sd-0.10436131162317831, 32'sd-0.02201802718105613, 32'sd-0.02913739614952896, 32'sd-0.22155838580053283, 32'sd-0.1305863047480233, 32'sd-0.09749654815692765, 32'sd0.03905627785588477, 32'sd0.003952529707783794, 32'sd0.08340861995837766, 32'sd0.13768143289593335, 32'sd0.07913240809484749, 32'sd0.10448114220670292, 32'sd0.057119208757658115, 32'sd0.012757279443057993, 32'sd-0.07658450788130655, 32'sd-0.11355105688264391, 32'sd-0.11187836952245087, 32'sd0.0022569824137020074, 32'sd-0.003228022457991782, 32'sd-0.029446679557388944, 32'sd-0.05701808396262041, 32'sd0.09535725659514589, 32'sd-3.113878589786602e-116, 32'sd2.5474174561831812e-126, 32'sd0.030821786735480403, 32'sd0.0476281071150474, 32'sd-0.06822698343181019, 32'sd-0.027110003542053503, 32'sd-0.05753933476875198, 32'sd-0.012980781618108601, 32'sd-0.022082264487872302, 32'sd-0.04422325315539074, 32'sd0.08987913204020355, 32'sd-0.055972654107333104, 32'sd-0.13313931166577408, 32'sd-0.07369754467403464, 32'sd0.15001165913802025, 32'sd0.08969163519787661, 32'sd0.05770286005324421, 32'sd0.08736345063344941, 32'sd0.1618335532106228, 32'sd0.08275634910856648, 32'sd0.11172593927143143, 32'sd-0.021935582412329617, 32'sd-0.1553863538598747, 32'sd-0.07686623453607756, 32'sd-0.09876062053177406, 32'sd-0.046867217651202504, 32'sd-0.007333251042576449, 32'sd0.03523468391522978, 32'sd0.05230569721391323, 32'sd-4.881649949808468e-127, 32'sd0.022601807698910036, 32'sd-0.050696634186418434, 32'sd0.06868393079359622, 32'sd-0.08312963392525041, 32'sd0.09346448870336616, 32'sd-0.004505237369017174, 32'sd-0.004205466953041034, 32'sd0.08322445078630304, 32'sd0.09677100640564944, 32'sd0.011106186087766855, 32'sd0.03244787557033476, 32'sd-0.06411698194417416, 32'sd-0.1269232766228097, 32'sd-0.17388053227271205, 32'sd-0.04741292276596659, 32'sd0.003536870929483268, 32'sd0.005906155115200797, 32'sd0.10005234439338986, 32'sd0.09069228732613055, 32'sd0.08608956539540617, 32'sd-0.03971517467982642, 32'sd-0.09311683992639098, 32'sd0.10954412918107281, 32'sd0.042484551441842634, 32'sd0.05471150770700494, 32'sd-0.01101146168113253, 32'sd-0.06586804792027151, 32'sd-1.4314695145460683e-118, 32'sd0.0161734907145677, 32'sd0.004882305171905778, 32'sd0.040105250747218005, 32'sd0.02044026285758903, 32'sd0.0534703476611465, 32'sd0.008301900228241902, 32'sd-0.02417571428753528, 32'sd0.1034995060690086, 32'sd0.0930403116426283, 32'sd-0.11631988350170483, 32'sd-0.09991691212517412, 32'sd0.010668268218005079, 32'sd-0.08973491958313899, 32'sd-0.10747717235699085, 32'sd-0.1510626073469719, 32'sd-0.19704959617219592, 32'sd0.06956424450549424, 32'sd0.1630918646750668, 32'sd0.1372270797751123, 32'sd0.06269540953499282, 32'sd0.08910510957694816, 32'sd0.03217232246639724, 32'sd0.014588189480649648, 32'sd0.039953323856976426, 32'sd0.052120179125650264, 32'sd-0.06148662962837978, 32'sd0.04504372282974708, 32'sd0.01159178283458728, 32'sd0.025260597585316902, 32'sd0.08988005734578149, 32'sd0.07483831747351348, 32'sd0.11814580409961016, 32'sd0.09249621772991601, 32'sd0.017293011876611124, 32'sd0.027179437736572682, 32'sd0.06875409288204365, 32'sd-0.0006938016078422791, 32'sd-0.0570405024191929, 32'sd0.06812893944824355, 32'sd0.13242596222451564, 32'sd-0.04523105781580674, 32'sd-0.15019600615249024, 32'sd-0.1823981098523429, 32'sd-0.17407061828181739, 32'sd-0.07658588279939388, 32'sd0.09969759869020514, 32'sd0.15470836644631739, 32'sd0.021952941331194572, 32'sd-0.01001585608763788, 32'sd0.06249313383116168, 32'sd-0.0693838885368964, 32'sd-0.03489331499151537, 32'sd-0.048251781443751814, 32'sd-0.0930970826883585, 32'sd-0.0830621548031874, 32'sd0.01393058089039377, 32'sd0.031913464343540844, 32'sd0.0544658729158023, 32'sd0.07526936261447394, 32'sd0.032634596679662, 32'sd0.07696810783163066, 32'sd0.008959524953827987, 32'sd0.10276623575537054, 32'sd-0.028217949313036457, 32'sd0.07234770623168958, 32'sd0.06393543942792906, 32'sd0.10197958689348754, 32'sd0.057487900084677884, 32'sd-0.06378293982379192, 32'sd-0.24011343705029356, 32'sd-0.3099359343535722, 32'sd-0.18062171361815357, 32'sd0.10348426793121816, 32'sd0.26374346066077986, 32'sd0.15606463907479567, 32'sd0.03958387472505519, 32'sd0.07553005309923042, 32'sd-0.0033876402847972144, 32'sd-0.015956896459144113, 32'sd-0.17682045768113822, 32'sd-0.10234347222548067, 32'sd-0.061518888066599, 32'sd0.0014465583760980914, 32'sd-0.04323431678859336, 32'sd0.03540530844687559, 32'sd-0.0349794173340523, 32'sd0.0053316627376147575, 32'sd0.1465559677993093, 32'sd-0.005199498540238997, 32'sd-0.06176812241880269, 32'sd0.11372936854769672, 32'sd0.11154163640650884, 32'sd0.016617505953506053, 32'sd0.008843808480641598, 32'sd0.10687800015106345, 32'sd0.06522843008639172, 32'sd-0.06520960225240059, 32'sd-0.1298337045127182, 32'sd-0.33551846618465264, 32'sd-0.1844603132296433, 32'sd0.1693060783594839, 32'sd0.2843777568553636, 32'sd0.17703369632984772, 32'sd0.16518127693240559, 32'sd0.061967358885662266, 32'sd-0.11615949343061843, 32'sd-0.06737488425191512, 32'sd-0.10923168143794966, 32'sd0.007064424356518627, 32'sd-0.048949398440124345, 32'sd0.05332485865155048, 32'sd0.052717544623042005, 32'sd-0.046403208968156126, 32'sd0.0799926157491696, 32'sd0.10050135031945101, 32'sd0.01868361296234344, 32'sd-0.05696257627557105, 32'sd-0.05195862819926091, 32'sd0.07232263383002933, 32'sd0.03235221093469006, 32'sd0.003535283293080192, 32'sd0.04970951314374913, 32'sd0.032065066727641894, 32'sd-0.05023178324644163, 32'sd-0.17783790135671218, 32'sd-0.13602834993465568, 32'sd-0.12623503883630988, 32'sd0.005548630463244788, 32'sd0.16486593540030994, 32'sd0.1946480625321643, 32'sd0.11278172105680906, 32'sd0.05308854932692427, 32'sd0.07092077066020439, 32'sd-0.09507916098974087, 32'sd-0.15988070277359, 32'sd-0.15641967070276497, 32'sd-0.013488379688216702, 32'sd-0.08122706546949104, 32'sd-0.0060417759924084125, 32'sd-0.03397325322703125, 32'sd0.05454088933263465, 32'sd0.04248543065747658, 32'sd0.0672099799451484, 32'sd0.025647789207464314, 32'sd-0.07472482980435895, 32'sd-0.024577916062966762, 32'sd0.0437189351899718, 32'sd0.13276625169509057, 32'sd-0.0809805771816341, 32'sd0.08774589029270974, 32'sd0.00392147827006212, 32'sd-0.03101548000645767, 32'sd-0.05050499223737986, 32'sd-0.08396099681096186, 32'sd0.019117532201763543, 32'sd0.027542665391195875, 32'sd0.16389987623381302, 32'sd0.1573678047551775, 32'sd-0.09073897320441177, 32'sd0.05892504430097047, 32'sd-0.05283631880033702, 32'sd-0.041370040337598786, 32'sd-0.08180069424087058, 32'sd0.029731421784150527, 32'sd-0.0027182177041784046, 32'sd-0.030813852994018457, 32'sd0.0012088093618834606, 32'sd0.013235289803907722, 32'sd0.06474360313734835, 32'sd-0.06650905164283759, 32'sd-0.031970279583853574, 32'sd-0.05388760188413382, 32'sd0.09917141565112873, 32'sd-0.0007692433212298233, 32'sd0.005174296469053022, 32'sd-0.05856655921654301, 32'sd0.09835941881929441, 32'sd0.0666149193321224, 32'sd0.05456750328519081, 32'sd-0.04128859139898677, 32'sd-0.016484610620990332, 32'sd0.009400532995324081, 32'sd-0.10539481587786881, 32'sd0.11602616327267869, 32'sd0.09504768886708186, 32'sd0.010529545738054069, 32'sd-0.017696131239497436, 32'sd-0.04785032594781084, 32'sd-0.07875536030164361, 32'sd-0.0202136931441945, 32'sd-0.06634217905937968, 32'sd0.1142382370838649, 32'sd-0.06696997331358595, 32'sd-0.07028481425470186, 32'sd0.028826281166981892, 32'sd-0.008336433634253218, 32'sd-0.011102243472507206, 32'sd0.07463747199136167, 32'sd0.0220498961138814, 32'sd-0.06667308949146843, 32'sd0.006542645424059625, 32'sd0.03461528871981339, 32'sd0.04095505916516433, 32'sd0.04344009462766256, 32'sd0.0852094008656369, 32'sd-0.05231216120179427, 32'sd0.0775981686448371, 32'sd-0.10667582760883221, 32'sd-0.09054624641658748, 32'sd-0.02619838867532626, 32'sd-0.021511463215552605, 32'sd0.004111661163235325, 32'sd0.1271664277180517, 32'sd0.03984438853771527, 32'sd-0.07531077951522638, 32'sd0.03616289250020605, 32'sd0.009593244013250127, 32'sd-0.0008787515250120664, 32'sd-0.080799843119898, 32'sd-0.0959749871908271, 32'sd-0.07701220003988733, 32'sd-0.007805526241471568, 32'sd0.029398267131085818, 32'sd-0.04066921159159943, 32'sd0.05730308378732014, 32'sd-0.04107686515955623, 32'sd-0.14129384786902136, 32'sd0.060445391421990895, 32'sd0.0792606825021833, 32'sd0.02200762102690149, 32'sd-0.07766344792520548, 32'sd-0.04979284470868645, 32'sd0.129117396192402, 32'sd0.10989187137389654, 32'sd0.05779302891548694, 32'sd0.01716338420142279, 32'sd0.02921380700128137, 32'sd0.05263835035921528, 32'sd-0.03562842563949458, 32'sd-0.11829340907522129, 32'sd0.038985702452810446, 32'sd0.049648659594656135, 32'sd-0.0023578259461756955, 32'sd0.0022871472310384026, 32'sd0.0898812822376806, 32'sd0.08865644708627608, 32'sd-0.032112658816472475, 32'sd0.03816351733823735, 32'sd-0.0028461506886693294, 32'sd0.03676373041177224, 32'sd0.07014497287200175, 32'sd-0.015055605581617072, 32'sd0.02343567823474372, 32'sd0.004393706218496335, 32'sd0.07679131258587432, 32'sd0.025665307373642237, 32'sd-0.110127971693363, 32'sd-0.06910169080312582, 32'sd0.01646277550364526, 32'sd0.14269245875111886, 32'sd0.09294796389876725, 32'sd0.13141023281424005, 32'sd0.040894334182397046, 32'sd-0.054198574249688686, 32'sd0.0998697215961593, 32'sd0.08744688318287934, 32'sd-0.020250582727113314, 32'sd-0.09656153337875675, 32'sd-0.07326458574057133, 32'sd0.013684087514761516, 32'sd0.12481486742410412, 32'sd-0.03499924958626444, 32'sd-0.009458068933675552, 32'sd0.04036608799200659, 32'sd-0.10242997841466743, 32'sd0.09307914414477134, 32'sd-0.07613224539094555, 32'sd-0.11982746959354647, 32'sd0.0016888728379723568, 32'sd0.007758147655622774, 32'sd-0.030297968092318165, 32'sd0.005925806656691578, 32'sd-0.05220460658998825, 32'sd-0.008618131166184683, 32'sd-0.10947848928471038, 32'sd-0.1740321610974758, 32'sd0.04185858709728103, 32'sd0.0995034077100811, 32'sd0.11915662869215614, 32'sd0.07181319567367729, 32'sd0.01848509888789417, 32'sd-0.05373873053341145, 32'sd0.07809425144191513, 32'sd0.13463941771248522, 32'sd0.02108615746817515, 32'sd0.00186847765463656, 32'sd-0.09651813534577672, 32'sd-0.06639965946334452, 32'sd0.07323827466557808, 32'sd-0.05539074989967529, 32'sd0.001211640730099517, 32'sd-0.04616329378425767, 32'sd-0.054879629051958076, 32'sd-0.023570694816646413, 32'sd-0.04990374396096231, 32'sd-0.031581873636944265, 32'sd0.022587896913830462, 32'sd2.162332669819092e-116, 32'sd0.03902711420711467, 32'sd0.02449918154750212, 32'sd0.07119556017149009, 32'sd-0.004506238866329782, 32'sd-0.04348910112109668, 32'sd-0.07097484260094739, 32'sd0.16738744956515159, 32'sd0.12933234705145386, 32'sd0.02202188521896352, 32'sd0.03472260436631295, 32'sd-0.05928797006470116, 32'sd0.007490422745744545, 32'sd0.009949336208944873, 32'sd0.08888804780903202, 32'sd0.04460059802558949, 32'sd-0.055006200258592715, 32'sd0.04156227726320748, 32'sd0.030765005122276725, 32'sd-0.03493002362068134, 32'sd-0.06956571366030787, 32'sd-0.06268965462812182, 32'sd0.010380248953735693, 32'sd-0.10175801881311487, 32'sd-0.0740408490913624, 32'sd-0.07495022266864194, 32'sd-0.04909706406205217, 32'sd0.09547492155378959, 32'sd-0.0077140252409563575, 32'sd0.05569870486034097, 32'sd0.032962669644410914, 32'sd0.1214530878398727, 32'sd-0.006223297790631117, 32'sd-0.04442811419825814, 32'sd-0.05853271365085662, 32'sd0.13853419828923388, 32'sd0.13625695777078234, 32'sd0.052856734146328264, 32'sd0.020721554978420754, 32'sd-0.060872797765154085, 32'sd-0.17215140882013205, 32'sd-0.1259226854228315, 32'sd-0.04492298244631273, 32'sd0.012733746039164953, 32'sd-0.0087316414504414, 32'sd-0.06781700844772391, 32'sd0.0751556901096825, 32'sd0.014852140702684534, 32'sd0.033229424134071026, 32'sd0.004770818478910886, 32'sd-0.037102973104221094, 32'sd-0.16993637099651263, 32'sd-0.04799219845360498, 32'sd0.08255623898871656, 32'sd-0.07432796795434672, 32'sd-0.003610135411423899, 32'sd0.021615865335674018, 32'sd-0.028310190383848986, 32'sd-0.05221710355795441, 32'sd0.14266624536445094, 32'sd-0.0745540592340664, 32'sd-0.034957557886825974, 32'sd-0.1266985607119646, 32'sd0.06520507765192408, 32'sd0.01889106020525566, 32'sd0.032908306866193476, 32'sd0.14403649021785414, 32'sd0.04058731562351648, 32'sd-0.25011205628969113, 32'sd-0.10042952771813914, 32'sd-0.02840687921616791, 32'sd0.13829311382835896, 32'sd0.11230766322159587, 32'sd0.0066656249210625, 32'sd-0.06764990101376522, 32'sd-0.05215326662222022, 32'sd-0.06270902401641539, 32'sd-0.05162562594059811, 32'sd-0.027747163779543088, 32'sd-0.09725488566978523, 32'sd-0.04547528302168458, 32'sd-0.01815543769381552, 32'sd-0.10751483515430688, 32'sd-0.016056297394320237, 32'sd-1.1615126248650844e-126, 32'sd0.046024574929966165, 32'sd0.029935860344710963, 32'sd0.06980145280417147, 32'sd0.019700187128748596, 32'sd-0.002748513894136766, 32'sd-0.05228121239600859, 32'sd-0.02574912717851307, 32'sd0.08413896120883115, 32'sd0.033461589578842224, 32'sd0.10485578384923096, 32'sd-0.0268019206836619, 32'sd-0.0653904454679373, 32'sd-0.049839809404705275, 32'sd-0.07878725327555786, 32'sd0.09759520717641407, 32'sd0.011589278376369081, 32'sd-0.06337928884438655, 32'sd-0.03246364133441326, 32'sd0.022845278539318236, 32'sd0.05748883534530698, 32'sd0.049351150504798755, 32'sd-0.11611891105257734, 32'sd0.04605093465511458, 32'sd-0.0208153553961492, 32'sd-0.025158374126814948, 32'sd0.05588511616930484, 32'sd-0.0408328219478117, 32'sd-0.020817922245245618, 32'sd0.04360733670512293, 32'sd0.08952886146523782, 32'sd0.05110561172808959, 32'sd-0.015178674397660661, 32'sd-0.05027007606399993, 32'sd0.03543256803044291, 32'sd0.026021166832439508, 32'sd0.03713901142791503, 32'sd0.09832534870030661, 32'sd0.06383143574422726, 32'sd-0.03304392785176828, 32'sd0.008191069850681302, 32'sd0.026929183112552477, 32'sd0.006231437488178438, 32'sd0.09951823959984278, 32'sd-0.017231441463136935, 32'sd-0.018373497268872434, 32'sd-0.05303669623729451, 32'sd-0.008465549095556702, 32'sd0.012787668911073942, 32'sd0.03331695491397525, 32'sd0.029753357558258576, 32'sd0.03740335327131758, 32'sd-0.07574631820202797, 32'sd0.07126119853562071, 32'sd0.09513814324596842, 32'sd0.02782521883697766, 32'sd-0.004692970375968324, 32'sd-0.061155732222431376, 32'sd0.03897785931096584, 32'sd0.06583361251146821, 32'sd0.042898582341277726, 32'sd0.013472066033900438, 32'sd0.015642030811562135, 32'sd-0.004516002200659402, 32'sd0.14018059355857923, 32'sd0.04557778170821452, 32'sd0.016378247942144264, 32'sd0.033520694592050905, 32'sd0.05826213249469878, 32'sd0.06485146042951037, 32'sd-0.048146793092739545, 32'sd0.08918466801693913, 32'sd0.039457264451948026, 32'sd-0.03731759726565273, 32'sd-0.02921125942589151, 32'sd0.008604261638352931, 32'sd0.003906378039715483, 32'sd-0.015370412008844685, 32'sd-0.09808475040281472, 32'sd-0.12259057028556312, 32'sd-0.010471413552592469, 32'sd-0.0036307987577115495, 32'sd0.006557397959788443, 32'sd-0.018093120934202515, 32'sd-1.949570953877882e-114, 32'sd-0.002600176479722669, 32'sd0.03207058560783643, 32'sd0.052105490971960135, 32'sd0.03210195640838894, 32'sd0.07236914740511566, 32'sd0.0685622729704911, 32'sd0.09776922577044135, 32'sd0.15918859161365614, 32'sd-0.0037079885140393, 32'sd-0.019269099341834336, 32'sd0.059378012057146594, 32'sd-0.06576917771090927, 32'sd-0.11191330072481484, 32'sd-0.022412065570501172, 32'sd-0.006117518305787568, 32'sd-0.029061927788875654, 32'sd-0.10922649786055595, 32'sd-0.007501302135146561, 32'sd-0.020103341422345572, 32'sd-0.05105496041071041, 32'sd0.04366676159985498, 32'sd-0.03929540639290479, 32'sd0.07194556439647215, 32'sd0.04971543554716559, 32'sd-0.09629679989198957, 32'sd0.022361226743718005, 32'sd-3.717434604448293e-119, 32'sd9.26127900375633e-125, 32'sd8.32197390084976e-118, 32'sd0.025893154180379758, 32'sd-0.03418558155010133, 32'sd0.07673165671301722, 32'sd0.09804887606546353, 32'sd-0.08209909178657833, 32'sd-0.018365945596022053, 32'sd-0.03545538730516042, 32'sd0.009780177396533987, 32'sd0.035299249403627914, 32'sd0.03946015782770099, 32'sd-0.08906459902218299, 32'sd-0.07089604342348074, 32'sd-0.031736364608775304, 32'sd-0.1033546656446385, 32'sd-0.029945345298312994, 32'sd-0.05101193119091556, 32'sd-0.07854782426543283, 32'sd0.044495967122616074, 32'sd0.06747982944985086, 32'sd0.03677999482021852, 32'sd-0.057291573322176916, 32'sd-0.04638893126436332, 32'sd-0.07393661230111866, 32'sd-0.012120080670698408, 32'sd0.04508737032235366, 32'sd2.715087841270808e-124, 32'sd-7.226003214604753e-122, 32'sd-1.1797890616858778e-126, 32'sd-0.018315744800942984, 32'sd0.056648165952088506, 32'sd-0.0037023287548768754, 32'sd-0.004948466790123369, 32'sd-0.06661167257259692, 32'sd-0.09798698811532215, 32'sd-0.03226766931012419, 32'sd0.008431177624642619, 32'sd0.04464537129745088, 32'sd-0.04729792897418718, 32'sd-0.1248339141296182, 32'sd-0.08759525034327062, 32'sd-0.12986872358023713, 32'sd-0.10419855581116157, 32'sd-0.054367878845111836, 32'sd0.029935549822893336, 32'sd0.017205434598169696, 32'sd-0.13803247303515281, 32'sd-0.020489158790458473, 32'sd-0.04285393983243698, 32'sd-0.058480327840460485, 32'sd0.08094765855182735, 32'sd-0.02643846808971099, 32'sd-0.009663627925652968, 32'sd-0.017000379342459196, 32'sd6.8578028149414925e-130, 32'sd1.9620143525542446e-122, 32'sd1.4213011602346988e-118, 32'sd-3.7617634908664094e-117, 32'sd0.02293859108457802, 32'sd0.003418223006930136, 32'sd-0.10341902665373524, 32'sd0.05108099536876334, 32'sd-0.0002613121915845099, 32'sd0.11385661959822786, 32'sd0.052347802949609036, 32'sd-0.042871995152202726, 32'sd-0.153755071738178, 32'sd0.09481754098255926, 32'sd-0.0015974471278362994, 32'sd-0.06974132520500646, 32'sd-0.05695737791958518, 32'sd-0.03360494887131511, 32'sd0.13279676727265888, 32'sd-0.05828371795710607, 32'sd-0.1300399219775685, 32'sd-0.08982956685815417, 32'sd-0.14183495214006822, 32'sd-0.13887456233494427, 32'sd0.054898290066397265, 32'sd0.0801072724739272, 32'sd0.04435563081873662, 32'sd-5.274689948526472e-128, 32'sd-6.729662882836487e-124, 32'sd-8.105536657520882e-122, 32'sd-1.1320535529285351e-123, 32'sd8.475353007169941e-117, 32'sd6.889508017510775e-124, 32'sd0.054163984507889146, 32'sd0.032416603399319094, 32'sd0.03750324577490273, 32'sd-0.04834299482053984, 32'sd-0.024166477425073583, 32'sd0.015255642057719633, 32'sd-0.04082351328962801, 32'sd-0.043695047554504145, 32'sd0.054740117157744156, 32'sd-0.015976692182229982, 32'sd-0.04890142815137024, 32'sd0.016282565363024342, 32'sd-0.045209847688443494, 32'sd-0.007189945661606101, 32'sd-0.0029458181008245356, 32'sd0.01940958165942145, 32'sd0.06420171205246486, 32'sd-0.01251983484717372, 32'sd-0.024907428148903045, 32'sd-0.011262132951270442, 32'sd9.730309804459176e-123, 32'sd5.100807233070979e-119, 32'sd-3.5022939834319244e-114, 32'sd1.242443846933822e-117},
        '{32'sd-2.8305786321247644e-117, 32'sd-6.954578517506293e-125, 32'sd9.743441883542399e-122, 32'sd-4.3048705691684965e-121, 32'sd3.910554215257819e-125, 32'sd-3.350479906853389e-123, 32'sd1.9638385510078748e-127, 32'sd3.0012878910012045e-127, 32'sd1.1126407711085365e-127, 32'sd-4.008166373908738e-118, 32'sd3.473318513558867e-127, 32'sd1.8185937759552755e-124, 32'sd-0.011855960507023363, 32'sd-0.011721382681874656, 32'sd-0.01817567925844555, 32'sd0.0022954256837078996, 32'sd1.7934899221310026e-120, 32'sd-1.260190597145556e-115, 32'sd-1.1330843045541984e-115, 32'sd4.380241174557339e-127, 32'sd-7.442544078711054e-116, 32'sd-3.6294934418730415e-123, 32'sd3.43575069822824e-118, 32'sd-2.0244795650061786e-122, 32'sd5.7614703821051875e-117, 32'sd-3.2482999408323503e-124, 32'sd2.254680912348497e-125, 32'sd-3.8990672635111245e-126, 32'sd-3.3303134740396105e-121, 32'sd1.2047074537489934e-118, 32'sd-2.532291699781704e-116, 32'sd2.020310489049299e-117, 32'sd0.03168192024925694, 32'sd0.06418676446040553, 32'sd-0.06322779835659277, 32'sd0.027179409247302454, 32'sd0.05303504020126848, 32'sd-0.06040078601722078, 32'sd0.08515001026163312, 32'sd0.015407671142257157, 32'sd0.01465357912264076, 32'sd-0.05849074436867022, 32'sd0.07471876929787001, 32'sd0.02284230579982396, 32'sd-0.06208629426502188, 32'sd0.06244200225457, 32'sd0.020607593413328178, 32'sd0.004118996721869672, 32'sd0.06885956511932462, 32'sd0.08475472845503432, 32'sd0.058960967927560316, 32'sd0.06095060266009999, 32'sd-3.274534084385783e-121, 32'sd-6.934818993118038e-121, 32'sd-1.0420738387924127e-121, 32'sd2.560330473267251e-118, 32'sd-2.950111095423232e-121, 32'sd-3.699361530831293e-120, 32'sd0.08600799048803412, 32'sd0.08838742924752026, 32'sd0.032592323711602554, 32'sd0.01015902438819096, 32'sd0.00431796104471295, 32'sd-0.05651242856100435, 32'sd-0.01302964405170337, 32'sd-0.021104269286147937, 32'sd0.10475731850170011, 32'sd0.038623677979700705, 32'sd0.007956110032695697, 32'sd-0.019568497708346153, 32'sd-0.1784612175928805, 32'sd-0.17163129085661835, 32'sd-0.11807385276188458, 32'sd0.051903005876648, 32'sd0.02777153967468095, 32'sd0.07818122960581092, 32'sd-0.017936725472474303, 32'sd0.004226559421312187, 32'sd0.09622213927824978, 32'sd-0.004578824621054973, 32'sd0.01995594686561516, 32'sd0.013589254406403597, 32'sd-2.0471864208050447e-124, 32'sd1.0899847197323793e-121, 32'sd-8.865779860529958e-120, 32'sd-3.412635929246258e-114, 32'sd0.11112308852533717, 32'sd0.10601609869064697, 32'sd-0.03602884908193726, 32'sd0.08249827704856942, 32'sd0.015171203810717016, 32'sd0.07870883557263864, 32'sd0.05706013631337836, 32'sd-0.12456067690534438, 32'sd-0.047998648072104196, 32'sd-0.04382577700726175, 32'sd0.030508309069771478, 32'sd-0.13404065276525257, 32'sd-0.10490149806618838, 32'sd-0.03588516049555314, 32'sd-0.07832139619473104, 32'sd0.03293982293190123, 32'sd-0.12244669442656772, 32'sd0.04756496976991551, 32'sd-0.017500337996295447, 32'sd-0.0329924426954327, 32'sd0.012922683945502686, 32'sd-0.039902341548745765, 32'sd-0.018755527017928545, 32'sd-0.06913857817031584, 32'sd-0.015406895933336945, 32'sd2.884325267163265e-124, 32'sd1.854493715003217e-116, 32'sd0.02009763428105314, 32'sd0.01627334457178977, 32'sd0.03924214623391566, 32'sd-0.061130816634123133, 32'sd0.03151049872170903, 32'sd-0.09173302383473256, 32'sd0.015962373186710458, 32'sd-0.028678114910065795, 32'sd-0.08971311084253863, 32'sd-0.07275844425880248, 32'sd-0.02679905875194334, 32'sd-0.09640812852812304, 32'sd-0.1438862355090499, 32'sd-0.04170492809513323, 32'sd-0.06890241553864873, 32'sd0.0289852963247729, 32'sd-0.03440796152173958, 32'sd0.002338059327356709, 32'sd-0.0351006681055551, 32'sd-0.03634177677565204, 32'sd0.056828908019298394, 32'sd-0.012624188750037374, 32'sd-0.07258961559823733, 32'sd-0.04263746369450945, 32'sd0.0682789558061717, 32'sd0.060543455045499975, 32'sd-0.05041487588949982, 32'sd3.4318701070745016e-122, 32'sd0.055795725926174634, 32'sd0.04985764959072256, 32'sd-0.09979312651203281, 32'sd-0.06705248465352898, 32'sd0.03310451727666974, 32'sd-0.02173579486220001, 32'sd-0.024965771208473334, 32'sd0.041963609579017, 32'sd0.0035348964939772264, 32'sd-0.03359638199644282, 32'sd-0.142650075623757, 32'sd-0.07186830578572205, 32'sd-0.08496989544557691, 32'sd0.058421192203072084, 32'sd0.05810967152634362, 32'sd0.06752834427000486, 32'sd0.005686760852402171, 32'sd-0.11563546912902051, 32'sd-0.15610698418547359, 32'sd-0.03651617665018042, 32'sd-0.0870813461290289, 32'sd0.017018653882347013, 32'sd0.14017239051859715, 32'sd-0.0020461605089361116, 32'sd0.02546047859174588, 32'sd0.055629085924128775, 32'sd-0.0012360396703585343, 32'sd-1.0239438907213519e-126, 32'sd0.022384922366569457, 32'sd0.05906168304726586, 32'sd0.044994835248529846, 32'sd0.06965545028686757, 32'sd0.004944649114332697, 32'sd-0.017074294370188564, 32'sd-0.049724992566509064, 32'sd0.07566650098921557, 32'sd-0.030057624742483482, 32'sd0.1112780220541847, 32'sd0.06850470575630734, 32'sd-0.08690212999516304, 32'sd-0.1247532022640691, 32'sd-0.05830146724364924, 32'sd-0.05894412354578568, 32'sd-0.03615443540975277, 32'sd-0.09529905994611153, 32'sd-0.001977143327859697, 32'sd0.05414807542723072, 32'sd0.044291149055460784, 32'sd-0.01586351061001977, 32'sd0.00026348710669421127, 32'sd0.07789396916024437, 32'sd0.11262182060026164, 32'sd-0.056810958156851284, 32'sd-0.009379106205467355, 32'sd0.07784090997298697, 32'sd0.02980998112607695, 32'sd0.01461005443421837, 32'sd0.013200306459619237, 32'sd0.02421484245404192, 32'sd-0.00029859842674927276, 32'sd-0.01078648514223111, 32'sd-0.03632767958542294, 32'sd0.030212490493968618, 32'sd-0.03477829002606513, 32'sd0.10468212729276756, 32'sd0.05058077091691972, 32'sd0.04405003605999084, 32'sd-0.09502285752726866, 32'sd-0.13153072100923352, 32'sd-0.014263892821605572, 32'sd0.04617809316866709, 32'sd0.0284138250628996, 32'sd0.11448781490299315, 32'sd-0.06387722837535467, 32'sd0.10133054039526225, 32'sd0.17913307938301515, 32'sd0.02928308017267868, 32'sd0.15220594389780193, 32'sd0.014013127908306099, 32'sd0.026527873358200345, 32'sd-0.04278652192018169, 32'sd-0.04305988187050207, 32'sd-0.05523331683402815, 32'sd0.05301303271054438, 32'sd0.02289564964094256, 32'sd-0.0702964850344031, 32'sd-0.007036714520463089, 32'sd-0.09906809423351601, 32'sd-0.0014407718019971373, 32'sd-0.01162174166071533, 32'sd-0.013609395835647523, 32'sd-0.019325512947905524, 32'sd0.05979023151363057, 32'sd-0.0472126215346612, 32'sd-0.10728484735891448, 32'sd0.013045581778403495, 32'sd0.08151685957728302, 32'sd0.014429791244257223, 32'sd0.04698921047160536, 32'sd0.08343528914545041, 32'sd0.11685779779026556, 32'sd0.15026529378606698, 32'sd0.15473712152640148, 32'sd0.09119430989383244, 32'sd0.09605132921660378, 32'sd0.054783085272965465, 32'sd0.09402074275664066, 32'sd0.09711947989917616, 32'sd0.034258001533127656, 32'sd0.015107781233251549, 32'sd0.040625296158554806, 32'sd0.10655356651137836, 32'sd-0.01639116531071647, 32'sd0.08004678490522248, 32'sd-0.08846153389036672, 32'sd-0.026144091518405153, 32'sd-0.06532866825847518, 32'sd-0.055602331418216286, 32'sd-0.039017045895333086, 32'sd-0.08224584446587055, 32'sd-0.04063061916830278, 32'sd-0.023564914469581935, 32'sd0.03578528877963677, 32'sd-0.05805902100833006, 32'sd-0.04455396881616435, 32'sd-0.15171530607249448, 32'sd-0.12729254532596662, 32'sd0.11123194206335842, 32'sd0.013614291212821981, 32'sd0.16722818398670924, 32'sd-0.053830330020577126, 32'sd0.028341709389729096, 32'sd0.055222144959970416, 32'sd0.05316156694506695, 32'sd0.03387372818396316, 32'sd0.13566117048673298, 32'sd0.07112610645531647, 32'sd0.02623712425672547, 32'sd-0.0380031472538485, 32'sd0.03340431470382849, 32'sd0.05955187943352371, 32'sd0.09696227601428876, 32'sd0.10700827769822671, 32'sd0.012120034520091565, 32'sd0.008543892768791193, 32'sd-0.05075686628928084, 32'sd-0.13019289035247103, 32'sd-0.055231148589345254, 32'sd0.04474511308445045, 32'sd-0.006121307755633353, 32'sd-0.09992682890292845, 32'sd-0.1427436525342623, 32'sd-0.15755661048944153, 32'sd-0.19166950634870572, 32'sd-0.056120797391001495, 32'sd-0.057720629093326495, 32'sd-0.03671588691664483, 32'sd-0.0876612287044685, 32'sd-0.19218031557118354, 32'sd0.00603773017402187, 32'sd0.04072117993075978, 32'sd0.12775371878422104, 32'sd0.025250195003501227, 32'sd0.04938525267042993, 32'sd0.09073176699125099, 32'sd0.05633530602395125, 32'sd-0.01535866014585016, 32'sd0.09180534690507326, 32'sd0.02368190366116781, 32'sd0.01594330814567886, 32'sd-0.052508561750578484, 32'sd-0.09629783393016529, 32'sd0.1001732803378876, 32'sd0.01265312085605902, 32'sd-0.07715685654942796, 32'sd-0.09191099686390766, 32'sd-0.023759561465833336, 32'sd-0.0345861300274217, 32'sd-0.06089458312577254, 32'sd-0.20439216799113416, 32'sd-0.15053271423807923, 32'sd0.009745487080016003, 32'sd-0.11604488724120401, 32'sd-0.19704890285036766, 32'sd-0.14914214917606536, 32'sd-0.15863290211212444, 32'sd-0.24254507454671229, 32'sd-0.1000478298685434, 32'sd-0.05450848110062674, 32'sd-0.1298805164430727, 32'sd-0.05672875334711284, 32'sd-0.018316667474169903, 32'sd0.022578580176886544, 32'sd-0.03865429986257474, 32'sd0.05522273453195924, 32'sd0.02507653063549432, 32'sd0.014200594468160068, 32'sd-0.01975531416431717, 32'sd-0.07559249602612374, 32'sd-0.04275217777820408, 32'sd-0.01679230090721523, 32'sd-0.04174268580454386, 32'sd-0.029849661942489458, 32'sd-0.09848394157540902, 32'sd-0.03774565182770124, 32'sd-0.05382725416667465, 32'sd-0.029766749942774094, 32'sd-0.09841864365588071, 32'sd-0.03537959942902661, 32'sd0.13333779531262777, 32'sd-0.04485122751944061, 32'sd-0.18399617675282817, 32'sd-0.21284685716956864, 32'sd-0.07475911352690004, 32'sd-0.20404451383934938, 32'sd-0.1437667677206585, 32'sd-0.1387161983790298, 32'sd-0.014411712074521814, 32'sd0.033547652491158285, 32'sd-0.057056377034765876, 32'sd-0.19185728366723523, 32'sd-0.14574604090231294, 32'sd0.04058073125680159, 32'sd0.03927535167482415, 32'sd0.030659438549080098, 32'sd-0.025665242079590825, 32'sd-0.08160913038865092, 32'sd-0.023534485033143853, 32'sd0.02891091052159565, 32'sd0.03425001457657709, 32'sd0.007677016233172979, 32'sd-0.07784590563552739, 32'sd0.05948307998310484, 32'sd-0.02850303576802166, 32'sd-0.08561289383714268, 32'sd-0.013582553195105, 32'sd-0.08747967761415881, 32'sd0.10945741948053066, 32'sd-0.018306049166606768, 32'sd-0.07971883542255627, 32'sd-0.1251754996054203, 32'sd-0.07056480069464668, 32'sd-0.1504549144577212, 32'sd-0.10487919669653431, 32'sd-0.08196707882997042, 32'sd-0.07778514158730696, 32'sd0.09311227293229941, 32'sd-0.02389923852904497, 32'sd0.02440348294401694, 32'sd-0.15368818225766812, 32'sd0.019962930869351726, 32'sd0.0708108395876402, 32'sd-0.0142908759067199, 32'sd-0.03735919052290351, 32'sd-0.004340296939365285, 32'sd0.12948131071598915, 32'sd-0.07093423399445624, 32'sd-0.0723976898055174, 32'sd0.05242226385276257, 32'sd0.12033651578625473, 32'sd0.035116376248629184, 32'sd-0.02687909310580883, 32'sd-0.09954454680796639, 32'sd-0.1540607737467008, 32'sd-0.08716534375179524, 32'sd0.09344352724514528, 32'sd-0.04070037518226952, 32'sd-0.09858578688176384, 32'sd-0.06304820915329525, 32'sd-0.07254973649318949, 32'sd-0.1545293126293037, 32'sd-0.11505405974247114, 32'sd-0.09405221546848326, 32'sd0.010090913664124478, 32'sd0.15703973407790986, 32'sd0.23644978624738125, 32'sd-0.012170525287512982, 32'sd-0.08150966238274006, 32'sd0.010150437332551773, 32'sd0.13164860895170002, 32'sd0.008671722421383013, 32'sd-0.11211556940798925, 32'sd-0.06042265572385482, 32'sd0.07326999003398406, 32'sd-0.033907354223163086, 32'sd-0.004568968812416214, 32'sd0.05007671280757906, 32'sd0.02313807257146131, 32'sd0.13618913401510718, 32'sd0.005987203589480702, 32'sd-0.002676459774578021, 32'sd-3.886991921451998e-05, 32'sd0.02967876125678235, 32'sd-0.051078486414652506, 32'sd-0.04721260392448711, 32'sd-0.06289897142629054, 32'sd-0.05577488200547267, 32'sd-0.10127357302209833, 32'sd-0.20487022963404553, 32'sd-0.18536766877144314, 32'sd-0.05187708617990208, 32'sd-0.06602033806162932, 32'sd0.09449477713900976, 32'sd0.17560888863153357, 32'sd-0.07343633019472708, 32'sd-0.11921095794944533, 32'sd0.027751082938154977, 32'sd0.026256472856616933, 32'sd-0.028887063591758768, 32'sd-0.03419095104178184, 32'sd-0.10389912580006108, 32'sd-0.06815805289093115, 32'sd-0.006629570880288324, 32'sd-0.08292290301680734, 32'sd-0.07044457034422928, 32'sd-0.09697586925803049, 32'sd0.035533008287325175, 32'sd0.105188874562213, 32'sd0.03271705222331111, 32'sd0.034767553431330096, 32'sd0.11709808276932994, 32'sd0.026420493328484927, 32'sd-0.07218714225795117, 32'sd-0.11998476429797235, 32'sd-0.10251608579385815, 32'sd-0.027990148501132434, 32'sd0.013959842230426478, 32'sd-0.19180308334385893, 32'sd0.04263290756689357, 32'sd0.09389097117030547, 32'sd0.08205679609299056, 32'sd0.19400936847817907, 32'sd0.045037922233727504, 32'sd-0.07257665267062097, 32'sd0.07265235419145841, 32'sd6.863952178805175e-118, 32'sd-0.014194110077261082, 32'sd-0.020953722817614588, 32'sd-0.08682788740705746, 32'sd-0.03747899981701976, 32'sd-0.0653014743499299, 32'sd-0.0725963209199962, 32'sd-0.10541163195092651, 32'sd-0.03618410988286211, 32'sd-0.07907206641002658, 32'sd-0.1539262537724354, 32'sd-0.03332469021338955, 32'sd-0.09067353997328745, 32'sd-0.0030130046613564923, 32'sd-0.149577224424685, 32'sd-0.1617649352095027, 32'sd-0.10274233523305634, 32'sd-0.055967350677347746, 32'sd-0.0595614345616347, 32'sd0.025039580331960094, 32'sd0.10044732075937632, 32'sd0.043303281087928025, 32'sd0.10055155405531577, 32'sd0.13600099169695082, 32'sd0.16664576880331108, 32'sd-0.005242786079984858, 32'sd0.06587675311565244, 32'sd-0.05156839817677852, 32'sd0.02632020733679763, 32'sd-0.016393148926369963, 32'sd0.005688717549394965, 32'sd0.002527747571655642, 32'sd0.049189812683665346, 32'sd0.006089786650396714, 32'sd-0.1644201485098171, 32'sd-0.14766192888468047, 32'sd-0.08997322345633497, 32'sd-0.23950802496881102, 32'sd-0.1374221530819711, 32'sd-0.14400394569326672, 32'sd-0.1007222717091425, 32'sd-0.0006826074539164258, 32'sd-0.2096573486948282, 32'sd-0.28392987697919203, 32'sd-0.0156438157402997, 32'sd-0.055959610785865595, 32'sd-0.017719479854457997, 32'sd0.02058723116869843, 32'sd0.09043482225156602, 32'sd-0.0495893321509339, 32'sd0.02481623962121427, 32'sd0.023500717707103522, 32'sd-0.0870863323666564, 32'sd0.04828462824807425, 32'sd0.04676797116301554, 32'sd-0.05628481663888952, 32'sd0.056311051242242546, 32'sd0.046413418244883764, 32'sd-0.06626123145553553, 32'sd0.0160475720861034, 32'sd-0.10022806175475657, 32'sd-0.017103161218331723, 32'sd-0.05478822205404969, 32'sd-0.08967218189626167, 32'sd-0.14276975539950124, 32'sd-0.18584360602114985, 32'sd-0.2395991528110678, 32'sd-0.2596688938573817, 32'sd-0.21810138155156553, 32'sd-0.04294595267116983, 32'sd-0.07345385220921609, 32'sd-0.1771031056555152, 32'sd-0.1083558446386377, 32'sd-0.06732706315227256, 32'sd0.07026838736500836, 32'sd0.06616424479935805, 32'sd0.17106814480314758, 32'sd-0.03426612665676455, 32'sd-0.03168506284101312, 32'sd0.05851265257617841, 32'sd0.039441415624550384, 32'sd-0.0034970417382156316, 32'sd0.05760755565245056, 32'sd-0.04330569985846195, 32'sd1.1305699280416377e-126, 32'sd0.01858485655175501, 32'sd-0.00785648591622771, 32'sd-0.05674997359583143, 32'sd0.0775585584040424, 32'sd0.007355553016333943, 32'sd0.002814610369376449, 32'sd-0.06777604423756055, 32'sd-0.003460874803051127, 32'sd-0.12528333796908867, 32'sd-0.12326593595361465, 32'sd-0.20104581791184656, 32'sd-0.1878638183037605, 32'sd-0.0726769697898964, 32'sd-0.06259928997064541, 32'sd-0.13812529540983234, 32'sd0.018972558884040217, 32'sd0.04635220570766192, 32'sd0.026117627869091033, 32'sd0.12589320710007254, 32'sd0.13695327674419508, 32'sd-0.0047912946819020545, 32'sd-0.013540543901397, 32'sd0.009633442093272559, 32'sd0.13388422866531613, 32'sd-0.029094999875697913, 32'sd0.03280867296137233, 32'sd0.07385551492313533, 32'sd0.04208087920783882, 32'sd0.05722943951677545, 32'sd0.080626037418798, 32'sd0.010020021211235549, 32'sd0.0530600377817826, 32'sd0.06312699865703411, 32'sd-0.06028301610507681, 32'sd0.024045357047578236, 32'sd0.11987231752060065, 32'sd0.06409926504029972, 32'sd-0.09705315224290045, 32'sd0.11598603467905998, 32'sd-0.004544181507026561, 32'sd0.018985472109060916, 32'sd-0.01734853209940978, 32'sd0.0657854563108093, 32'sd0.0822464743431196, 32'sd-0.08095306912831819, 32'sd0.11120752806850366, 32'sd0.038160052016296526, 32'sd0.06107802171911753, 32'sd-0.02604328868267845, 32'sd0.020987425791942446, 32'sd-0.0143942159192854, 32'sd0.035738741648846155, 32'sd-0.1111373973148194, 32'sd0.07341942475817764, 32'sd0.022663866313672957, 32'sd0.09200070941601153, 32'sd0.06670167302676465, 32'sd0.07631172612262448, 32'sd0.08946294100546885, 32'sd-0.04218440188541717, 32'sd0.13937807606142544, 32'sd0.08179610768934015, 32'sd0.050044676916020964, 32'sd0.038989831547409703, 32'sd0.006050279621832077, 32'sd0.04846507026141364, 32'sd0.1297510861882551, 32'sd-0.04722359100681894, 32'sd0.05108005127306201, 32'sd-0.033579169127449945, 32'sd0.012700435117027325, 32'sd-0.025721451131863724, 32'sd0.05265985654224162, 32'sd0.032565563800368985, 32'sd0.08812175649364519, 32'sd0.10603572328010946, 32'sd0.013030095576257771, 32'sd0.03302143236832143, 32'sd0.018037081752955635, 32'sd-0.12123212338819979, 32'sd-0.14860856444029383, 32'sd-0.0214054459530561, 32'sd0.06466770005214134, 32'sd-3.201136145475745e-121, 32'sd0.028337714501950377, 32'sd-0.06503680977516652, 32'sd-0.0017863442114039775, 32'sd0.011841095471398186, 32'sd0.0852007810956584, 32'sd-0.027506911224981362, 32'sd0.028869432871674677, 32'sd-0.04568814058030643, 32'sd0.12311255678574934, 32'sd0.07783175766717108, 32'sd0.01834197883925749, 32'sd-0.04334084924602415, 32'sd-0.019250385010135134, 32'sd0.04530349460314113, 32'sd0.05305458078406667, 32'sd0.1554862967749139, 32'sd0.08097650976617089, 32'sd-0.1401075098439156, 32'sd-0.1293665572312889, 32'sd-0.06115106913796901, 32'sd0.020183095201163827, 32'sd0.030608104786631465, 32'sd-0.06145192881670707, 32'sd-0.020584007710902862, 32'sd0.035360939656058944, 32'sd-0.08299775662261229, 32'sd1.791943804669301e-114, 32'sd-3.554346915417648e-119, 32'sd-1.0317568290705167e-119, 32'sd-0.010792515102826222, 32'sd0.04012417366936665, 32'sd0.021805886008160406, 32'sd0.019139525382628177, 32'sd0.023753609629070076, 32'sd-0.0010049629295968642, 32'sd-0.016518929205336198, 32'sd0.041838780920129943, 32'sd-0.07138705970690827, 32'sd-0.015666380016648083, 32'sd-0.05723992050539396, 32'sd0.000803065078903178, 32'sd0.02598536128092204, 32'sd0.020136497062778185, 32'sd-0.05302862692735251, 32'sd0.08628243808494562, 32'sd-0.04193672350909738, 32'sd-0.1598716875660703, 32'sd-0.04875590024680989, 32'sd0.044368184049938, 32'sd-0.05983685678134398, 32'sd-0.1033834007678296, 32'sd0.0010710248069025975, 32'sd0.07164501644981128, 32'sd0.009978662563467702, 32'sd-2.568642427502078e-121, 32'sd9.19364665920665e-124, 32'sd9.573561068101052e-119, 32'sd0.057505194945491264, 32'sd-0.01980869164474648, 32'sd0.0331535296361127, 32'sd-0.03831477907265942, 32'sd-0.03874013585853568, 32'sd0.0033433975405329037, 32'sd0.08821287714973317, 32'sd0.03118068484778069, 32'sd-0.013215629218132805, 32'sd-0.009858019627844725, 32'sd0.008324740255835412, 32'sd0.05482409349891188, 32'sd0.042862586207135615, 32'sd0.07253027910783852, 32'sd-0.045966376679903984, 32'sd-0.030184254492849387, 32'sd0.018742274469543647, 32'sd0.06545223269560634, 32'sd0.05787280932872885, 32'sd0.03959686145023106, 32'sd0.005803968621518142, 32'sd-0.14930870782799444, 32'sd-0.013161096646641161, 32'sd0.03276409024989066, 32'sd0.028139071496301894, 32'sd5.498039199718548e-119, 32'sd2.794460891348377e-119, 32'sd5.262577924258268e-118, 32'sd-1.2241346447401446e-116, 32'sd0.08204619103585979, 32'sd-0.07241195715988509, 32'sd-0.017747172732363328, 32'sd-0.0583903173084532, 32'sd-0.021302183791125515, 32'sd-0.13616202781603337, 32'sd-0.05410994847297444, 32'sd0.019962269300803918, 32'sd0.03929634734042255, 32'sd-0.07756236866949393, 32'sd-0.04614156087942834, 32'sd-0.008244528121516536, 32'sd-0.0017179945926410073, 32'sd-0.11177800926719852, 32'sd0.02895820854716888, 32'sd0.05136837491582511, 32'sd0.024932542461458967, 32'sd-0.058466749092641726, 32'sd0.02729752811137576, 32'sd-0.11058236259951959, 32'sd-0.005274198392146075, 32'sd0.026036077843200833, 32'sd0.05447443272064671, 32'sd-4.870901353715272e-121, 32'sd-8.619874287124936e-119, 32'sd-8.667146538125154e-121, 32'sd-5.452681151898624e-126, 32'sd3.942252081899293e-129, 32'sd-3.239780545644096e-121, 32'sd0.09164082859297602, 32'sd0.07053683402945969, 32'sd0.03142056103110519, 32'sd0.013065907674948625, 32'sd-0.001766152925181976, 32'sd0.023786095823692188, 32'sd0.007872567684914178, 32'sd0.05416408512393782, 32'sd0.05285882987629375, 32'sd0.00014244354866896298, 32'sd-0.07561850240958451, 32'sd0.05747860442648717, 32'sd-0.004629380085812346, 32'sd-0.016786525216323556, 32'sd0.007674019374247939, 32'sd-0.04123648949560787, 32'sd0.028811611555399675, 32'sd-0.025064549116870734, 32'sd-0.10274642998154566, 32'sd0.07373190507890034, 32'sd-1.8189153971892786e-117, 32'sd-5.813758430303762e-126, 32'sd-1.8814063074689888e-122, 32'sd-2.8824214275379375e-124},
        '{32'sd6.786855388706412e-123, 32'sd1.430096698225036e-116, 32'sd-2.288209980949085e-115, 32'sd4.346013637621439e-123, 32'sd-1.268581852084597e-122, 32'sd-3.859769074387711e-125, 32'sd5.782476987805661e-127, 32'sd1.5402124042925615e-115, 32'sd1.4926777965923237e-127, 32'sd8.574262629363782e-127, 32'sd-1.0133250685658237e-115, 32'sd2.514696984001712e-119, 32'sd0.010122813816647602, 32'sd-0.07149981181931019, 32'sd-0.013965143372469206, 32'sd-0.023007183575485434, 32'sd2.510955916449098e-126, 32'sd-5.261980445532858e-118, 32'sd-4.022929497772973e-123, 32'sd3.0875906150192982e-115, 32'sd3.788925831713331e-122, 32'sd1.0021630198112888e-119, 32'sd8.517956273311381e-117, 32'sd-1.0624019290903499e-121, 32'sd1.0385085923525017e-123, 32'sd1.8005343396825494e-123, 32'sd3.3650569009343364e-120, 32'sd2.5637069952619405e-114, 32'sd1.3400414366938915e-116, 32'sd-1.2135234910133097e-115, 32'sd-5.426174164650551e-123, 32'sd1.1019097162992581e-121, 32'sd0.0476554571554093, 32'sd0.0640631323277492, 32'sd0.0381162610010756, 32'sd0.010730658642161025, 32'sd0.09824482406650935, 32'sd0.065450457735608, 32'sd-0.03216802319292027, 32'sd0.08226867120931099, 32'sd0.02236863095521316, 32'sd-0.03829428990995865, 32'sd0.03307083005242918, 32'sd0.08089594571419348, 32'sd0.02518496380712078, 32'sd-0.010907749327849247, 32'sd0.05675534291348675, 32'sd0.02385365001499255, 32'sd0.06878369039762981, 32'sd0.06611532121396603, 32'sd-0.025264595969789295, 32'sd0.02018847031163666, 32'sd-6.807259920003558e-120, 32'sd6.847673653471731e-124, 32'sd-1.6397630734295954e-124, 32'sd2.1784369445335643e-119, 32'sd3.603230316524803e-119, 32'sd7.424984122515955e-115, 32'sd-0.01085498929741223, 32'sd-0.01507335541313462, 32'sd0.011435577575779109, 32'sd-0.015488084897354164, 32'sd0.025279922351520722, 32'sd0.007378181161434078, 32'sd-0.04012770025665326, 32'sd-0.10254403351106112, 32'sd0.00780034506360782, 32'sd-0.04238268545831855, 32'sd0.0486398736486804, 32'sd0.014139796926045367, 32'sd0.037834906774990865, 32'sd-0.048668432723935166, 32'sd-0.12412797145287106, 32'sd-0.028224222752981247, 32'sd0.010433265362981047, 32'sd0.02298068648146877, 32'sd-0.057641234884276596, 32'sd0.12466232623412511, 32'sd-0.011578821176215172, 32'sd0.099393619692312, 32'sd0.030211868951033755, 32'sd-0.017560221473883104, 32'sd1.8317669163681057e-127, 32'sd9.936317662792719e-125, 32'sd6.925991203000479e-117, 32'sd-3.453108231333495e-118, 32'sd-0.020873953648824575, 32'sd-0.04084516234595973, 32'sd-0.0839560382492172, 32'sd0.018301140643500795, 32'sd-0.022551378876269425, 32'sd-0.11426442959983123, 32'sd0.06486150635563498, 32'sd-0.004149638814594299, 32'sd-0.06490149134787476, 32'sd0.009723837385039307, 32'sd-0.031744801253913976, 32'sd0.05280099358567453, 32'sd-0.02107025218467237, 32'sd-0.017380882459084188, 32'sd0.0040947705313479806, 32'sd-0.1267083387320252, 32'sd-0.16345136753204925, 32'sd-0.12283231265657335, 32'sd-0.1901630993194442, 32'sd-0.04004012356018303, 32'sd-0.05862988947566287, 32'sd0.06527356372953674, 32'sd-0.031124505511130114, 32'sd-0.004734258751196493, 32'sd-0.009780064231679526, 32'sd1.253507021283253e-118, 32'sd1.1872346457819095e-127, 32'sd0.008204190186526327, 32'sd-0.0016907850128717475, 32'sd-0.0834413097328133, 32'sd0.026613994743910387, 32'sd-0.048595996669759535, 32'sd0.02158419430269815, 32'sd-0.00551181314886011, 32'sd-0.0524081448071729, 32'sd-0.06082150521859154, 32'sd0.08595870847245934, 32'sd-0.0048498916862646175, 32'sd0.10972895411982121, 32'sd0.12118033184951545, 32'sd0.11985403036054086, 32'sd-0.04050718273185787, 32'sd-0.0802130079848741, 32'sd-0.08017393318766912, 32'sd-0.04968214322647351, 32'sd0.025961166695996293, 32'sd0.11378298978487777, 32'sd-0.04493678058893193, 32'sd0.0035410269678170696, 32'sd-0.12104761026745452, 32'sd0.04499068775318351, 32'sd0.027908587978051482, 32'sd0.057079185859998, 32'sd-0.011620703915080455, 32'sd1.616701683327917e-125, 32'sd-0.021274937634249428, 32'sd0.04272024209707586, 32'sd-0.03688049663556611, 32'sd0.02124752166915722, 32'sd0.01278426305503142, 32'sd0.0686204772310265, 32'sd0.058504206332765006, 32'sd0.013741279468288466, 32'sd-0.08244359767832032, 32'sd-0.01171490575352822, 32'sd-0.07675262715333013, 32'sd0.10722568475597183, 32'sd0.07167446235206247, 32'sd-0.10301361574235059, 32'sd-0.008875043220774825, 32'sd0.006554905356744429, 32'sd-0.05852604786616362, 32'sd-0.08268732920756038, 32'sd-0.05554464290419977, 32'sd-0.12051225880439981, 32'sd-0.05805019759548999, 32'sd-0.0008281534170321266, 32'sd0.034419339095412185, 32'sd-0.10502413244086378, 32'sd-0.03754119464985884, 32'sd0.0031322463979348856, 32'sd-0.0055434136977175995, 32'sd3.0449610515314262e-121, 32'sd0.03253981129041678, 32'sd-0.002105685983400086, 32'sd-0.1242774892949984, 32'sd-0.0012328708792812256, 32'sd-0.05334416732978792, 32'sd0.03161493311984678, 32'sd0.08464816951579864, 32'sd0.013331590254653976, 32'sd-0.061447030333319365, 32'sd-0.09292245786287176, 32'sd-0.05718301938628292, 32'sd-0.05658287735457321, 32'sd-0.05406178730219367, 32'sd0.04371013308478994, 32'sd0.05503705094087104, 32'sd0.05327756809178911, 32'sd-0.04625811256767851, 32'sd-0.02185435812700046, 32'sd-0.00734727967641047, 32'sd0.00866569809089768, 32'sd0.013264755500259849, 32'sd0.03412237461628468, 32'sd-0.07652183288158937, 32'sd-0.17072726731590995, 32'sd-0.14820251048661714, 32'sd0.10294579975797559, 32'sd-0.0017101741263492714, 32'sd0.020932608183029434, 32'sd0.01596477390039271, 32'sd-0.08720366232640187, 32'sd0.07310533207685356, 32'sd0.01872676215716174, 32'sd-0.06378879122718747, 32'sd-0.013844871105382876, 32'sd-0.07750184337923235, 32'sd-0.027571475605986336, 32'sd-0.08690107793113477, 32'sd-0.10763310429447631, 32'sd-0.020854238779229057, 32'sd-0.0923544873037395, 32'sd-0.0552892278222588, 32'sd0.06672364405731103, 32'sd0.15579268151975048, 32'sd0.04187061217608983, 32'sd-0.021023972271007843, 32'sd-0.027389301731822656, 32'sd-0.11299059216785469, 32'sd-0.07694825006140968, 32'sd0.041898950278039374, 32'sd-0.011824440352683603, 32'sd-0.09003263657099438, 32'sd-0.1691854087066896, 32'sd-0.13086774006179794, 32'sd-0.038176665467940366, 32'sd-0.02213289498308603, 32'sd-0.02099932474057831, 32'sd0.05618777004282555, 32'sd-0.03417900059650044, 32'sd-0.07280882787614966, 32'sd0.08849137441880772, 32'sd-0.08539452116665566, 32'sd-0.059349390564217626, 32'sd-0.05454524759685151, 32'sd-0.060605853489896694, 32'sd-0.0803086328540793, 32'sd-0.12988163299468233, 32'sd-0.08880939901030604, 32'sd-0.07164532253447084, 32'sd-0.12880438082183457, 32'sd-0.032479362919185975, 32'sd-0.06251756870871038, 32'sd-0.11077266077549403, 32'sd-0.03605654717048937, 32'sd0.062405017382544406, 32'sd-0.043758979664079836, 32'sd-0.03278456123918408, 32'sd0.06262452656249017, 32'sd-0.046148115605358246, 32'sd-0.16869120723825565, 32'sd-0.18957014267894884, 32'sd-0.0357781999408815, 32'sd0.03911831631681599, 32'sd-0.002132054723580903, 32'sd0.09417505763676064, 32'sd-0.01527119591291948, 32'sd-0.09696495123269301, 32'sd-0.012291793211885185, 32'sd-0.05246976717026951, 32'sd-0.16674129285625613, 32'sd-0.06820003755713494, 32'sd-0.07075741664236626, 32'sd-0.015348058096716959, 32'sd0.01262759257045037, 32'sd0.04252275543436608, 32'sd-0.02118554236461988, 32'sd-0.08224518538466725, 32'sd-0.06034054974084421, 32'sd-0.09121859719848666, 32'sd-0.050342224232186185, 32'sd0.07234475599480773, 32'sd0.11132974421444189, 32'sd-0.10245716003960047, 32'sd-0.02487835776528925, 32'sd-0.06392556982842235, 32'sd-0.011521618457691073, 32'sd-0.12901895045825482, 32'sd0.0010176273071855584, 32'sd0.039759737313419384, 32'sd-0.05392161680117097, 32'sd-0.04936137459987185, 32'sd-0.024617921208619872, 32'sd-0.013044591950936059, 32'sd-0.0013099198095413188, 32'sd-0.03202151825459122, 32'sd0.01789655596609336, 32'sd-0.024055361906186384, 32'sd-0.18485573933178623, 32'sd-0.22919041986989794, 32'sd0.007697033854757775, 32'sd-0.01690749783280672, 32'sd0.1339968966089032, 32'sd0.06521739527202142, 32'sd0.04505314011483015, 32'sd0.03051241049194369, 32'sd-0.10248969115799615, 32'sd0.0342147383571332, 32'sd-0.17038739760431498, 32'sd-0.046072143663138554, 32'sd0.06635235747091836, 32'sd0.11249807557815727, 32'sd-0.013681238304692927, 32'sd-0.1294924108089704, 32'sd-0.23743640925694326, 32'sd-0.086961523090135, 32'sd-0.13269387352480333, 32'sd-0.009295175372771294, 32'sd-0.1757960431533713, 32'sd-0.04179727333632416, 32'sd-0.016711237360789975, 32'sd0.03879838447341166, 32'sd0.07299344657297026, 32'sd0.032741585644871396, 32'sd-0.05023055346362203, 32'sd-0.08888581021356715, 32'sd-0.1573650827977609, 32'sd-0.1337823299400177, 32'sd0.06476137757599061, 32'sd0.08905619833020084, 32'sd0.04725119814818222, 32'sd0.028085044768722343, 32'sd0.10167048017439956, 32'sd-0.026758097228074443, 32'sd0.06761394748874658, 32'sd0.014040485443485955, 32'sd-0.17822137353975534, 32'sd-0.03542116770562462, 32'sd0.10661330308953297, 32'sd0.19593548734458302, 32'sd0.10362576121557099, 32'sd0.0005617086584171587, 32'sd-0.06739218254185758, 32'sd-0.0721453404036407, 32'sd-0.11052789632303288, 32'sd-0.16828789972712152, 32'sd-0.02833407267404102, 32'sd0.005055407322430092, 32'sd0.07500359447644908, 32'sd-0.020127412731152924, 32'sd-0.09625767781250053, 32'sd-0.01941579114042517, 32'sd-0.07841610356081168, 32'sd0.00407926024127069, 32'sd-0.06075947751039878, 32'sd-0.10639093251664487, 32'sd-0.041772863793459535, 32'sd0.05264929474454605, 32'sd0.09307533110633544, 32'sd-0.051049247080584115, 32'sd0.005965487233875887, 32'sd-0.1375496295237458, 32'sd-0.10586920652636973, 32'sd-0.012487579815380305, 32'sd0.007132427860125101, 32'sd0.08162869663187941, 32'sd0.09598801146540234, 32'sd0.19066355080336136, 32'sd0.060621909040494464, 32'sd0.04040577425466986, 32'sd-0.03771108271785066, 32'sd-0.06159526327250588, 32'sd-0.12163730631727405, 32'sd-0.020948652834046, 32'sd0.005983609852343829, 32'sd0.010913589492463358, 32'sd0.07477791129975407, 32'sd-0.019918300110420877, 32'sd-0.011124674114945726, 32'sd0.01324608185083033, 32'sd-0.024431637245334318, 32'sd-0.010063401789675939, 32'sd-0.12223486311138315, 32'sd0.03189306770557398, 32'sd-0.007240834456466445, 32'sd0.03711179522798892, 32'sd0.04967394795661941, 32'sd-0.038224600425656494, 32'sd-0.04291605138399471, 32'sd-0.15314711339221762, 32'sd-0.029770240355016055, 32'sd0.08037333632852883, 32'sd0.03501768418871414, 32'sd0.036218705260149794, 32'sd0.12127484342640565, 32'sd0.14878178210128443, 32'sd0.11724807258966767, 32'sd-0.012179972348298393, 32'sd-0.03455817889179121, 32'sd-0.1056583818940511, 32'sd-0.00023827929097897614, 32'sd-0.11109227976804158, 32'sd-0.10358461796789234, 32'sd-0.057810735359315316, 32'sd0.06876961468812195, 32'sd0.005121240376727465, 32'sd-0.027459104320562425, 32'sd-0.05160087230601, 32'sd0.038207878984944245, 32'sd-0.073412477774106, 32'sd-0.1345278586052511, 32'sd-0.1759956703036181, 32'sd-0.05687716358874183, 32'sd0.07820923794773192, 32'sd-0.024299766767278085, 32'sd-0.031030364237149062, 32'sd-0.10852567891245882, 32'sd0.04036636268884159, 32'sd0.08570283850391622, 32'sd0.008622663288394273, 32'sd0.07097837041923886, 32'sd0.10113098271489311, 32'sd-0.008769900747239047, 32'sd-0.035641183840146265, 32'sd0.16316895022377056, 32'sd0.0618114931682269, 32'sd-0.1263429905720531, 32'sd-0.12809633744905147, 32'sd-0.11244640103778356, 32'sd0.0024548070359056424, 32'sd-0.04831391565822934, 32'sd0.047376093835308254, 32'sd0.023232368150637287, 32'sd-0.019750213611601453, 32'sd-0.05924398288401103, 32'sd0.01425229359911471, 32'sd-0.004147761157378456, 32'sd-0.0877656364551878, 32'sd-0.06936656150209371, 32'sd-0.19456556411490725, 32'sd0.08390892197605321, 32'sd0.08567575362615734, 32'sd-0.13599977027511767, 32'sd-0.04340515543500736, 32'sd-0.04582976189207888, 32'sd0.12032186150327069, 32'sd0.07429290594468141, 32'sd0.03333764177711924, 32'sd-0.07600265282041696, 32'sd-0.014637554405716569, 32'sd0.04533559143732177, 32'sd0.018954914798582367, 32'sd0.04629378399120684, 32'sd-0.07279831643815556, 32'sd-0.10468616105051474, 32'sd-0.09540686207106205, 32'sd-0.13541218632960758, 32'sd0.011867418140612419, 32'sd-0.07286525494534755, 32'sd-0.02847020098763591, 32'sd-0.03693045658307003, 32'sd0.011502622370319264, 32'sd0.033301483889349816, 32'sd-0.003698481112576945, 32'sd-0.06083881437349862, 32'sd-0.013404891238716226, 32'sd-0.05153282338659402, 32'sd-0.22228378684099873, 32'sd0.008319932896730784, 32'sd-0.032103455488601315, 32'sd-0.11907812477587336, 32'sd-0.03269714996572106, 32'sd0.06120098732812529, 32'sd0.07827978524571365, 32'sd0.005100156444480912, 32'sd0.04468206448897835, 32'sd-0.07929316700190724, 32'sd0.09661648007689513, 32'sd0.09980373427384794, 32'sd-0.0704467649343089, 32'sd-0.0979905169599086, 32'sd-0.07099542566982836, 32'sd-0.1888863207062558, 32'sd-0.1845398530693163, 32'sd-0.09424348722020484, 32'sd0.04746447289557822, 32'sd-0.05280230511772882, 32'sd-0.012074194917492401, 32'sd0.03237052000762245, 32'sd-5.541658998858824e-122, 32'sd-0.013333321335899423, 32'sd-0.008579960849136379, 32'sd-0.027132857792966845, 32'sd-0.07703021642667295, 32'sd-0.11740396765296196, 32'sd-0.10828107380697871, 32'sd-0.09370787022473934, 32'sd-0.15932615876712178, 32'sd-0.16503474214915784, 32'sd0.02545549452161826, 32'sd0.10808862577765388, 32'sd0.06949855355865271, 32'sd0.017560610287626052, 32'sd-0.1058905698152694, 32'sd0.020753998172364327, 32'sd0.04763063176810449, 32'sd0.016908477671338164, 32'sd-0.004975387638855183, 32'sd-0.10016486477290233, 32'sd-0.02384060144092344, 32'sd-0.040745747237959304, 32'sd-0.035587585638672974, 32'sd-0.034937173778, 32'sd0.03920808563130634, 32'sd-0.08767328270173338, 32'sd0.05482352991185266, 32'sd0.023068943966878176, 32'sd-0.0233247931099274, 32'sd0.019471854508902906, 32'sd-0.09023695587620512, 32'sd-0.07745502277951495, 32'sd-0.07147221218078234, 32'sd-0.22655777123450213, 32'sd-0.17394501519734965, 32'sd-0.13453361745665834, 32'sd-0.045836301934481766, 32'sd0.016513305076174427, 32'sd0.17203100945779087, 32'sd0.09430410206955239, 32'sd0.03701178930632897, 32'sd0.0643829516293901, 32'sd-0.032743209381754915, 32'sd0.061654051297413415, 32'sd-0.037645243551481085, 32'sd-0.04902295067216435, 32'sd-0.09616392912419786, 32'sd-0.037357815797266304, 32'sd0.0065765983783515015, 32'sd-0.09135682008037999, 32'sd-0.11647944065934561, 32'sd-0.06633844557226211, 32'sd0.03245093662297748, 32'sd-0.09793751483680775, 32'sd-0.02924600639017424, 32'sd0.06865364022791647, 32'sd-0.011049124811317569, 32'sd0.059780290161855626, 32'sd0.024359831942508656, 32'sd-0.01292062573835082, 32'sd-0.09490985845473213, 32'sd-0.15497979126693762, 32'sd-0.1884643978277601, 32'sd-0.17748453684503723, 32'sd-0.018422768047809974, 32'sd0.06360596010742009, 32'sd0.08167426848363997, 32'sd0.021296872095389493, 32'sd0.11621760144442556, 32'sd0.010886828022662947, 32'sd-0.04104575250154487, 32'sd0.07287759109610725, 32'sd-0.004767514835717295, 32'sd-0.03523962375233823, 32'sd-0.1322695454489399, 32'sd-0.02578659585146464, 32'sd-0.09099498470668195, 32'sd-0.09409245966522067, 32'sd-0.032611127052983926, 32'sd-0.04222346583426636, 32'sd-0.021477670177080452, 32'sd0.007760334029800435, 32'sd0.037644659605470296, 32'sd-0.04541818292525556, 32'sd-4.704539803318957e-123, 32'sd-0.025744131390969267, 32'sd-0.12898900434751087, 32'sd-0.0029527084813202754, 32'sd-0.1545375511384996, 32'sd-0.08251735997521205, 32'sd-0.14078953690100962, 32'sd-0.055553783390074385, 32'sd-0.13903436317956128, 32'sd0.12011117517112206, 32'sd0.18127033221206962, 32'sd0.02452260373910957, 32'sd-0.11669094627028563, 32'sd-0.13645316049598594, 32'sd-0.022708115781518188, 32'sd-0.041688370877566217, 32'sd0.020475149448395073, 32'sd-0.05100379388812989, 32'sd-0.03770285628620837, 32'sd0.012444334394386065, 32'sd0.025540135340216902, 32'sd0.044850417120834846, 32'sd-0.14287664530721894, 32'sd-0.0029521209755818878, 32'sd0.0024715931932872653, 32'sd-0.08122670956690993, 32'sd-0.02698254564781458, 32'sd0.03263005195199183, 32'sd-0.008977097417361784, 32'sd-0.011366017759930755, 32'sd-0.09806068250447662, 32'sd-0.004325733654399395, 32'sd-0.08200603004182794, 32'sd0.01802370595046869, 32'sd-0.13594750858714372, 32'sd-0.08426409213092599, 32'sd-0.014582583031085694, 32'sd0.04140985414252167, 32'sd0.09864165311362856, 32'sd-0.10818261444780272, 32'sd-0.011713838134337334, 32'sd0.06541291265255239, 32'sd0.07648256149465396, 32'sd0.0019066078505907459, 32'sd-0.00819130849682884, 32'sd0.061071106435756556, 32'sd-0.05950465683854232, 32'sd0.0611122161513572, 32'sd-0.11542104000299251, 32'sd-0.13720848279948003, 32'sd-0.07696053319602274, 32'sd-0.04772736031735073, 32'sd0.103703474359256, 32'sd0.09078056266074006, 32'sd0.0882899429908954, 32'sd0.03886046400659127, 32'sd-0.0004959765559509503, 32'sd-0.05192877150483532, 32'sd0.04635000951421572, 32'sd-0.04572580452150517, 32'sd-0.006715609960335114, 32'sd-0.09695087880066022, 32'sd-0.11866204188748708, 32'sd-0.15034244007619132, 32'sd-0.06531058599461992, 32'sd-0.08210095459641052, 32'sd-0.006336517275612485, 32'sd-0.030585980847495427, 32'sd0.027451961433078896, 32'sd0.030281416963103148, 32'sd0.14832518059526936, 32'sd-0.05272480295082466, 32'sd0.051040777768993094, 32'sd0.06294464978815842, 32'sd-0.04811100960965999, 32'sd0.03227273144958218, 32'sd-0.13535249955719506, 32'sd-0.18005408073031243, 32'sd-0.0871960625290965, 32'sd-0.07223608989072977, 32'sd0.028926049038067017, 32'sd0.0554580759047453, 32'sd0.11109026540359503, 32'sd0.02115012183026562, 32'sd-3.980787647144935e-125, 32'sd-0.018506435896592125, 32'sd-0.02039318356151193, 32'sd0.03677195739491104, 32'sd-0.05002817824572904, 32'sd-0.06085182988473241, 32'sd-0.07743623400784841, 32'sd-0.12501362363952617, 32'sd-0.03918159606310272, 32'sd0.04289944828998437, 32'sd-0.09510163222755329, 32'sd-0.03813049956232122, 32'sd0.08659954716003748, 32'sd0.09795276083220862, 32'sd0.07099770106914499, 32'sd-0.13274609015795008, 32'sd-0.01655656030650911, 32'sd0.0031045211977144597, 32'sd0.04375958098365635, 32'sd0.033453596421243854, 32'sd-0.01885226061127927, 32'sd-0.002489240849219716, 32'sd-0.008532484052545607, 32'sd-0.16905045127320076, 32'sd-0.06458459536335498, 32'sd-0.06696457495100522, 32'sd-0.07089133206922292, 32'sd-1.050517525533108e-114, 32'sd-1.0073170175776623e-122, 32'sd-7.202389122531899e-120, 32'sd0.0035506228832035617, 32'sd0.01160723046259102, 32'sd0.03156365588494595, 32'sd0.016205799476308416, 32'sd-0.04460705548264866, 32'sd-0.06986378015616844, 32'sd-0.08733254454669495, 32'sd-0.06827349548029425, 32'sd0.002333841120483705, 32'sd-0.055068794242409326, 32'sd-0.07193259277868197, 32'sd-0.09097547336942834, 32'sd-0.06706491097673323, 32'sd-0.11572513948011924, 32'sd0.05455288566988301, 32'sd-0.05677939739862827, 32'sd-0.0027040335962306558, 32'sd-0.05974676479631385, 32'sd-0.049120526104060376, 32'sd-0.04357286747049573, 32'sd0.044311944424871685, 32'sd-0.047432570182842686, 32'sd-0.01798381141001665, 32'sd0.019018842095491834, 32'sd-0.013921100576244457, 32'sd1.0920152307793366e-119, 32'sd2.070010422938204e-120, 32'sd3.0148623616500537e-121, 32'sd-0.029008193951109876, 32'sd-0.0009081648947853276, 32'sd-0.14234945937628, 32'sd0.034490961792796766, 32'sd0.10021711534259185, 32'sd0.07884070777235419, 32'sd0.02824944734640752, 32'sd0.02728427614869622, 32'sd-0.10056396139753063, 32'sd-0.06284315639802196, 32'sd-0.011802301139160802, 32'sd0.06898872135856435, 32'sd0.14137537151084728, 32'sd0.019473985372673794, 32'sd0.11619687388847362, 32'sd0.06731185382983941, 32'sd0.05016157302876528, 32'sd0.03417009355819826, 32'sd0.06372654584696943, 32'sd-0.007975749754454668, 32'sd-0.004906914106448114, 32'sd-0.01671242138384563, 32'sd-0.030935189809540346, 32'sd0.03388909281202435, 32'sd-0.014106730997955074, 32'sd3.510822594355708e-116, 32'sd5.022833473909399e-119, 32'sd-2.5223712068545935e-126, 32'sd-1.808333835329254e-123, 32'sd0.004016542573946687, 32'sd-0.08582685180919172, 32'sd0.023895266182034084, 32'sd-0.005511761910490817, 32'sd0.09705334229951065, 32'sd0.027614813337045983, 32'sd0.043492542490860625, 32'sd-0.0355066930703924, 32'sd-0.020025595921640243, 32'sd0.036606846190068196, 32'sd-0.062093370783583623, 32'sd-0.02187910891896531, 32'sd0.03321782955942005, 32'sd0.018519160105406062, 32'sd0.11386583987831472, 32'sd0.13756557466208358, 32'sd-0.005402942523059922, 32'sd0.019953463779258558, 32'sd0.005240206840198828, 32'sd0.002480662124212073, 32'sd-0.07498778142615226, 32'sd0.05388184302631361, 32'sd0.0036344349660154948, 32'sd2.958680402721841e-123, 32'sd-3.7997133107594994e-122, 32'sd-3.4633637940279163e-116, 32'sd2.2209125995401356e-129, 32'sd-5.630990390238486e-124, 32'sd1.2559458484777917e-117, 32'sd-0.00811874398663734, 32'sd-0.028625812914567887, 32'sd-0.029917275188820456, 32'sd0.05559956409117904, 32'sd0.12190291187562581, 32'sd0.058527845732770534, 32'sd0.08929660894105275, 32'sd-0.020527688244365343, 32'sd0.07894075192140419, 32'sd0.03669198975252563, 32'sd0.08813525510675094, 32'sd0.0713320069896689, 32'sd0.077495469537608, 32'sd0.08046001855006693, 32'sd-0.04705387607661276, 32'sd-0.07884796983227789, 32'sd0.024403699336231092, 32'sd-0.011047641221224662, 32'sd-0.014653087077744023, 32'sd0.04712374916089242, 32'sd-3.0846506254022987e-120, 32'sd6.2635756281030235e-121, 32'sd-1.60087317410271e-118, 32'sd2.1104980980613028e-119},
        '{32'sd5.339711057777611e-118, 32'sd1.5857372979527998e-125, 32'sd-2.6391418638967014e-124, 32'sd-7.200851426485423e-121, 32'sd-2.7867899948759697e-123, 32'sd-3.935289916766793e-128, 32'sd-3.639994021342185e-115, 32'sd4.0573668926397466e-119, 32'sd1.672086557550253e-123, 32'sd-3.0346711058468058e-121, 32'sd7.5005837921469196e-118, 32'sd-3.103550563391294e-115, 32'sd0.023687165502535256, 32'sd0.07572449858645164, 32'sd-0.006969077554002364, 32'sd0.08108541837571341, 32'sd-7.482215964329381e-125, 32'sd1.4606216725741035e-116, 32'sd-7.80514353068421e-124, 32'sd3.175242978148507e-117, 32'sd-1.1098290783918146e-119, 32'sd4.630957107546843e-115, 32'sd-1.6039677112360113e-117, 32'sd-5.273485930584587e-117, 32'sd-1.3527154708856737e-116, 32'sd-4.7997222124122004e-123, 32'sd1.1366431556699404e-119, 32'sd-7.998212974873708e-125, 32'sd-1.3079071953087704e-123, 32'sd7.564457791516022e-115, 32'sd-2.00808807206865e-118, 32'sd-2.3430713089285502e-122, 32'sd0.0018977148523223778, 32'sd-0.029696991536113816, 32'sd0.0026034469030469074, 32'sd0.0682803759710657, 32'sd-0.003961981989699244, 32'sd-0.014388772000559266, 32'sd0.08827376747327655, 32'sd0.04079722866618252, 32'sd0.011214757589358365, 32'sd-0.04918992216313782, 32'sd-0.08381266062107018, 32'sd-0.03132366108816414, 32'sd-0.1263813078957052, 32'sd-0.0018502982371975934, 32'sd-0.10710719232568382, 32'sd0.07108110505161591, 32'sd-0.020993628160293924, 32'sd0.0023092200797114396, 32'sd-0.011961051547147451, 32'sd-0.020162485307377458, 32'sd-1.859025231262598e-123, 32'sd-5.11636890206181e-124, 32'sd-8.98477539268092e-124, 32'sd5.8425976935031624e-126, 32'sd-7.559769230174402e-124, 32'sd-3.401142917198249e-122, 32'sd0.0427835582798757, 32'sd-0.03104933473945966, 32'sd0.005906609433565447, 32'sd0.0585365972112175, 32'sd0.06936100854027101, 32'sd0.04314071346929779, 32'sd0.01800528674520794, 32'sd0.0752415727557643, 32'sd0.009269558369106234, 32'sd0.052933302275926415, 32'sd0.0969097880143829, 32'sd0.10004715029521422, 32'sd-0.024053985955758538, 32'sd0.05335079989460842, 32'sd0.05546150380541798, 32'sd0.04526130574545812, 32'sd-0.018286867838750644, 32'sd0.008062842739286393, 32'sd0.006019860368154024, 32'sd0.003984734305646077, 32'sd0.0776861899055089, 32'sd0.06027673024198203, 32'sd0.03482552844331357, 32'sd-0.023201331038045482, 32'sd-1.0546505985751095e-121, 32'sd-6.524779459550834e-117, 32'sd-9.953562713434635e-126, 32'sd6.563538695789389e-124, 32'sd-0.0540432883551178, 32'sd-0.03142877579752049, 32'sd0.053982399890818496, 32'sd0.010123671241157402, 32'sd-0.07720952686173053, 32'sd0.061940804123862006, 32'sd-0.010784585259140805, 32'sd0.06855863065321151, 32'sd0.006346168157367641, 32'sd0.22301626433055283, 32'sd0.1731893909724685, 32'sd0.09597328193281443, 32'sd0.032060177441210314, 32'sd0.10566148404946359, 32'sd0.12170989720126152, 32'sd0.04900015793419266, 32'sd0.08618933328025581, 32'sd-0.0026785003514788216, 32'sd-0.10345193560592415, 32'sd0.05730162896877577, 32'sd-0.004334016651347323, 32'sd-0.06206640970140028, 32'sd0.0342636784250179, 32'sd-0.01947838982462081, 32'sd-0.03016106890901362, 32'sd1.4182398931509063e-118, 32'sd3.271244708668074e-116, 32'sd-0.004319502408883464, 32'sd0.028368791187698784, 32'sd-0.12199459696240561, 32'sd0.011240220794025214, 32'sd0.15002519223085778, 32'sd-0.06489483922176355, 32'sd0.014999999362360048, 32'sd0.008342220229379709, 32'sd0.03304301718257519, 32'sd0.1348760217643398, 32'sd0.13787971911333155, 32'sd-0.017689495589277304, 32'sd0.12347000892261188, 32'sd0.0570199339551693, 32'sd-0.013628664819064615, 32'sd-0.01143604573832394, 32'sd-0.03840731988447062, 32'sd-0.06471997399620746, 32'sd0.0806420637391622, 32'sd0.03844225949809589, 32'sd-0.04610545828226635, 32'sd-0.004332746154747987, 32'sd0.04420050775823739, 32'sd0.04893472748277101, 32'sd-0.019698513194624376, 32'sd-0.09466231070558269, 32'sd-0.04432408887639467, 32'sd9.50076368318694e-125, 32'sd0.0019284258811272212, 32'sd-0.06705945173760652, 32'sd0.011125388944507316, 32'sd-0.04199137591373227, 32'sd0.14689557252125932, 32'sd0.03825645610815151, 32'sd0.10019276893263802, 32'sd-0.058658909538389925, 32'sd0.09170541236348358, 32'sd0.09374707784471548, 32'sd-0.05709017886839968, 32'sd-0.2014508186185827, 32'sd-0.1318638261122439, 32'sd-0.10323251114888733, 32'sd0.02195338562862326, 32'sd-0.04428916432370121, 32'sd-0.13656784980676628, 32'sd0.003997139384959973, 32'sd-0.0044432459709633524, 32'sd0.0969091955336074, 32'sd0.04014303433336099, 32'sd0.05855317152367401, 32'sd0.04848700043328233, 32'sd-0.02325641480764066, 32'sd0.012209365646976344, 32'sd-0.127407571942325, 32'sd-0.003176612003215761, 32'sd-3.715675276563002e-122, 32'sd-0.04231044501540596, 32'sd0.03517880339772157, 32'sd-0.040265697983987936, 32'sd-0.014887465822651678, 32'sd0.0039025140855200756, 32'sd-0.04475375790237698, 32'sd-0.08152684883173854, 32'sd0.08466496794039956, 32'sd-0.02616056401829457, 32'sd0.0292370004759688, 32'sd-0.06924401410892403, 32'sd-0.23084043104917562, 32'sd-0.20956636244524468, 32'sd-0.036562077346550585, 32'sd-0.0762698810251955, 32'sd0.006324688796959768, 32'sd-0.09570780442794471, 32'sd-0.13630099922739178, 32'sd-0.01482604581199407, 32'sd0.024991297531664857, 32'sd-0.014286484865097978, 32'sd0.0009606240384486223, 32'sd-0.09725114702836594, 32'sd0.11272453195705859, 32'sd0.12304264182072305, 32'sd-0.05059837154916129, 32'sd0.047390969838421775, 32'sd0.02474190413155082, 32'sd-0.00799795969497519, 32'sd-0.043265218364957087, 32'sd0.04454975386426808, 32'sd-0.05866456885999797, 32'sd-0.11471531189671759, 32'sd-0.12749742556407942, 32'sd0.04965541001736562, 32'sd0.0432176645316911, 32'sd0.1427810260923124, 32'sd-0.025330426373005702, 32'sd-0.04629990461150956, 32'sd-0.17276475899652532, 32'sd-0.1864288332919055, 32'sd-0.17648149271430827, 32'sd-0.14271745732991362, 32'sd-0.08312871006592763, 32'sd-0.08664874951498916, 32'sd-0.028890514333291574, 32'sd-0.11094757962502091, 32'sd-0.010188104539918, 32'sd-0.04794245802636918, 32'sd0.0047038397407139585, 32'sd-0.08652242063470986, 32'sd-0.0012545947525959978, 32'sd-0.07804343611500292, 32'sd0.09807814524973923, 32'sd-0.09331459389494895, 32'sd0.005617483650312982, 32'sd-0.033172974568163614, 32'sd0.03827687792568008, 32'sd0.07589368957915278, 32'sd-0.10948631193378955, 32'sd-0.1545415102227933, 32'sd-0.08028769087473737, 32'sd-0.05646532725286661, 32'sd0.13794110918609712, 32'sd0.06240538037463205, 32'sd0.04331789380654199, 32'sd0.004413864684237786, 32'sd-0.11425324227732755, 32'sd-0.1347638082308559, 32'sd-0.09718386853618799, 32'sd0.02399360392385993, 32'sd-0.01719643650352322, 32'sd0.03758821715800072, 32'sd-0.08272857917495428, 32'sd-0.049449378308918164, 32'sd0.0523329542424027, 32'sd-0.07009227846011118, 32'sd-0.04505858195234356, 32'sd0.049090571403493, 32'sd-0.07360079479544153, 32'sd-0.022429449048778423, 32'sd0.09588319879685234, 32'sd-0.009880335229229521, 32'sd-0.001242314408301146, 32'sd-0.0351154290168725, 32'sd0.03969482733194129, 32'sd0.054757473698985176, 32'sd0.05459465293720852, 32'sd0.09551395917273423, 32'sd-0.12500989025700696, 32'sd-0.05065088445283874, 32'sd-0.10120090514893224, 32'sd-0.026814662432293322, 32'sd-0.018594220475087478, 32'sd-0.06744906506101506, 32'sd0.007027054154802754, 32'sd-0.06573820574754323, 32'sd-0.10142424515975147, 32'sd0.007429727877210749, 32'sd0.13801123841291638, 32'sd0.07362949813124355, 32'sd0.05616441733038019, 32'sd-0.032679250623775684, 32'sd0.059049319903715244, 32'sd-0.06735496212767413, 32'sd-0.031107270478930336, 32'sd-0.18481027899084718, 32'sd-0.10386648824173218, 32'sd0.022549323408375295, 32'sd0.043209250542724516, 32'sd0.030989697445831108, 32'sd-0.007046518758803798, 32'sd-0.0664553257081466, 32'sd-0.022483259902801294, 32'sd0.05411069994324926, 32'sd0.11184367519286775, 32'sd0.11133161601535811, 32'sd-0.05292061388614098, 32'sd-0.12113616022353742, 32'sd-0.10338607734008212, 32'sd-0.049477831221330336, 32'sd-0.02406753893400926, 32'sd-0.02065839693284734, 32'sd-0.19340199209545905, 32'sd-0.1476555892359128, 32'sd-0.09552167002767337, 32'sd-0.027073428374036618, 32'sd0.07583945238577205, 32'sd0.07630458605624452, 32'sd0.001669131167794029, 32'sd-0.017775687107090318, 32'sd0.018299899747617816, 32'sd0.08606071938248289, 32'sd-0.11818384401626708, 32'sd0.028125708302642473, 32'sd0.1038628239243745, 32'sd-0.020985318828388996, 32'sd0.013889251217522627, 32'sd-0.08124782517202161, 32'sd0.056015945035126385, 32'sd0.048909909796337726, 32'sd-0.03445263815911733, 32'sd0.03480536770100598, 32'sd0.11189902880873456, 32'sd0.11448496110939729, 32'sd-0.04428656325487814, 32'sd-0.04143887868847172, 32'sd-0.12226680669231517, 32'sd-0.016297443086299757, 32'sd-0.13470545470554082, 32'sd-0.12127570146898806, 32'sd-0.014475523710512311, 32'sd-0.2214191692719369, 32'sd-0.24621801375085856, 32'sd-0.07122339348660964, 32'sd-0.12268932830391113, 32'sd-0.07531799225651456, 32'sd-0.18021434412456358, 32'sd-0.07670172678974822, 32'sd-0.08698202847839291, 32'sd0.05617555289656177, 32'sd-0.062117300952603344, 32'sd0.026904416817052777, 32'sd-0.06416813457796118, 32'sd-0.04607584255227171, 32'sd0.019839213934197908, 32'sd-0.07125791299464015, 32'sd-0.02912280620080518, 32'sd-0.04898110303844971, 32'sd0.039562481241443036, 32'sd-0.05770426071008529, 32'sd-0.04820671706691642, 32'sd-0.005175939965850542, 32'sd-0.03170281680232166, 32'sd-0.0220402809652149, 32'sd-0.09247007941284442, 32'sd-0.1316877714502413, 32'sd-0.01652666586243425, 32'sd0.055088140803169344, 32'sd-0.024599218936881544, 32'sd-0.024734593518848543, 32'sd-0.041653737169490744, 32'sd-0.11186777019622915, 32'sd-0.04051703244389159, 32'sd-0.14606986385144713, 32'sd-0.13977634166974304, 32'sd-0.2594668554390556, 32'sd-0.12043973768073127, 32'sd-0.010700408996584723, 32'sd0.11294321479931925, 32'sd-0.09877141300821178, 32'sd0.02615741365253767, 32'sd-0.015807662278496976, 32'sd0.04581952621950069, 32'sd-0.07088266397318131, 32'sd-0.010643287012658981, 32'sd0.030321710895810535, 32'sd-0.061350852800144864, 32'sd-0.04998950393981407, 32'sd-0.04970826181867735, 32'sd-0.05596204037289472, 32'sd-0.04727156633142348, 32'sd-0.06101273587980386, 32'sd-0.12351619889702195, 32'sd-0.01130264021222038, 32'sd0.10611408140708771, 32'sd0.11611991161124136, 32'sd-0.02764669310549026, 32'sd0.09878303675646263, 32'sd0.0197060799591179, 32'sd-0.12486910849294058, 32'sd-0.030980182366731914, 32'sd-0.10040089176714749, 32'sd-0.10434889252553022, 32'sd-0.13930100981203225, 32'sd-0.021765571425795605, 32'sd-0.027672589796279838, 32'sd-0.07181787238006312, 32'sd-0.02029398358815629, 32'sd0.03893182315187008, 32'sd-0.03846123699374203, 32'sd0.010118589626005581, 32'sd-0.04756861287158732, 32'sd0.00758769032111285, 32'sd0.006005656233817846, 32'sd0.003291978417193353, 32'sd-0.03416744804969568, 32'sd-0.11018119097744608, 32'sd0.015511298455502205, 32'sd0.08105877405461763, 32'sd-0.1133338984127098, 32'sd-0.16168973557408933, 32'sd0.0006259339603731885, 32'sd0.12597455830786597, 32'sd0.10385476699279243, 32'sd0.1451388211898213, 32'sd0.09796755220376452, 32'sd0.056189269862246524, 32'sd-0.04971264348595675, 32'sd-0.019350918152770194, 32'sd-0.1526959229098626, 32'sd-0.038762622761997836, 32'sd-0.10124953462748267, 32'sd-0.14805299226484633, 32'sd0.013633582194842255, 32'sd-0.011709956372401804, 32'sd0.04870400159709345, 32'sd0.18542698025591253, 32'sd0.07302209539945304, 32'sd0.038160765776137084, 32'sd0.018248116548728516, 32'sd0.07673089036934062, 32'sd0.03690904537116564, 32'sd-0.07149761106307506, 32'sd-0.024474085254839986, 32'sd0.029292600264789772, 32'sd0.15842000848599472, 32'sd0.020040344533721905, 32'sd0.021544380240791434, 32'sd0.019030295938593948, 32'sd0.08571295670523602, 32'sd0.044038215165042686, 32'sd0.13291604566701548, 32'sd0.2192807215442879, 32'sd0.18902650810431185, 32'sd0.09851062467030375, 32'sd-0.08330950078002536, 32'sd-0.06300642304218566, 32'sd0.05580781953419489, 32'sd0.059482756541276285, 32'sd-0.028549232718639524, 32'sd-0.11964446760512784, 32'sd-0.054894128037153496, 32'sd0.06506284191807107, 32'sd0.031993103680298764, 32'sd0.1441465212856664, 32'sd0.010954468496801808, 32'sd-0.05088155230824928, 32'sd-0.04822977858424395, 32'sd-0.027353872982782804, 32'sd-0.025524229051349635, 32'sd-0.08396070001044753, 32'sd0.08384745670856361, 32'sd0.04247706931359966, 32'sd0.07539862801536462, 32'sd0.0849436715287504, 32'sd0.0021474269910685562, 32'sd-0.07200934625799595, 32'sd0.13205358367616138, 32'sd0.10351416566506699, 32'sd0.10184620706744585, 32'sd0.24989721629532066, 32'sd0.16587683342145063, 32'sd0.09791716599993396, 32'sd0.04680954719920349, 32'sd0.09125092530075939, 32'sd0.09699424115488393, 32'sd0.06840894507576632, 32'sd0.009911414021296682, 32'sd-0.10258274349930656, 32'sd-0.0018115478243733245, 32'sd0.0828872142306306, 32'sd0.16268217906343346, 32'sd0.13182087440943474, 32'sd-0.06854248496962853, 32'sd-0.05221878098398027, 32'sd-0.055359929657916425, 32'sd1.5280487181426321e-124, 32'sd-0.04662618598748678, 32'sd-0.057570677920734746, 32'sd0.03824128573371484, 32'sd-0.011889710931754893, 32'sd-0.004214062484219329, 32'sd0.08618410292035783, 32'sd0.05894887604507503, 32'sd0.0611141874408034, 32'sd0.0619937589390373, 32'sd0.026821895370636107, 32'sd0.13626872965528275, 32'sd0.06498346335987419, 32'sd0.01350943643262288, 32'sd0.00957821469834236, 32'sd-0.06497031056936853, 32'sd0.10096083045217827, 32'sd-0.003443904429796283, 32'sd0.06768639489407369, 32'sd0.005721320057730188, 32'sd0.0194729527526091, 32'sd0.017546707001278437, 32'sd0.09726831655711572, 32'sd0.034739288779862335, 32'sd-0.050069983485398845, 32'sd-0.024602836642574885, 32'sd-0.12823205427410597, 32'sd0.029697723475242552, 32'sd-0.0016438002408305501, 32'sd0.004346308375506011, 32'sd0.095982159007083, 32'sd-0.04482830442626985, 32'sd-0.051602998072023634, 32'sd0.07590927566374825, 32'sd0.08659302586817187, 32'sd0.021192499145903067, 32'sd0.08711291128732451, 32'sd0.022436072116479668, 32'sd0.09487381214211944, 32'sd0.10024312253424825, 32'sd0.08528809926820957, 32'sd0.07832419828623811, 32'sd0.05907225052064392, 32'sd0.1061570038136063, 32'sd-0.020810391293806907, 32'sd0.13476862489939812, 32'sd0.12340658739573299, 32'sd0.03976766229167858, 32'sd-0.03234346429555681, 32'sd0.006097041008507118, 32'sd-0.041654809740652755, 32'sd-0.1021963160010634, 32'sd-0.045625690118157376, 32'sd0.09885889190589137, 32'sd-0.09077678029405432, 32'sd-0.014127022735688905, 32'sd0.03392377640215083, 32'sd-0.0066448056919039935, 32'sd0.015627149811182676, 32'sd-0.15852495073846923, 32'sd0.024282971230269665, 32'sd-0.04497908137349934, 32'sd-0.01957587118600158, 32'sd-0.07023246836405733, 32'sd-0.039981188008249596, 32'sd0.0021509058016483808, 32'sd0.15902523810648145, 32'sd0.05869405223829628, 32'sd0.08639512117886489, 32'sd0.06697912171740239, 32'sd0.08818320135633802, 32'sd0.069212397143605, 32'sd0.016321884415901225, 32'sd0.08034748346417697, 32'sd0.1892699527382712, 32'sd0.00828929459778996, 32'sd0.08946623906316756, 32'sd0.15406617037271939, 32'sd0.054894661022786395, 32'sd0.05639635675318851, 32'sd-0.23699919678562165, 32'sd0.026582867372100055, 32'sd-0.0015676184697289912, 32'sd-0.062996396195567, 32'sd-3.7376055657890486e-116, 32'sd-0.07509816885996204, 32'sd-0.01616249875449674, 32'sd-0.16948256166753545, 32'sd0.1448939056728887, 32'sd-0.10221334807776773, 32'sd-0.03604225404339849, 32'sd0.016235824116312716, 32'sd0.08369434429545296, 32'sd0.20352747975120664, 32'sd0.16865575050426931, 32'sd0.12132628658503354, 32'sd0.013783033218090664, 32'sd-0.010355336823392363, 32'sd0.02998848790475986, 32'sd-0.0789612990406552, 32'sd-0.10651079444270564, 32'sd0.037264838745802324, 32'sd0.16135240673358464, 32'sd0.010753386113687135, 32'sd0.06237434608435253, 32'sd0.143609763044366, 32'sd0.06513987287157438, 32'sd0.01773130021979622, 32'sd-0.1332943897015288, 32'sd0.0045608924009578845, 32'sd0.06839948262645162, 32'sd-0.05552809240643663, 32'sd-0.05325660349104722, 32'sd0.08208229218517778, 32'sd0.058816486792377484, 32'sd-0.0443431161999028, 32'sd0.0990761048530884, 32'sd0.04570134224930809, 32'sd-0.020057420107986265, 32'sd0.030341775692063633, 32'sd0.0062952704415490226, 32'sd0.13900997893492423, 32'sd0.09380384474911174, 32'sd0.0035135322926170957, 32'sd0.07815207112192431, 32'sd0.0919148611396223, 32'sd-0.03719015212649714, 32'sd-0.07788843250392319, 32'sd0.016631542303609755, 32'sd-0.030462262659570884, 32'sd0.0825416354944531, 32'sd0.12892844396128544, 32'sd0.13086207485480886, 32'sd0.09872129943157308, 32'sd0.02754545822487003, 32'sd0.0052153714553113085, 32'sd-0.12760829803320628, 32'sd-0.09941628970062127, 32'sd0.07664323148919347, 32'sd-0.019476654669795715, 32'sd-0.004128594581474114, 32'sd-0.055918968263121184, 32'sd-0.07040487422805805, 32'sd0.007911806773442021, 32'sd-0.10072725661876351, 32'sd-0.005582990275344186, 32'sd-0.049550245055169286, 32'sd-0.09032352229939791, 32'sd-0.07172549495266481, 32'sd0.014402172656174972, 32'sd0.015449229882188564, 32'sd-0.08395097205154825, 32'sd-0.04528472116582439, 32'sd-0.030039718192787453, 32'sd-0.04378602284949525, 32'sd-0.02171689248906169, 32'sd0.01864369417889069, 32'sd-0.14232296805641556, 32'sd-0.007677354843305884, 32'sd0.062332972877760864, 32'sd0.06162007822680512, 32'sd-0.03961664276286354, 32'sd-0.035668679637856554, 32'sd-0.06950507328881306, 32'sd0.0027960235973623405, 32'sd-0.01658511889104804, 32'sd-0.015318141711675353, 32'sd-0.008350559806673414, 32'sd-6.586294350899677e-126, 32'sd-0.0033711802205700367, 32'sd0.15691003022776617, 32'sd0.03186562780327329, 32'sd0.004844236345943974, 32'sd-0.049125937747807734, 32'sd-0.00935165924439968, 32'sd-0.07548263325449185, 32'sd-0.08161621616063157, 32'sd-0.01763772635281841, 32'sd-0.027690738889871638, 32'sd-0.13923356764590614, 32'sd-0.007952546567497755, 32'sd-0.10285784825481165, 32'sd-0.03062822546081809, 32'sd-0.04604481936031858, 32'sd-0.18828333072353748, 32'sd-0.1408340313215266, 32'sd0.03784508924097004, 32'sd-0.019408826546838773, 32'sd-0.04869720906717577, 32'sd0.03614657347525536, 32'sd-0.033827031819961675, 32'sd-0.13584960456570663, 32'sd-0.07537860316078827, 32'sd0.03851105992256829, 32'sd0.04145391202301601, 32'sd-8.628711549205293e-125, 32'sd-4.495774720266755e-116, 32'sd8.563877923837628e-129, 32'sd0.033841415366262576, 32'sd-0.12237465654529008, 32'sd0.029820030541016423, 32'sd-0.10229856441806764, 32'sd-0.06967790394810747, 32'sd-0.13313925781893773, 32'sd-0.23001802343905556, 32'sd-0.15824218638387147, 32'sd-0.15913510644218812, 32'sd-0.22325349834053146, 32'sd-0.13235035658594124, 32'sd-0.020877890517312925, 32'sd-0.1409984141576003, 32'sd-0.047050115756090964, 32'sd0.0436636072423389, 32'sd0.016268396095594544, 32'sd-0.05990992367443223, 32'sd-0.10298002469307456, 32'sd-0.11242918951716505, 32'sd-0.004001064599521882, 32'sd-0.056907796898694865, 32'sd0.011073780166258257, 32'sd-0.006248159893756262, 32'sd-0.013390294538939165, 32'sd0.027296195736205356, 32'sd5.898534815728622e-128, 32'sd-4.2264960539764735e-118, 32'sd-3.091466193874744e-119, 32'sd-0.04340701981415327, 32'sd-0.02778095707383992, 32'sd-0.07191121550090815, 32'sd-0.0382617806753321, 32'sd-0.05436009597776779, 32'sd-0.0499284549878508, 32'sd-0.06707453856499836, 32'sd-0.04218283330230872, 32'sd-0.14778771127708246, 32'sd-0.07420365686517705, 32'sd0.0016276762282030324, 32'sd-0.19995566725244598, 32'sd-0.04814275584563002, 32'sd0.033195274983084666, 32'sd0.06694886830976064, 32'sd-0.08868249276600883, 32'sd0.041314759512111554, 32'sd-0.15217187140739571, 32'sd-0.0005265428813886134, 32'sd-0.13078695016273326, 32'sd-0.05425979255727488, 32'sd-0.06643478681490222, 32'sd0.02867024185104131, 32'sd0.03152383016623849, 32'sd0.07442531817985294, 32'sd-1.82568606746161e-121, 32'sd2.1569631715655265e-128, 32'sd-2.245794154884428e-129, 32'sd2.7081519197431783e-122, 32'sd-0.026111642362493227, 32'sd0.01189450315529031, 32'sd0.006107665960492689, 32'sd-0.0009567729740243922, 32'sd-0.06391489480820729, 32'sd-0.062299657579732715, 32'sd0.03459017169318379, 32'sd0.035712466149523905, 32'sd0.026978927104621696, 32'sd-0.06887238523020893, 32'sd0.07334962983380201, 32'sd0.00454240656654558, 32'sd-0.004933024548006611, 32'sd0.0562989703163448, 32'sd-0.03274106205821807, 32'sd-0.11884984029876372, 32'sd-0.043922413795911955, 32'sd-0.05381346698790111, 32'sd-0.04617493695458609, 32'sd0.0019745721416909454, 32'sd-0.08814285861434175, 32'sd0.028043280271290924, 32'sd-0.03474339528707758, 32'sd5.118414291162176e-127, 32'sd-3.09473546951713e-125, 32'sd-5.8744173637735945e-120, 32'sd-1.6629883463751507e-126, 32'sd-3.460522364713417e-123, 32'sd3.56596231280227e-117, 32'sd-0.043626177438427075, 32'sd-0.04618701850601129, 32'sd-0.032500170439689016, 32'sd0.015994039410384332, 32'sd-0.058327263268048754, 32'sd-0.04496971451585103, 32'sd0.0035023184099593208, 32'sd0.0667879005025078, 32'sd0.023389108530660917, 32'sd-0.012765416560297097, 32'sd0.059202047378677805, 32'sd0.0407139953031874, 32'sd-0.028301269294461265, 32'sd-0.05387176042581296, 32'sd-0.04256217892135088, 32'sd-0.021684950708587555, 32'sd0.03423152823237915, 32'sd-0.0931056328921562, 32'sd-0.002409351897933465, 32'sd0.013329994703478157, 32'sd-8.73351281261785e-117, 32'sd-3.145727078243268e-120, 32'sd1.5249958814118951e-125, 32'sd-4.84860544602373e-123},
        '{32'sd-7.501859578027104e-115, 32'sd-7.87141542599156e-124, 32'sd6.770414920059848e-119, 32'sd-3.7189744812885716e-126, 32'sd-5.106949483661508e-117, 32'sd-4.65139753287769e-120, 32'sd-1.8081359821222793e-124, 32'sd-1.978408533004626e-121, 32'sd1.8974773880212057e-126, 32'sd-9.180922923123877e-122, 32'sd-1.2551484885815442e-127, 32'sd-3.0892719691608865e-122, 32'sd-0.011245649145183657, 32'sd0.013081991847505466, 32'sd-0.03890823202854701, 32'sd-0.05022455191695397, 32'sd3.9025582755931823e-123, 32'sd-2.6854192533309494e-123, 32'sd-2.25822265692397e-124, 32'sd3.6647101654423554e-122, 32'sd-5.309193075186135e-118, 32'sd6.832669261842394e-118, 32'sd5.270888529663458e-125, 32'sd1.0008655906842718e-122, 32'sd-1.6296058098394563e-115, 32'sd3.0575433274712164e-114, 32'sd3.575351158724034e-123, 32'sd-1.1013105069737328e-119, 32'sd1.0714135519648082e-121, 32'sd3.5150114342492394e-122, 32'sd6.366399972304188e-115, 32'sd-1.0354775829250456e-124, 32'sd-0.004449085641649436, 32'sd-0.09459253682869344, 32'sd-0.005806340651972763, 32'sd-0.10068076828703511, 32'sd-0.0772088677392096, 32'sd-0.1096487434235764, 32'sd-0.1288575936569958, 32'sd-0.0178015252035871, 32'sd0.03089403324934105, 32'sd-0.05896943411044926, 32'sd-0.03906768855022665, 32'sd0.009099810508914377, 32'sd-0.07471369108776518, 32'sd-0.12134772780779514, 32'sd-0.02594074123014919, 32'sd-0.04520695748010205, 32'sd0.023420716881229483, 32'sd-0.07210232262269244, 32'sd0.00914161518630209, 32'sd-0.016358456270082034, 32'sd7.043476758485086e-118, 32'sd6.582389183628244e-126, 32'sd3.868205873414594e-123, 32'sd1.1355339657167074e-119, 32'sd-3.088235372967573e-118, 32'sd3.0261321684211435e-117, 32'sd-0.04604834193315149, 32'sd-0.01148760751076642, 32'sd-0.08078230307024373, 32'sd-0.09626434588436723, 32'sd-0.053269137863239405, 32'sd-0.06808867499087273, 32'sd-0.045648810167138065, 32'sd-0.09800858106066168, 32'sd-0.06093361317872106, 32'sd-0.14835653058371864, 32'sd-0.12464148075647856, 32'sd-0.1299089603785456, 32'sd-0.11012958248845284, 32'sd-0.11282014021061891, 32'sd-0.034968941087035105, 32'sd-0.08897729280186348, 32'sd0.02812558705633985, 32'sd0.01540742143502955, 32'sd0.01693229241233515, 32'sd-0.06779043240233772, 32'sd0.0360217043067774, 32'sd-0.08407869902110168, 32'sd-0.08407075614363319, 32'sd-0.08195465162395146, 32'sd-2.1529610788469817e-127, 32'sd2.496516796840765e-118, 32'sd2.033955665996611e-127, 32'sd-1.1056761709924232e-122, 32'sd-0.011440413112794421, 32'sd-0.03617875849051429, 32'sd-0.08356436980999161, 32'sd0.033565993020482236, 32'sd-0.007726614555400575, 32'sd-0.09983499495324918, 32'sd-0.03573096633041894, 32'sd-0.14418660076093373, 32'sd-0.04755114047552422, 32'sd-0.16368362851558152, 32'sd-0.09865364330856141, 32'sd-0.2651062128466459, 32'sd-0.10907717013184574, 32'sd-0.020735484115607803, 32'sd0.0312405589612119, 32'sd-0.15787000953658148, 32'sd-0.03334491231048087, 32'sd-0.12194307632340914, 32'sd-0.12556159755089533, 32'sd0.056003760414897394, 32'sd0.07166906112225943, 32'sd0.03220577517539175, 32'sd-0.04391601798477257, 32'sd-0.04467783377585325, 32'sd-0.05526777120805822, 32'sd1.7688631637801839e-121, 32'sd-8.760990380909167e-129, 32'sd0.029509325821853852, 32'sd-0.10570554667248526, 32'sd-0.031085503492706508, 32'sd-0.0795521759498281, 32'sd-0.023777081025630618, 32'sd-0.03592928271379124, 32'sd-0.046275850455768874, 32'sd-0.11882191164338424, 32'sd-0.257582131571407, 32'sd-0.04319308833945085, 32'sd-0.06912671844677115, 32'sd-0.11807723061938147, 32'sd-0.24534107749977987, 32'sd-0.182176431478226, 32'sd0.03818950777692557, 32'sd-0.036488039328124534, 32'sd-0.044073940631647116, 32'sd0.0039463621426999735, 32'sd-0.1635230758657547, 32'sd-0.010356678717550532, 32'sd0.0048933695515543775, 32'sd-0.009888938703483022, 32'sd-0.01706307618075172, 32'sd-0.0667442547369841, 32'sd-0.0664692899376241, 32'sd-0.0010655831043921114, 32'sd-0.022684335022404606, 32'sd-1.8396783790257642e-121, 32'sd-0.009286357939563044, 32'sd-0.12175873302071574, 32'sd-0.15864848018167818, 32'sd-0.08377402083855107, 32'sd0.06403289210548127, 32'sd0.051505980863367204, 32'sd0.008547880805965687, 32'sd0.03558088357770602, 32'sd0.025854557793999124, 32'sd0.02656223152463129, 32'sd0.10021043842489946, 32'sd0.027988205061161908, 32'sd-0.10138193890029404, 32'sd-0.009752360914388162, 32'sd0.062049280176615755, 32'sd-0.04782191560560577, 32'sd-0.008934417747134134, 32'sd0.000592581376320811, 32'sd0.02686597214568141, 32'sd-0.14903508896151652, 32'sd-0.10708435427396341, 32'sd-0.10791858144863177, 32'sd-0.1790092175743308, 32'sd-0.04787199201213387, 32'sd-0.1097401454396883, 32'sd-0.005205121354058454, 32'sd-0.10702978066850449, 32'sd-2.0958164927020113e-127, 32'sd0.011826812608201258, 32'sd0.09389544191588756, 32'sd0.06605350795436757, 32'sd0.08410304794305451, 32'sd0.10980414496512769, 32'sd-0.023380807888730426, 32'sd-0.022082549991381033, 32'sd0.08219490484144748, 32'sd0.16772332280992566, 32'sd0.1208176268003192, 32'sd0.05199011972327136, 32'sd0.023020086765346764, 32'sd-0.04241686883130952, 32'sd-0.1045953340150634, 32'sd0.058606612286541966, 32'sd0.11552892851343881, 32'sd0.1640987696521925, 32'sd0.13320293803675679, 32'sd0.06892126190859008, 32'sd0.0022238748258630297, 32'sd0.05837216607798287, 32'sd-0.020926860673557618, 32'sd-0.18134229816776856, 32'sd-0.1354920674826524, 32'sd-0.07375028607061365, 32'sd-0.13910228543830522, 32'sd-0.1123540396627147, 32'sd-0.04638260198732827, 32'sd0.03972216896781398, 32'sd0.0543075820404834, 32'sd0.024239607587607775, 32'sd0.19439073139004998, 32'sd-0.03776105004203423, 32'sd0.09852970048883851, 32'sd0.1398001512658042, 32'sd0.02425746033579015, 32'sd0.06628095511069267, 32'sd-0.02551724628357074, 32'sd-0.03333727889195055, 32'sd-0.14660955368667644, 32'sd-0.12289325119264037, 32'sd-0.037641263416526696, 32'sd-0.03652773405893026, 32'sd0.023046102220872715, 32'sd-0.035978494100190564, 32'sd0.06602310189892249, 32'sd0.021639148855171778, 32'sd0.046257412573878685, 32'sd0.07448542237336359, 32'sd-0.02432855171437253, 32'sd-0.019004327744558038, 32'sd0.019089200016987017, 32'sd-0.04937578504791485, 32'sd-0.20938222943816012, 32'sd-0.05528685963550189, 32'sd0.00760535943027603, 32'sd0.06922631011054488, 32'sd0.06879709353135431, 32'sd-0.04444071546605361, 32'sd-0.01792576843110172, 32'sd-0.021188404199778504, 32'sd-0.011699564221833577, 32'sd0.08105300364061489, 32'sd0.075883850342042, 32'sd0.054396534966491814, 32'sd0.08688764262358342, 32'sd-0.013053265123769179, 32'sd-0.07067429783817365, 32'sd-0.17375323875461265, 32'sd0.009779153308010734, 32'sd0.042687160685538586, 32'sd0.020107134982248535, 32'sd-0.10094532861786068, 32'sd0.06659564499094156, 32'sd-0.014949858631954294, 32'sd-0.061327026205140626, 32'sd0.0011971540036740454, 32'sd-0.14707737078827665, 32'sd-0.07587995350547601, 32'sd0.05166126876268073, 32'sd-0.03899061510492032, 32'sd-0.09339911559064683, 32'sd-0.10281367301364933, 32'sd-0.005775565097942107, 32'sd-0.04122837172582431, 32'sd-0.01017061761232883, 32'sd-0.03159150593543162, 32'sd0.10734809169394692, 32'sd-0.034892968497597945, 32'sd0.019317456530869633, 32'sd-0.007288655797270277, 32'sd0.06287148735367043, 32'sd0.13916191193784733, 32'sd0.0937930214443614, 32'sd0.0935097447785593, 32'sd0.105855412323804, 32'sd-0.0877124595390822, 32'sd0.12006267166604537, 32'sd-0.03939664568334953, 32'sd-0.14450488535662082, 32'sd-0.03814281434235918, 32'sd-0.05215400836346439, 32'sd-0.02846048054728048, 32'sd-0.056741797877763366, 32'sd-0.06307430398835943, 32'sd-0.13580800928043127, 32'sd-0.1607806759956948, 32'sd0.04611368742358447, 32'sd0.00024099392242105968, 32'sd-0.026128022579098135, 32'sd0.03857943380884972, 32'sd-0.0010432905346498204, 32'sd0.016868574694374167, 32'sd0.05213100078116877, 32'sd-0.04457618973188618, 32'sd0.11500146442811185, 32'sd-0.04031348000600359, 32'sd-0.02015884353403313, 32'sd-0.10372485840332804, 32'sd0.12246973670721428, 32'sd0.2189052497340157, 32'sd0.041249259120630634, 32'sd0.04701572944779736, 32'sd-0.06312960638709537, 32'sd0.061178966772093155, 32'sd0.1143022304431199, 32'sd-0.10944152909130225, 32'sd-0.12365163886129744, 32'sd-0.1366833687073825, 32'sd-0.09300135847180722, 32'sd0.01039225911965487, 32'sd-0.04449771870340981, 32'sd-0.08933777185558453, 32'sd-0.1862706946096562, 32'sd-0.12319614730727853, 32'sd0.006717542141780678, 32'sd0.019344428169691896, 32'sd-0.013820264248560997, 32'sd-0.0676575411056263, 32'sd-0.05161259024960751, 32'sd-0.051978725860470296, 32'sd0.11441952136627356, 32'sd0.0672294692083555, 32'sd-0.040991476528266665, 32'sd-0.17493312069233508, 32'sd-0.10511388252477127, 32'sd-0.031014378362292882, 32'sd0.13025744010639598, 32'sd0.1445339019665557, 32'sd0.028572001495222897, 32'sd0.061071908380787236, 32'sd-0.07932364598277976, 32'sd-0.07014524187716593, 32'sd0.03638848965446044, 32'sd0.058046799700078026, 32'sd-0.10630794124381308, 32'sd-0.0064165765191454395, 32'sd0.026780282783070614, 32'sd0.14098345888038394, 32'sd0.08680240543468164, 32'sd-0.035458411070748375, 32'sd0.020532036862299003, 32'sd-0.021118161765176058, 32'sd0.005317273063804903, 32'sd-0.02688019895468632, 32'sd-0.001100386283907286, 32'sd-0.020495895955859777, 32'sd-0.0633399802748079, 32'sd-0.06847873262148559, 32'sd0.08388800596457102, 32'sd-0.052481372168466864, 32'sd0.11409138321006597, 32'sd-0.0045007234997253886, 32'sd0.08145624448825213, 32'sd0.07677672804011605, 32'sd0.12041858209992876, 32'sd0.028899522762644195, 32'sd0.09623992237111598, 32'sd-0.013561700899178419, 32'sd-0.16601683723997748, 32'sd-0.0780521623465462, 32'sd-0.12084427952555934, 32'sd-0.05837894527940068, 32'sd-0.024919577719634482, 32'sd-0.04077673997145846, 32'sd0.12530751826235997, 32'sd0.12775458528419245, 32'sd-0.033303451007184716, 32'sd0.037350639259828324, 32'sd0.03023777210283482, 32'sd-0.07433326382383496, 32'sd-0.05615862455371501, 32'sd0.03404402551667504, 32'sd-0.021594680181170285, 32'sd0.041459391224896926, 32'sd-0.04890591151431397, 32'sd-0.0356943589403271, 32'sd-0.047143110810849785, 32'sd-0.06722913597923029, 32'sd-0.013063952915489896, 32'sd-0.03960568027028386, 32'sd0.09872442893057395, 32'sd0.07126451268603053, 32'sd0.0782467760923891, 32'sd-0.02913398337597926, 32'sd0.08488923103745541, 32'sd0.0777796335580121, 32'sd-0.08936016283371127, 32'sd0.0739849935967449, 32'sd-0.05359539634749899, 32'sd0.07405296644651765, 32'sd0.015271582831060086, 32'sd0.0013165635879624424, 32'sd0.13291510098506018, 32'sd0.043475189853386935, 32'sd0.04381339455554564, 32'sd0.02603024877754512, 32'sd-0.042346168186955795, 32'sd-0.09210813457204463, 32'sd-0.0857265551988919, 32'sd-0.05814187706510871, 32'sd-0.002806496469024295, 32'sd-0.05046022621240607, 32'sd-0.05418841973997525, 32'sd-0.06314115483258223, 32'sd-0.08056814587937192, 32'sd-0.0627953308252353, 32'sd-0.022813444093628663, 32'sd0.020301001920529884, 32'sd0.052980668224175444, 32'sd0.05333758334528172, 32'sd0.003616709218501499, 32'sd0.06313923032298362, 32'sd0.08866995517057513, 32'sd0.11378684066506871, 32'sd0.031036339855261382, 32'sd0.12053503348492448, 32'sd0.14518015454565653, 32'sd0.12754659574162872, 32'sd0.007458597087416054, 32'sd0.1474244168593776, 32'sd0.23273658183805532, 32'sd0.18575786158646054, 32'sd-0.0034663718902097503, 32'sd-0.03689025767955956, 32'sd-0.17912801438100748, 32'sd-0.17348900228660405, 32'sd-0.10996884332048071, 32'sd0.023048916286731187, 32'sd-0.14124290569770104, 32'sd-0.04106690810085661, 32'sd-0.07496697669235952, 32'sd-0.06333772078852865, 32'sd-0.06184911088639148, 32'sd-0.06252492674920992, 32'sd0.008149579961481251, 32'sd-0.010675490944913317, 32'sd-0.0284126121309941, 32'sd0.11047267327932135, 32'sd-0.03578057033642891, 32'sd0.07433233181409028, 32'sd0.07948448644588241, 32'sd0.01741342187807481, 32'sd0.028846506248162374, 32'sd0.03955493137556708, 32'sd0.11789571369869624, 32'sd0.11447963938266065, 32'sd0.08983019047641902, 32'sd0.23725191133517337, 32'sd0.17960390501809287, 32'sd0.016975718717721668, 32'sd0.003105185425399436, 32'sd-0.030569905202765556, 32'sd-0.0237806667115684, 32'sd-0.12625103046127864, 32'sd-0.10365008035355901, 32'sd-0.10107443339053111, 32'sd-0.06155159957366046, 32'sd0.05002926594240907, 32'sd0.026224739128929024, 32'sd-0.022311624556098635, 32'sd-0.025976808001655673, 32'sd-0.007977522247280239, 32'sd-0.08667623305714882, 32'sd-0.1331159826677382, 32'sd0.04334287958699453, 32'sd0.06919637169569823, 32'sd0.02931163742012188, 32'sd0.03919181214495793, 32'sd0.056956341542875925, 32'sd0.05886227876757966, 32'sd0.049944053804057524, 32'sd0.11390123747195725, 32'sd0.06395997186293334, 32'sd0.10193275256956624, 32'sd0.062238588015201976, 32'sd0.05509341799731934, 32'sd-0.027128115583397585, 32'sd0.007257413185256397, 32'sd-0.028411548398765554, 32'sd0.0021835137142235516, 32'sd-0.009715071047285724, 32'sd-0.16346095700246438, 32'sd-0.1383944199524746, 32'sd-0.12975710643063307, 32'sd-0.15946635675358217, 32'sd-0.052116068583958786, 32'sd-4.7282870366858844e-123, 32'sd-0.11227634002662999, 32'sd0.011986986887051902, 32'sd-0.12909192263547836, 32'sd-0.13473408687552552, 32'sd-0.03564473254993946, 32'sd0.08322779863882405, 32'sd0.105855990110296, 32'sd0.006896696647853839, 32'sd0.10254243393882637, 32'sd-0.006983631688108341, 32'sd0.05660231151371746, 32'sd-0.02169783408048203, 32'sd0.015000925163388294, 32'sd0.06371408999005211, 32'sd0.03518767797305607, 32'sd0.06238353153466717, 32'sd0.056943853250754364, 32'sd0.03386267529766456, 32'sd-0.00016760421790281902, 32'sd-0.12781718332618758, 32'sd-0.056115006554931304, 32'sd0.017127187435476712, 32'sd0.004033378544251672, 32'sd-0.049933328069844726, 32'sd0.05809037478624168, 32'sd-0.1706973781616159, 32'sd-0.05328496326873782, 32'sd-0.07771136235744781, 32'sd-0.009942566901719272, 32'sd0.04380052466484801, 32'sd-0.12677367769107487, 32'sd-0.019414163765332323, 32'sd-0.17369863274635763, 32'sd-0.04644632650552765, 32'sd0.11548700501429218, 32'sd0.11278364641392334, 32'sd0.03339112903650464, 32'sd0.038524131483995444, 32'sd-0.024206231370039993, 32'sd0.026750895601871896, 32'sd0.061119576073932445, 32'sd0.021213111958968005, 32'sd0.11692948901424231, 32'sd-0.053890304378622696, 32'sd0.05219830375887923, 32'sd-0.07395306178150693, 32'sd-0.05218183867394915, 32'sd-0.15336855980912018, 32'sd-0.049740624270923295, 32'sd0.11693540532691656, 32'sd0.08407773132562055, 32'sd-0.11126467103246056, 32'sd-0.03577561772946766, 32'sd-0.009268947641783312, 32'sd-0.11978610035941398, 32'sd-0.0394377141432891, 32'sd-0.0013917736630315422, 32'sd-0.015148069327946554, 32'sd-0.05654842560755849, 32'sd-0.0859264479477369, 32'sd-0.1225631884395704, 32'sd-0.19786060151438134, 32'sd-0.05575062208832911, 32'sd0.04985509490928479, 32'sd-0.004638078640112825, 32'sd0.001531824531508912, 32'sd0.022597357742472266, 32'sd-0.06461337646066304, 32'sd-0.11760748358203031, 32'sd0.14979244801149696, 32'sd0.07757278931074471, 32'sd0.0256292191969691, 32'sd0.029073590171955543, 32'sd-0.060052192307691175, 32'sd-0.09003352167064636, 32'sd-0.15824785551231652, 32'sd-0.1067851741807727, 32'sd-0.015389935790503977, 32'sd-0.04614981412272042, 32'sd0.02549761904797028, 32'sd0.03410220924011184, 32'sd0.0017753568350738107, 32'sd-0.06915390819752501, 32'sd1.1452727232014644e-115, 32'sd-0.0036193977945654467, 32'sd-0.08159458836216808, 32'sd-0.04936526297349568, 32'sd-0.17181327260973672, 32'sd-0.25421897972937235, 32'sd-0.2673149876356845, 32'sd0.007023598148576314, 32'sd-0.12962002016776394, 32'sd-0.06630979538063103, 32'sd0.03194147323115578, 32'sd-0.10843780574478248, 32'sd-0.12706905687567474, 32'sd-0.08050140110121727, 32'sd0.09823300152541864, 32'sd0.026034345955887803, 32'sd0.03928945718363466, 32'sd0.009324230568574895, 32'sd-0.14001902625970197, 32'sd-0.17448655855463865, 32'sd-0.2005726547701972, 32'sd-0.028460867452257135, 32'sd-0.01183791112217382, 32'sd0.03316910644753526, 32'sd-0.012675865489488704, 32'sd0.048669011388258854, 32'sd-0.05966781287969063, 32'sd-0.0030753446310791605, 32'sd-0.013768917759720072, 32'sd-0.11449099148713285, 32'sd-0.04063729711755649, 32'sd-0.021324720488118225, 32'sd-0.025342949649064774, 32'sd-0.15981941411640632, 32'sd-0.09945302438997018, 32'sd-0.13831577005599255, 32'sd-0.11164870483008613, 32'sd-0.03310997995621079, 32'sd0.008120912306589954, 32'sd-0.02386881434322756, 32'sd-0.10752681119035183, 32'sd-0.13302832432278483, 32'sd-0.1434724469195615, 32'sd-0.10242203475336194, 32'sd0.10524752200261074, 32'sd0.03519871112382813, 32'sd-0.149941920715084, 32'sd-0.14123084450896267, 32'sd-0.1832399380457748, 32'sd-0.05795906659232447, 32'sd-0.1567238729684451, 32'sd-0.01661831073299643, 32'sd-0.06126059041250628, 32'sd-0.0008708442673382967, 32'sd0.05468423557468918, 32'sd0.0172181958677316, 32'sd-0.08372634150111066, 32'sd-0.09661345962742501, 32'sd-0.04304067305123124, 32'sd-0.057501000207022465, 32'sd0.0010320562598685739, 32'sd-0.006851374074503352, 32'sd-0.04320297546696786, 32'sd-0.16373306161403695, 32'sd-0.20610237154505198, 32'sd-0.07141346573589319, 32'sd0.03816447025744691, 32'sd-0.09992019491848157, 32'sd0.014549801174472812, 32'sd-0.0975630483620912, 32'sd-0.06850761311139461, 32'sd-0.17739756148802197, 32'sd-0.023403513220634106, 32'sd-0.11776958693182162, 32'sd-0.04887465925483076, 32'sd-0.14131097854825012, 32'sd-0.0929038898490622, 32'sd-0.2453752363142225, 32'sd-0.048510298009598114, 32'sd-0.10664729616104272, 32'sd-0.06429241545997844, 32'sd0.03506756004701615, 32'sd-0.0002381797777925515, 32'sd0.02095378219967855, 32'sd-3.1548150918112604e-116, 32'sd-0.03989780540614907, 32'sd-0.12368980223011704, 32'sd-0.05737257088179148, 32'sd-0.04775588476418063, 32'sd-0.01721797673531769, 32'sd-0.00642610263487012, 32'sd-0.029156184726089544, 32'sd-0.11279108538052016, 32'sd-0.09976933016026485, 32'sd-0.10078604061125514, 32'sd-0.14455994260826976, 32'sd-0.08494908187102367, 32'sd0.05980869011428235, 32'sd0.02802479848865856, 32'sd-0.0959269553437601, 32'sd-0.018144397481625982, 32'sd-0.12047738584862286, 32'sd0.009836900908842209, 32'sd-0.047980591427158374, 32'sd-0.11799029681856113, 32'sd-0.1754712677901055, 32'sd-0.047969889267796904, 32'sd-0.11424012917629342, 32'sd-0.13212512364943496, 32'sd0.01451685766739067, 32'sd0.0426773391686469, 32'sd1.0577235694145982e-121, 32'sd2.5386656372390023e-124, 32'sd-1.040276434379248e-124, 32'sd0.002494262915887243, 32'sd-0.06823869195481959, 32'sd0.1140217065563652, 32'sd0.07526037427107705, 32'sd-0.02953349404406909, 32'sd-0.00390613798734157, 32'sd0.012892104587563737, 32'sd-0.06565866738591633, 32'sd-0.011853242435129134, 32'sd-0.014708334739864593, 32'sd-0.01433125989568823, 32'sd0.04079769721612083, 32'sd-0.06159410954309708, 32'sd-0.04736649570685052, 32'sd0.033909626698676226, 32'sd0.04347630629998271, 32'sd0.0223187721495191, 32'sd-0.02096734088877137, 32'sd-0.06695053347426047, 32'sd-0.20055748675273663, 32'sd-0.06013748974253262, 32'sd-0.06473519770262261, 32'sd-0.05828391648351364, 32'sd-0.08930925007366762, 32'sd-0.04714302704046019, 32'sd8.349586348430501e-128, 32'sd2.7066768179194987e-118, 32'sd3.0673610186090494e-120, 32'sd0.025258960723948676, 32'sd0.016921199588873607, 32'sd0.034415709548063805, 32'sd0.04206612982726869, 32'sd0.06091780085185494, 32'sd-0.03527602546653375, 32'sd-0.03317597615545614, 32'sd-0.05802514066172307, 32'sd0.0702439527956827, 32'sd0.009555294839016779, 32'sd0.003011714127232169, 32'sd-0.02584506220994238, 32'sd-0.1026764094277249, 32'sd0.024908343881147352, 32'sd0.17588674380994956, 32'sd0.12142421531034753, 32'sd0.04434833001996123, 32'sd-0.05287299694790256, 32'sd-0.039668018680974027, 32'sd-0.20133701022234884, 32'sd-0.022120808378512675, 32'sd0.0021540263007605513, 32'sd-0.008811042525462151, 32'sd0.02259950406505506, 32'sd-0.019892961516803788, 32'sd1.5998719293680003e-124, 32'sd1.1978487151778057e-125, 32'sd2.088527169266794e-117, 32'sd-6.49508462902838e-117, 32'sd-0.041153924817800266, 32'sd-0.0624096494959056, 32'sd-0.09181779133383992, 32'sd0.04179956346552513, 32'sd0.19110796485785736, 32'sd0.03312526958946505, 32'sd0.024069885405981654, 32'sd-0.014507784436327267, 32'sd-0.06525221997874611, 32'sd-0.05948036017826212, 32'sd0.16705393718448824, 32'sd0.012565091716983614, 32'sd-0.045930822318606616, 32'sd0.051730337743985354, 32'sd0.07512606192969604, 32'sd-0.009998695611975543, 32'sd-0.001723966549910332, 32'sd-0.022847087346233353, 32'sd-0.08977816252558812, 32'sd0.0671592721514234, 32'sd0.03978006701957332, 32'sd-0.022970698931115405, 32'sd-0.00395936768431105, 32'sd4.9092692809175006e-120, 32'sd-3.1922539998268663e-119, 32'sd-6.7687589287401815e-124, 32'sd2.0471326974722576e-124, 32'sd-3.90271626997293e-116, 32'sd1.5658960238891723e-125, 32'sd-0.08776293795439918, 32'sd0.025518114759200232, 32'sd0.006641448357399528, 32'sd-0.07692815670957104, 32'sd-0.1121996616925034, 32'sd-0.039397886120653335, 32'sd0.010844209383573658, 32'sd0.08993536641169926, 32'sd-0.027933048685676285, 32'sd0.029123249082317337, 32'sd0.0055044329802887565, 32'sd-0.02599438753214766, 32'sd0.013188822378247216, 32'sd-0.04972209556640978, 32'sd0.08252730655910001, 32'sd-0.0685618186861817, 32'sd-0.07778411240849797, 32'sd-0.045206057422537735, 32'sd-0.03040216158992981, 32'sd-0.086359290635071, 32'sd4.235991759533093e-123, 32'sd5.892652529236034e-124, 32'sd1.0394508529106024e-120, 32'sd7.872213359391296e-123},
        '{32'sd-5.263926889808709e-115, 32'sd-8.24293090874901e-117, 32'sd-3.13646715000778e-123, 32'sd1.1249466390369564e-125, 32'sd5.369750603848782e-126, 32'sd-3.0884463375683036e-116, 32'sd5.916718489689415e-124, 32'sd-9.955040758127744e-124, 32'sd1.2526866760974636e-122, 32'sd1.0788330141206058e-125, 32'sd-9.452197410797237e-125, 32'sd-4.115196726103565e-115, 32'sd-0.0551092127226398, 32'sd0.04409896104405732, 32'sd0.02982060523066259, 32'sd-0.038230310738363735, 32'sd-1.2435384910182725e-117, 32'sd-7.689407655335075e-126, 32'sd8.123288321721642e-121, 32'sd-2.031666108635048e-117, 32'sd8.161436996900524e-117, 32'sd3.993655795280269e-116, 32'sd7.373959123592324e-127, 32'sd-1.0155986541842356e-124, 32'sd-3.3664685644502844e-122, 32'sd-5.882363567005767e-126, 32'sd1.8026165095095595e-123, 32'sd3.161705761963288e-123, 32'sd-1.132282558309215e-119, 32'sd1.472487116226112e-125, 32'sd-3.076698703060799e-121, 32'sd3.2862049468954684e-126, 32'sd-0.03160547520526079, 32'sd0.004854333096918809, 32'sd0.03715858493575159, 32'sd-0.01957994254446379, 32'sd-0.07197228406637599, 32'sd0.07478620787987279, 32'sd0.0545041054819804, 32'sd-0.0294364273086644, 32'sd-0.029377980573248766, 32'sd-0.1263917085856154, 32'sd-0.02933194134809297, 32'sd0.00278982832907289, 32'sd0.02439625054728296, 32'sd0.029605503040192185, 32'sd-0.008169386939807954, 32'sd-0.0010343796924234924, 32'sd-0.016704869941440995, 32'sd0.03554297512954272, 32'sd0.08777112663828027, 32'sd0.024209858672025953, 32'sd3.3605676464929984e-120, 32'sd-3.0019475983791758e-120, 32'sd2.0108860948320745e-126, 32'sd-8.81868105137292e-122, 32'sd4.060830755119979e-127, 32'sd5.156798484694313e-124, 32'sd0.060889993152136584, 32'sd0.04745618885317919, 32'sd0.011917708945885024, 32'sd0.00016411807817929368, 32'sd0.024090230622358006, 32'sd-0.011733804315747472, 32'sd0.005114697479965163, 32'sd-0.09039757185141069, 32'sd-0.05029398246937462, 32'sd0.03933777142992332, 32'sd0.06150974205768643, 32'sd0.022381240116456976, 32'sd-0.05944976707113393, 32'sd-0.032112718086731974, 32'sd0.01895800030864601, 32'sd0.01472312760653399, 32'sd-0.017811547397850513, 32'sd0.11395846468778012, 32'sd-0.0034732925368447308, 32'sd-0.06882528271727185, 32'sd-0.06599499592201212, 32'sd0.00902761773267355, 32'sd0.019809018574437155, 32'sd0.08645532528214259, 32'sd1.076176561327363e-124, 32'sd1.166702432760019e-115, 32'sd2.750628909049046e-119, 32'sd3.424395126074099e-114, 32'sd-0.06403836662931596, 32'sd0.06643678160223834, 32'sd-0.03736870365155746, 32'sd-0.014536022652842758, 32'sd-0.12289902692377101, 32'sd-0.13161457053495848, 32'sd-0.11843850978689117, 32'sd-0.09342247309478707, 32'sd-0.007040853369730223, 32'sd-0.032165019783435736, 32'sd0.08377357577486012, 32'sd-0.12029196184037627, 32'sd0.08316161077652362, 32'sd-0.13756130670698485, 32'sd-0.054719558154062924, 32'sd-0.020382386983614165, 32'sd-0.14610694907217284, 32'sd-0.06303704408489158, 32'sd0.022978275846314185, 32'sd0.012512495983399858, 32'sd-0.005175251763165415, 32'sd-0.07535440457660744, 32'sd-0.0670926945494857, 32'sd-0.11640136061475076, 32'sd-0.01290833107715935, 32'sd-8.749754300045531e-119, 32'sd8.010477264792291e-122, 32'sd0.0652095960592489, 32'sd0.0436257364035775, 32'sd0.012519611548992138, 32'sd0.04468770685813488, 32'sd0.07093608832014697, 32'sd-0.028404611089911817, 32'sd-0.09208535801752428, 32'sd-0.030121181439916697, 32'sd-0.08015356568689395, 32'sd-0.05400471152840516, 32'sd-0.1123743996920566, 32'sd-0.037293186728734405, 32'sd0.0207892752874982, 32'sd-0.06430302868890837, 32'sd-0.0028965439960909754, 32'sd-0.18132815838624763, 32'sd-0.022724078534510892, 32'sd-0.1848942985154906, 32'sd-0.046839101928941224, 32'sd-0.011233561671051847, 32'sd-0.0673199042420611, 32'sd-0.039868288261761954, 32'sd0.012462260750859568, 32'sd0.08398693682129732, 32'sd0.005519042141686691, 32'sd0.02562328663622383, 32'sd-0.028087523187153948, 32'sd-2.30449939747056e-116, 32'sd0.07587947808702851, 32'sd-0.045693593257833016, 32'sd0.09572642976268475, 32'sd0.0591641070027313, 32'sd-0.07712943509289184, 32'sd0.0206801124580954, 32'sd0.03630379549543165, 32'sd0.01912450840263124, 32'sd-0.02409876471338087, 32'sd-0.020502837242429676, 32'sd-0.11359025528308479, 32'sd-0.007113597504050421, 32'sd-0.026398808325642457, 32'sd-0.034492146788900106, 32'sd0.05613037644472739, 32'sd-0.05219821281611972, 32'sd-0.12630435049601887, 32'sd-0.11590453188959486, 32'sd-0.08918163848211794, 32'sd-0.05421360881377214, 32'sd-0.09748206037280385, 32'sd-0.03880961751918176, 32'sd-0.14542719602404436, 32'sd-0.09862802115780385, 32'sd-0.07355298782236601, 32'sd-0.06798236083069333, 32'sd0.009719758923591441, 32'sd1.9131651713890361e-121, 32'sd0.03368271980788151, 32'sd0.034677987943635025, 32'sd-0.12221218994389615, 32'sd-0.04558600972792653, 32'sd-0.04937253086481022, 32'sd0.025249939233799826, 32'sd-0.11090608587720174, 32'sd-0.0831700350069509, 32'sd-0.06464867620000855, 32'sd-0.1489193410079738, 32'sd-0.03915970843618824, 32'sd0.01641361622585587, 32'sd-0.053000904806274916, 32'sd-0.02149949152610375, 32'sd-0.0627109580625437, 32'sd-0.13429950071870478, 32'sd-0.14089867588849062, 32'sd-0.058362761451175485, 32'sd-0.20577851224486296, 32'sd-0.09280983991102693, 32'sd-0.04721178714612366, 32'sd0.01674743512818699, 32'sd0.06086858191248344, 32'sd-0.1562529420799832, 32'sd-0.19638923868146674, 32'sd-0.05798913814462729, 32'sd-0.033872229769849174, 32'sd0.03665809431650155, 32'sd-0.00754285517766876, 32'sd-0.10781307511659634, 32'sd0.0384249920993479, 32'sd0.0033240086626030404, 32'sd0.004985990091819301, 32'sd-0.024476459968210802, 32'sd-0.016171320904961407, 32'sd-0.18045834641159275, 32'sd-0.17985282198472055, 32'sd-0.10040678725797697, 32'sd-0.06613049702974498, 32'sd-0.1083318243284266, 32'sd-0.028993267614593202, 32'sd-0.2101785197852157, 32'sd-0.059180352023720906, 32'sd-0.026315961583062732, 32'sd0.05284901320930335, 32'sd0.02093912077610014, 32'sd-0.045605819306523465, 32'sd-0.05337852698680822, 32'sd0.05257072357041439, 32'sd-0.03904933782282619, 32'sd0.014803647384092282, 32'sd-0.020350667488700385, 32'sd-0.06304575269583725, 32'sd0.0013583238020505488, 32'sd0.08964090509304064, 32'sd-0.046142093165598794, 32'sd-0.0677143550130433, 32'sd0.08572882980619997, 32'sd-0.02976235591844916, 32'sd0.009162318170285413, 32'sd-0.0635262587539342, 32'sd-0.03647689750805537, 32'sd0.035976875292399964, 32'sd-0.0630908972489639, 32'sd-0.10422754305810632, 32'sd-0.10036365969368591, 32'sd-0.05550533860666681, 32'sd-0.05145223428882168, 32'sd-0.07166647426340658, 32'sd-0.058379105052765466, 32'sd-0.006250607452206301, 32'sd0.0774096757221699, 32'sd0.13280934870423827, 32'sd-0.014653932072227873, 32'sd-0.12065127115851695, 32'sd-0.08523391348662862, 32'sd-0.07359142798634327, 32'sd0.0303454710942952, 32'sd-0.05567868011636601, 32'sd0.10766608077363242, 32'sd-0.01982555802876622, 32'sd0.07831924075649052, 32'sd-0.003560027914161654, 32'sd0.02603339859972843, 32'sd-0.009363443404526375, 32'sd0.0616653617994965, 32'sd-0.014842826059902997, 32'sd-0.025413379439012503, 32'sd-0.10137534999779023, 32'sd0.016272950215314663, 32'sd0.009540277390660719, 32'sd-0.09599575188479742, 32'sd-0.13068151711116055, 32'sd-0.030645251285639493, 32'sd0.05369876839501573, 32'sd-0.03666085562162158, 32'sd-0.03361068782832972, 32'sd-0.11991543777604227, 32'sd0.0010133110294637381, 32'sd0.08124750393106156, 32'sd0.08577541516798358, 32'sd0.16052088397458564, 32'sd0.09575858079846686, 32'sd-0.0035677667253250916, 32'sd-0.08871212983961049, 32'sd-0.08954416131641556, 32'sd0.03472378211162437, 32'sd0.0956941192396265, 32'sd0.0324296209689417, 32'sd0.02367300481190952, 32'sd0.0443707285059434, 32'sd-0.019845015102989357, 32'sd0.03983375721993836, 32'sd0.08729326779255485, 32'sd0.022712627650094276, 32'sd0.0645366359785258, 32'sd-0.019674360866822515, 32'sd-0.009293433850779425, 32'sd-0.039186289860936634, 32'sd-0.11289239860169442, 32'sd0.0571566634258872, 32'sd0.036437257561506266, 32'sd0.10553838639412776, 32'sd-0.07417284743480378, 32'sd-0.02456999796603894, 32'sd0.030354983730509485, 32'sd0.1707261272517961, 32'sd0.14586926285638024, 32'sd0.08611004316889145, 32'sd0.15633857719279173, 32'sd0.16146941265256798, 32'sd-0.04902009178290462, 32'sd-0.10895394468120449, 32'sd-0.1832307042075823, 32'sd-0.0505807293410299, 32'sd0.018457806205679196, 32'sd0.05196753072172059, 32'sd-0.05263217702225185, 32'sd-0.08603820803151185, 32'sd-0.04770748071136164, 32'sd0.0899940240617564, 32'sd0.13054134723999875, 32'sd0.022235941887248055, 32'sd-0.06639886461062748, 32'sd-0.06735424780114103, 32'sd0.08786962034007074, 32'sd0.038881220041316465, 32'sd-0.02498615713102381, 32'sd-0.00031419865941755725, 32'sd-0.06379174235806523, 32'sd0.021727563898401168, 32'sd0.11066652570926394, 32'sd0.0027366124247201026, 32'sd-0.11971089168656435, 32'sd-0.05815270222659133, 32'sd0.12760916410922454, 32'sd0.10283297552931564, 32'sd0.23300657171967878, 32'sd0.10480927592464923, 32'sd-0.0024052933444454307, 32'sd0.041076688169387914, 32'sd-0.010410556407955001, 32'sd-0.015050138808315449, 32'sd-0.04577090855448951, 32'sd-0.004663817353553893, 32'sd-0.061003570305883825, 32'sd-0.002843618708759866, 32'sd0.07102156196002596, 32'sd0.017113753405684842, 32'sd0.012874319433749998, 32'sd0.025055324625148635, 32'sd0.01585420467137763, 32'sd-0.106393613448076, 32'sd0.0708042488508493, 32'sd-0.02102447402903246, 32'sd0.03247266041306938, 32'sd0.07133630471441138, 32'sd0.08897146347548754, 32'sd0.11647312614102898, 32'sd0.12093021025289054, 32'sd-0.07507870181328552, 32'sd-0.11464705376019231, 32'sd-0.021551775863381015, 32'sd-0.0062597369601038785, 32'sd0.004687606047509404, 32'sd0.07589206074931071, 32'sd0.17326730613780653, 32'sd0.029870175091613493, 32'sd-0.05129287738256729, 32'sd0.0615073578561074, 32'sd-0.06894540562140063, 32'sd0.0328098794855822, 32'sd0.040601933047221775, 32'sd-0.036634030137519244, 32'sd0.016420093916930927, 32'sd0.0349124888377658, 32'sd0.03174779133445272, 32'sd-0.017864974460960758, 32'sd-0.016315854902561953, 32'sd0.03306067665314339, 32'sd0.004337859141504834, 32'sd0.05548902580433976, 32'sd0.04525538096233613, 32'sd0.06952244866657287, 32'sd-0.05802030315538263, 32'sd0.018742217121913613, 32'sd0.13141010103051579, 32'sd0.13661483725593648, 32'sd-0.02114853471633469, 32'sd-0.09441457305045918, 32'sd-0.05219319273331733, 32'sd-0.07768862254476329, 32'sd0.16307860584663333, 32'sd0.1543720854443496, 32'sd0.18451578134049315, 32'sd0.013859207840421823, 32'sd0.03917231302681227, 32'sd-0.014944374528228386, 32'sd0.0704052687237586, 32'sd-0.0626807051367687, 32'sd0.0432299544454946, 32'sd0.039587179268236614, 32'sd-0.040473771245328694, 32'sd-0.04448614653421319, 32'sd-0.04555469230824873, 32'sd-0.013614203905023436, 32'sd-0.05747037046328634, 32'sd-0.09412508140729595, 32'sd-0.020304688496701234, 32'sd0.07934612427283566, 32'sd0.05629771834980753, 32'sd-0.044524924681501175, 32'sd0.1132851229760029, 32'sd-0.00386116457396437, 32'sd-0.013004051660099195, 32'sd0.0622289263364848, 32'sd-0.08614476923919341, 32'sd-0.07008815195561718, 32'sd0.0848547340891139, 32'sd0.039226608800046796, 32'sd0.2531251452371165, 32'sd0.12619578854693128, 32'sd0.2187275175969397, 32'sd0.04010999289928234, 32'sd-0.12083190558211665, 32'sd-0.08643436287419397, 32'sd-0.03308944478457015, 32'sd-0.10174550626386399, 32'sd0.09441087718901589, 32'sd-0.1080552181874344, 32'sd0.11481084291020868, 32'sd0.004190749705362977, 32'sd-0.01705857901210155, 32'sd0.05900694987171991, 32'sd0.026514943510128508, 32'sd0.09704040080320153, 32'sd0.07775221946036161, 32'sd-0.034658138216999736, 32'sd0.03717826106443337, 32'sd0.08429341638524042, 32'sd0.10006135996761994, 32'sd-0.005512736334569413, 32'sd0.035249990046265674, 32'sd0.13992138326786033, 32'sd-0.11207932283731327, 32'sd-0.1105245560750305, 32'sd0.04411248906203984, 32'sd-0.012688023708203988, 32'sd0.11365638928065176, 32'sd0.28137373542200467, 32'sd0.010382285368388347, 32'sd-0.15633745657180065, 32'sd-0.03850446238056873, 32'sd-0.015410956869005843, 32'sd-0.027196650829082365, 32'sd0.0068042318156296515, 32'sd-0.028807286375963085, 32'sd0.07633472963694517, 32'sd-0.04789772284221013, 32'sd0.04809778137143213, 32'sd-0.03007040636347464, 32'sd0.02242299625534227, 32'sd-0.0539314648736927, 32'sd-0.06645520556028625, 32'sd0.07836002169152632, 32'sd-0.0601290420243181, 32'sd0.08206059997308253, 32'sd0.06567596500027327, 32'sd0.14191136186701905, 32'sd0.08555180564108464, 32'sd0.10301166613051127, 32'sd0.09345463879653276, 32'sd-0.16798181278915744, 32'sd-0.2131426897682306, 32'sd-0.06460985191783837, 32'sd0.06834224208675964, 32'sd0.24327630735501685, 32'sd0.13071672284194502, 32'sd-0.08062811822390721, 32'sd-0.14173811213099832, 32'sd-0.09965287451229712, 32'sd-0.07013360348827337, 32'sd-0.0365517809205508, 32'sd-0.1266804536779932, 32'sd-0.09866014268242741, 32'sd0.039004963531570375, 32'sd-0.045397876597541575, 32'sd-1.479152378559295e-125, 32'sd0.06599608208497669, 32'sd0.07876376018952666, 32'sd-0.13198676241811683, 32'sd0.03853717637519005, 32'sd-0.008873748391999553, 32'sd0.08103484562334765, 32'sd0.017592681538277505, 32'sd0.07267290531653538, 32'sd0.17808726334447023, 32'sd0.0811646734311074, 32'sd0.17537612339313455, 32'sd-0.012483921104002378, 32'sd-0.06656922073600485, 32'sd-0.04193682116812234, 32'sd0.1670419534025754, 32'sd0.10599880084825912, 32'sd0.012910470131574774, 32'sd0.07690808202026968, 32'sd-0.052350071746282006, 32'sd-0.16042328674603393, 32'sd-0.061061921976369365, 32'sd-0.018186229018094434, 32'sd0.024031193589931873, 32'sd-0.028993906565085034, 32'sd0.0030803758608995164, 32'sd0.06208937080193523, 32'sd-0.023052772170821488, 32'sd-0.06921502335817604, 32'sd-0.03944111131275594, 32'sd0.042293615978515886, 32'sd-0.06893016337830422, 32'sd-0.020361335675801184, 32'sd-0.08259772222352364, 32'sd-0.03962551001599827, 32'sd0.05568713816985873, 32'sd0.16581025597783666, 32'sd0.11330898190274415, 32'sd-0.018071976292825497, 32'sd0.033911722841252497, 32'sd-0.04758347937533762, 32'sd-0.11189772332314553, 32'sd0.05076394932457521, 32'sd0.0991542906018735, 32'sd-0.00300984515701971, 32'sd-0.04484760403501851, 32'sd-0.035464872343652754, 32'sd-0.0679086018588768, 32'sd-0.114750497038665, 32'sd-0.1132042985112277, 32'sd-0.021019053558625603, 32'sd0.04540782598374374, 32'sd-0.14684643601139816, 32'sd0.07653511196124771, 32'sd-0.047309023419239045, 32'sd-0.05231388291438817, 32'sd0.0033657510147295316, 32'sd0.007731596545178209, 32'sd0.03936120669814466, 32'sd0.07300342890442398, 32'sd0.030128113231028, 32'sd-0.03809158928663128, 32'sd-0.039628330938298706, 32'sd0.14769362890184537, 32'sd0.11098186813915135, 32'sd-0.11446750833742152, 32'sd-0.04667109861203734, 32'sd-0.02397329303557828, 32'sd-0.06457355385201051, 32'sd-0.126118368433454, 32'sd-0.05821298223171111, 32'sd0.030977026110510106, 32'sd-0.15531294152786354, 32'sd0.003375665191289512, 32'sd-0.05809048492091402, 32'sd0.04831312570558538, 32'sd-0.08537495211020113, 32'sd-0.006210592133695408, 32'sd-0.01923145867740314, 32'sd-0.10566529764310349, 32'sd-0.03791739320648553, 32'sd0.06988180710594201, 32'sd-0.0826900540364695, 32'sd0.09208242727465893, 32'sd-3.287318264752704e-120, 32'sd-0.019763954991611748, 32'sd0.049048463791466275, 32'sd0.02154677953239834, 32'sd0.01374715006746928, 32'sd-0.03454240739392816, 32'sd-0.057389901659938417, 32'sd0.05853106897083664, 32'sd-0.10973007608358333, 32'sd-0.1744044390935668, 32'sd-0.07263771053810814, 32'sd-0.09990597060337075, 32'sd-0.020708695468597424, 32'sd-0.05647121861041701, 32'sd-0.12855110027175995, 32'sd-0.2264404787188142, 32'sd-0.06158820202088788, 32'sd-0.019750643977779207, 32'sd0.039159790724173235, 32'sd-0.051936529078285394, 32'sd-0.058309283655944136, 32'sd0.013046286082470231, 32'sd-0.04567359426484543, 32'sd-0.025244862182556844, 32'sd0.02772399670690892, 32'sd-0.007941085229918014, 32'sd-0.05898208796284483, 32'sd0.03236939773097875, 32'sd-0.0063849920832099605, 32'sd0.03780759206596789, 32'sd-0.023748027977180015, 32'sd-0.014708391722865718, 32'sd-0.03744824967114816, 32'sd0.13130584556072955, 32'sd0.01065586514557806, 32'sd-0.024993853412654126, 32'sd-0.06984340769571148, 32'sd-0.061808767994283594, 32'sd-0.12911916448260738, 32'sd-0.14396900527496398, 32'sd-0.08015667661387452, 32'sd-0.12544463990541593, 32'sd-0.14273832299755326, 32'sd-0.19793614786642688, 32'sd-0.039098669711479565, 32'sd-0.04027960444339744, 32'sd-0.10585977852706754, 32'sd0.09051864532887978, 32'sd-0.005739725669075579, 32'sd-0.04209927957855819, 32'sd0.05872942912669139, 32'sd-0.0049804800900627956, 32'sd-0.003615560736713647, 32'sd0.06095964998773856, 32'sd0.05302005250214482, 32'sd0.05399655144841009, 32'sd0.03943809848377017, 32'sd0.0010596631922221605, 32'sd0.09951777207351895, 32'sd-0.03310071044885431, 32'sd-0.005364535098605942, 32'sd-0.003403699372518006, 32'sd0.02357848478973234, 32'sd-0.09296568305176893, 32'sd-0.18362292238157393, 32'sd-0.05610744605508335, 32'sd-0.06562581080724615, 32'sd0.02628916524126509, 32'sd-0.054470640463382444, 32'sd-0.1276970639294364, 32'sd-0.015155382286953116, 32'sd-0.09351518688055359, 32'sd-0.0652503049802693, 32'sd-0.11634985232729103, 32'sd-0.10347152447067175, 32'sd0.009820898419617018, 32'sd-0.06669866625820667, 32'sd0.04912444013798914, 32'sd0.06124060818452001, 32'sd-0.06002846557332493, 32'sd-0.021101341454105527, 32'sd0.044908129363038896, 32'sd0.005923312481234222, 32'sd0.14548348864972485, 32'sd8.421617093478989e-127, 32'sd0.03661272616407123, 32'sd-0.034157377344734896, 32'sd-0.01908198147507559, 32'sd-0.13955432441972818, 32'sd-0.1257454795677626, 32'sd-0.08811332841454698, 32'sd-0.052153123665553726, 32'sd-0.038869505272701534, 32'sd-0.01508863493817185, 32'sd0.04209990966479477, 32'sd-0.058400424354516874, 32'sd-0.036697658398952254, 32'sd-0.04874614060667324, 32'sd0.006836860369689648, 32'sd-0.039959462842219184, 32'sd-0.01547756894176529, 32'sd-0.08962644086355534, 32'sd-0.11914585605142336, 32'sd0.00749596722298069, 32'sd0.039532885868894384, 32'sd-0.002479980179871928, 32'sd0.04397440313222116, 32'sd0.037139900999988096, 32'sd0.0999260640453057, 32'sd0.005655978829883985, 32'sd-0.07538231738518818, 32'sd2.5906278386657816e-126, 32'sd3.41066987179848e-123, 32'sd1.3776266542436078e-115, 32'sd0.0019889803194092868, 32'sd-0.04965671393322106, 32'sd-0.04364129954243651, 32'sd-0.05636044901497588, 32'sd-0.15585025014239262, 32'sd-0.010110511679115817, 32'sd0.038202083407678555, 32'sd0.0021750746878813516, 32'sd-0.046755168607142086, 32'sd-0.09663857166293371, 32'sd0.002400476616652002, 32'sd0.02467964134817065, 32'sd-0.06317814246487717, 32'sd-0.07567245181590622, 32'sd0.0019095096341725352, 32'sd-0.03314171250058368, 32'sd-0.05867442529643541, 32'sd0.08715395897218892, 32'sd-0.00044721954044746424, 32'sd0.0743135989070539, 32'sd0.11330955958995276, 32'sd0.10446336502392368, 32'sd0.002533047632103832, 32'sd0.0037530664028421045, 32'sd0.05398296860215872, 32'sd-1.7271197436740438e-115, 32'sd1.2669757681576118e-124, 32'sd2.273047804790221e-122, 32'sd0.07803194742217022, 32'sd-0.07583227611713697, 32'sd-0.03355152575042925, 32'sd-0.012093763733565592, 32'sd-0.04637266787949, 32'sd-0.04926730583146873, 32'sd0.014580501539976915, 32'sd0.0036092508138385773, 32'sd-0.05944134921615302, 32'sd-0.010610947940857977, 32'sd0.025840526954149057, 32'sd-0.0677705656766706, 32'sd0.02392314390770421, 32'sd0.04479317924072936, 32'sd-0.029316796555399968, 32'sd-0.06098503900747095, 32'sd0.06255465079686474, 32'sd-0.021798281807284024, 32'sd0.07054043583005594, 32'sd0.021806234538078218, 32'sd0.0787492330841642, 32'sd-0.02707146875144971, 32'sd-0.07673280253067105, 32'sd0.0980060234644198, 32'sd-0.013016184109293154, 32'sd-1.6287548189172979e-115, 32'sd-3.8760977004588374e-116, 32'sd-8.061107194841005e-117, 32'sd2.511695612241006e-123, 32'sd0.08915103143847945, 32'sd-0.023738120272121074, 32'sd0.08391320098868615, 32'sd0.0980003489075742, 32'sd0.055731616560191065, 32'sd-0.019832619662895207, 32'sd0.030138492209600305, 32'sd-0.07835056068079975, 32'sd0.10638970684877981, 32'sd0.05157004294402406, 32'sd0.05094332162526945, 32'sd-0.04024880484726777, 32'sd0.02945888427516064, 32'sd-0.0061845104624702425, 32'sd-0.07774199142627806, 32'sd-0.025406030956928217, 32'sd-0.05041266150573462, 32'sd-0.07517713566279861, 32'sd0.025541006014886396, 32'sd-0.01856301314992299, 32'sd0.015163160030196151, 32'sd0.08260010197835906, 32'sd0.04437078449518911, 32'sd-1.0575819915692394e-121, 32'sd-8.500253087984227e-115, 32'sd1.0006652960965699e-122, 32'sd2.394138614296869e-122, 32'sd-7.004102312299173e-129, 32'sd-1.4646097280026863e-123, 32'sd0.09503445889844887, 32'sd0.05166024748786588, 32'sd0.006821045517839897, 32'sd0.05195197993672068, 32'sd-0.07529098565630239, 32'sd0.04543350831035879, 32'sd0.09034319546316058, 32'sd0.015237857265632693, 32'sd-0.012528538909810944, 32'sd0.09874573189785145, 32'sd0.013821888406244535, 32'sd0.02128495517806199, 32'sd0.03441907921168712, 32'sd-0.02877479131722105, 32'sd-0.003096589445678131, 32'sd0.06062976707338678, 32'sd0.05170160801920298, 32'sd-0.04196911691304015, 32'sd0.1257866237581155, 32'sd-0.0052955813493535545, 32'sd2.3988552452219473e-129, 32'sd-1.1949199160610653e-124, 32'sd2.0365320829009052e-129, 32'sd-5.06233137898076e-126},
        '{32'sd-3.7735319074526255e-115, 32'sd3.601170337179253e-114, 32'sd-4.2653022316177344e-123, 32'sd1.0861396543703802e-119, 32'sd9.801262863765513e-121, 32'sd-1.333605755665669e-122, 32'sd-2.083046540234263e-121, 32'sd3.554097754636047e-116, 32'sd-2.3072855259736344e-123, 32'sd-1.2429974490510821e-126, 32'sd9.538814978223286e-123, 32'sd1.2325824441155171e-123, 32'sd0.035631847526699775, 32'sd0.016057277790392625, 32'sd-0.052001825682859625, 32'sd0.00969292764756304, 32'sd8.275300512247037e-126, 32'sd1.7756767844984482e-125, 32'sd6.822982287174913e-116, 32'sd3.614992898257507e-125, 32'sd-1.0714329896853253e-119, 32'sd-1.1084266916627316e-121, 32'sd-9.344340092364044e-116, 32'sd3.426241100707322e-122, 32'sd-1.996002826699719e-117, 32'sd5.354364987419895e-118, 32'sd-9.264880165375155e-119, 32'sd3.392957528614752e-119, 32'sd-9.362298457619838e-116, 32'sd-3.7946684410092256e-122, 32'sd3.5607801752764384e-114, 32'sd1.0140970353004184e-124, 32'sd0.1139367258272079, 32'sd-0.02589062627873409, 32'sd-0.007123928929326378, 32'sd0.09184974832054332, 32'sd0.02374036470630391, 32'sd0.03784344282627861, 32'sd0.0505141905188072, 32'sd-0.0904029876326093, 32'sd-0.008657939984605411, 32'sd0.11500881294033947, 32'sd-0.006294978520597279, 32'sd0.02677247132268363, 32'sd0.05836070347770698, 32'sd0.01638544703943008, 32'sd0.10948711181491902, 32'sd-0.02740866707856906, 32'sd0.04985244668224314, 32'sd0.14868695945401578, 32'sd0.14647336919312604, 32'sd0.04728503864116639, 32'sd5.034925006538676e-124, 32'sd-4.7324083370084304e-123, 32'sd1.3970668521279631e-118, 32'sd3.851037782539609e-124, 32'sd-1.1091153773385893e-121, 32'sd5.357334031904003e-118, 32'sd0.09846108964412618, 32'sd0.0525253663823429, 32'sd0.053582035048772375, 32'sd0.013017788867702315, 32'sd-0.1074265681499867, 32'sd0.014003897902167974, 32'sd0.01184139784371571, 32'sd0.13185090273202613, 32'sd-0.0028281415000159468, 32'sd0.05105766552023713, 32'sd0.029711308203653437, 32'sd0.04598142137217764, 32'sd-0.09653314457390888, 32'sd0.005234915608072376, 32'sd0.0663539029844965, 32'sd0.14313780612526492, 32'sd0.0908933693164628, 32'sd0.072612033919204, 32'sd0.05313641502645146, 32'sd-0.01688366568625487, 32'sd0.17895394316170818, 32'sd0.09118448594150441, 32'sd0.0692777354381368, 32'sd0.19197284743954626, 32'sd3.379604517319038e-116, 32'sd8.061173820857132e-127, 32'sd3.321714214420801e-122, 32'sd-5.749448023445312e-121, 32'sd0.1438303567509534, 32'sd-0.02719442515308864, 32'sd0.06914006933990323, 32'sd-0.038851109093144855, 32'sd-0.03395026033093301, 32'sd0.0545383962831532, 32'sd0.01648162313360331, 32'sd0.0023355561946660514, 32'sd0.125927585349629, 32'sd-0.000526168073417238, 32'sd0.08430073076107737, 32'sd-0.0407032699557384, 32'sd-0.0009459490670258447, 32'sd0.050669050502402696, 32'sd0.005468500438016683, 32'sd-0.019039176845434182, 32'sd-0.07821463150895334, 32'sd-0.009729591474897884, 32'sd-0.02581999358888027, 32'sd-0.023154637529107888, 32'sd-0.05627987074492405, 32'sd0.0366727342181682, 32'sd-0.03995458459692098, 32'sd-0.025014257631661048, 32'sd0.001026635134380713, 32'sd-8.209720109004927e-120, 32'sd6.167860116822603e-124, 32'sd0.028851217750284767, 32'sd0.10703358847833985, 32'sd-0.031027865635793978, 32'sd-0.006753968808346675, 32'sd-0.18521717790009953, 32'sd-0.10196642161886461, 32'sd0.12056957661735723, 32'sd0.030747112307616436, 32'sd0.04350564000652125, 32'sd-0.012048556380901486, 32'sd-0.09772869465448704, 32'sd0.01494336037736812, 32'sd0.004618252481027651, 32'sd0.06543464073211949, 32'sd-0.021575678037186106, 32'sd-0.022847443480698552, 32'sd-0.04861869317397633, 32'sd0.05952578674665436, 32'sd0.057666245826352214, 32'sd0.009379198608883425, 32'sd-0.08228896793355565, 32'sd-0.005501990055139351, 32'sd-0.05078871831819624, 32'sd-0.0018443332121837299, 32'sd-0.057151645312262626, 32'sd0.06106211231850813, 32'sd0.08725091837816053, 32'sd1.2674009630101592e-120, 32'sd-0.02887696633758235, 32'sd-0.018726303967867248, 32'sd-0.10796957096022562, 32'sd0.05137377642359106, 32'sd0.06675115474900703, 32'sd0.01639773029566134, 32'sd-0.053857844071693535, 32'sd-0.014646023126669419, 32'sd0.005738362041858623, 32'sd-0.17258671615089585, 32'sd-0.1077099733758143, 32'sd-0.10864674750343759, 32'sd0.03235401186980588, 32'sd0.14639976618238054, 32'sd0.07916512783647713, 32'sd0.07492686628355642, 32'sd0.06803721038296627, 32'sd-0.13757491290887358, 32'sd-0.036166800544177105, 32'sd0.013761028320677895, 32'sd-0.08091791905190376, 32'sd-0.0663059652515276, 32'sd0.03701190491902043, 32'sd0.11774551654382476, 32'sd-0.03432071526751069, 32'sd-0.11315124989372245, 32'sd0.022237521559159115, 32'sd3.4523426701503065e-116, 32'sd0.09050317670186249, 32'sd0.08558920351701088, 32'sd-0.08648952533273112, 32'sd0.07507342544392917, 32'sd0.030331974341354633, 32'sd-0.037691833914016086, 32'sd0.013029492564065506, 32'sd-0.021703330796145823, 32'sd-0.10479037874099938, 32'sd-0.10669202407789855, 32'sd0.07125796040689272, 32'sd0.014061991348213123, 32'sd0.055049945143738996, 32'sd0.1669976564975726, 32'sd-0.025678158013789306, 32'sd0.01289702354886273, 32'sd-0.07136736577527793, 32'sd-0.06481943794931792, 32'sd0.013484883096423667, 32'sd-0.11392713270952799, 32'sd-0.09345160610985226, 32'sd0.037474247766040615, 32'sd-0.03270238898726068, 32'sd0.029737134568102327, 32'sd-0.13192061333354957, 32'sd0.030565023983417188, 32'sd-0.019270397080701527, 32'sd0.12935661762792597, 32'sd0.12114604903150879, 32'sd-0.03691747438508499, 32'sd0.04004160827672496, 32'sd0.0851968897507448, 32'sd0.07490841602459317, 32'sd-0.07767987101460849, 32'sd0.09047477609090829, 32'sd0.01714794854666384, 32'sd0.08180567643616417, 32'sd-0.07957492561163189, 32'sd-0.08039932823566669, 32'sd-0.05020021966922686, 32'sd-0.05483306782629195, 32'sd0.10623099068859371, 32'sd-0.09619167630211307, 32'sd-0.24463738745018754, 32'sd-0.12511156251667946, 32'sd-0.11161619518832598, 32'sd-0.162316165675372, 32'sd-0.14139642254211277, 32'sd-0.13373007971219894, 32'sd-0.04473253648641873, 32'sd-0.07087791048280971, 32'sd-0.16353814177137657, 32'sd-0.14437777751304798, 32'sd0.0022128485666493614, 32'sd0.069626413808306, 32'sd0.09339179586705636, 32'sd0.02034449127256603, 32'sd-0.03724539451258374, 32'sd-0.04240703086852082, 32'sd0.10546410682075705, 32'sd0.01908353788910511, 32'sd-0.025512559955794854, 32'sd-0.013376288322526887, 32'sd0.023236154629314137, 32'sd-0.0027795403029606184, 32'sd-0.00516646697486641, 32'sd4.882217383471513e-05, 32'sd-0.015925421301297277, 32'sd-0.09313959277958889, 32'sd-0.12112531692492774, 32'sd-0.08848255855812243, 32'sd-0.25754476148543554, 32'sd-0.3020564095575101, 32'sd-0.1955003362825758, 32'sd-0.23241093691690512, 32'sd-0.24407350079003567, 32'sd-0.017562034927470556, 32'sd-0.054822868612447416, 32'sd-0.08415859918375813, 32'sd-0.06927146311207005, 32'sd-0.0717062924945359, 32'sd0.09643426487115939, 32'sd-0.026832512888142198, 32'sd0.030545639937697457, 32'sd0.11376217358003583, 32'sd-0.09345069280830713, 32'sd0.059565037000448746, 32'sd0.06754692027629691, 32'sd0.07538988549431473, 32'sd0.006791133359992035, 32'sd0.010066721946437759, 32'sd0.052849362395612394, 32'sd-0.048838408616623884, 32'sd-0.021095506896819174, 32'sd0.024061306926431346, 32'sd0.03897005842363294, 32'sd-0.016850220633077947, 32'sd0.08083280098744018, 32'sd-0.16993729705958996, 32'sd-0.3655741448096484, 32'sd-0.13900989461346586, 32'sd-0.04469241218521941, 32'sd-0.06501573057675271, 32'sd-0.03504635470199442, 32'sd-0.012032316584784852, 32'sd-0.005240662828579973, 32'sd0.07793309827440205, 32'sd0.004494229248230324, 32'sd0.03135182918780186, 32'sd0.08793894891182508, 32'sd0.0913628799929035, 32'sd0.05719055865876513, 32'sd0.06857755869738062, 32'sd-0.02013751356313878, 32'sd-0.08221223331828652, 32'sd0.032802503027450275, 32'sd0.02986102321488767, 32'sd0.007671221170531423, 32'sd-0.033253870696019594, 32'sd-0.0465982384767763, 32'sd-0.006046550473143218, 32'sd0.05604146191891162, 32'sd0.1839299964135318, 32'sd0.0971250897135955, 32'sd0.1101924681326981, 32'sd0.17143374236229994, 32'sd-0.02525964215318636, 32'sd-0.16299021659254428, 32'sd-0.03794895995822854, 32'sd0.021550709984836297, 32'sd-0.01686716927524593, 32'sd0.10629981303262867, 32'sd0.07224068271987748, 32'sd0.1015216863498035, 32'sd0.049583148322879154, 32'sd0.10659218857670594, 32'sd0.04754505498598053, 32'sd-0.05220332572842994, 32'sd-0.08563678201267381, 32'sd0.09166935124623704, 32'sd0.04950549765768017, 32'sd-0.03902513607632688, 32'sd0.055576358116504444, 32'sd-0.010234141002594887, 32'sd-0.03173627288459905, 32'sd0.08151111835287478, 32'sd-0.05014050092702394, 32'sd-0.050827813458040376, 32'sd0.13077184346103615, 32'sd0.025821644476766156, 32'sd0.14136466792066893, 32'sd0.06128909731707228, 32'sd0.2649599241386808, 32'sd0.24262604324630616, 32'sd0.0010070522518500346, 32'sd-0.11329210266226566, 32'sd0.05969176916662708, 32'sd0.20020675285165704, 32'sd0.06458196133295324, 32'sd0.07134910674679464, 32'sd0.16175215013058702, 32'sd0.11888488823104608, 32'sd0.09081160595438857, 32'sd-0.04952223500622704, 32'sd0.01318606998631208, 32'sd-0.02895593346151167, 32'sd0.04410189410368562, 32'sd0.0472367707141899, 32'sd0.04423251530633482, 32'sd0.09454192602964544, 32'sd0.09339656928807852, 32'sd-0.00047494818444786296, 32'sd0.025803775416198514, 32'sd-0.06889847698776999, 32'sd-0.15212163171019405, 32'sd0.027524456671574726, 32'sd0.08160862164860753, 32'sd-0.08828188705115833, 32'sd0.09440143598565127, 32'sd0.19017157152047723, 32'sd0.2329756127672917, 32'sd0.20539822514472453, 32'sd-0.02190239095539121, 32'sd-0.13624159821829673, 32'sd0.047009591198508505, 32'sd0.022109808640216406, 32'sd0.09830165631613665, 32'sd0.1865763455708145, 32'sd0.09474125276749235, 32'sd0.2442121753832177, 32'sd0.13406095354098602, 32'sd-0.10288274715963772, 32'sd-0.08577850263483533, 32'sd0.08553785136961473, 32'sd0.13918438257128407, 32'sd0.08850337731710937, 32'sd0.08563255999252914, 32'sd0.04144782414029423, 32'sd0.03714237597934343, 32'sd-0.10810159939037091, 32'sd0.1397410434229348, 32'sd-0.08478344759180897, 32'sd-0.049263596858228474, 32'sd-0.06110242278409409, 32'sd-0.11223933561007148, 32'sd-0.09862600615938122, 32'sd-0.03703180364031733, 32'sd0.08544650130010666, 32'sd0.1304605299126953, 32'sd0.008527684544020402, 32'sd0.08054734077925328, 32'sd-0.010444129971889279, 32'sd0.05198007853585466, 32'sd-0.021257277760924745, 32'sd0.05333697103930622, 32'sd0.09306965844348691, 32'sd0.22760898147113337, 32'sd0.08301428517712092, 32'sd0.15421200907609667, 32'sd-0.021663778684061476, 32'sd-0.017431164592822516, 32'sd-0.00035677776974181414, 32'sd-0.03314273495128881, 32'sd0.13289301124788805, 32'sd-0.02316126888342225, 32'sd0.029379912649601363, 32'sd0.07912509373477263, 32'sd-0.10376128924653187, 32'sd-0.01080910689033077, 32'sd0.020661444749350753, 32'sd0.0012370055350992885, 32'sd-0.005789376820746528, 32'sd0.009100461967216426, 32'sd0.06385336923322926, 32'sd-0.04279510768886937, 32'sd0.09336426205848405, 32'sd-0.0004970703887429301, 32'sd0.09170152276363516, 32'sd0.09043317399867841, 32'sd0.12414056945224212, 32'sd0.01771740000524246, 32'sd0.07449695142552268, 32'sd-0.011162280777246753, 32'sd0.09057593750169878, 32'sd0.16458765433198513, 32'sd0.06623112490248931, 32'sd-0.0032966425558638227, 32'sd-0.028669680215004316, 32'sd-0.03137229473079852, 32'sd-0.09184986795383343, 32'sd-0.05560564852437025, 32'sd0.038936640923072655, 32'sd-0.006798541974640502, 32'sd0.04418602587432152, 32'sd-0.021290009607560466, 32'sd-0.058492510632934806, 32'sd-0.0669579768660537, 32'sd-0.01846383655819584, 32'sd0.11058560627331591, 32'sd0.08274303893947489, 32'sd0.004062582610531655, 32'sd0.02098649218399534, 32'sd-0.05298087098878738, 32'sd0.0023376003805066297, 32'sd0.13576927752697387, 32'sd0.15191774276842393, 32'sd0.0974663810169902, 32'sd-0.03721892984208294, 32'sd-0.015860825838059926, 32'sd0.06604411497365714, 32'sd0.043403249584129784, 32'sd0.05158905283875848, 32'sd0.07415722255228681, 32'sd0.06309502593132627, 32'sd-0.007837841076374485, 32'sd0.002618916794472587, 32'sd0.041521923513766275, 32'sd-0.0032478056757973372, 32'sd0.04050231739428812, 32'sd0.035819911364233584, 32'sd-0.050763063148541065, 32'sd0.02921086141044669, 32'sd0.06285509631714971, 32'sd0.01429744912655916, 32'sd0.07150707995009419, 32'sd0.09100965572463895, 32'sd0.06578913651794507, 32'sd0.06562087317741434, 32'sd-0.06471765121123375, 32'sd-0.029556259628668292, 32'sd-0.0637405769922881, 32'sd-0.025030815012529597, 32'sd-0.023800860265384135, 32'sd0.10797255222058097, 32'sd-0.028153923593963254, 32'sd-0.16106952789735351, 32'sd-0.09609219796402084, 32'sd-0.03225469260973946, 32'sd-0.08150636042491029, 32'sd0.0008655805665560932, 32'sd0.02802588208471755, 32'sd-0.08654230612479452, 32'sd-0.06895748892430834, 32'sd-0.020500884559379984, 32'sd-0.053232664164581514, 32'sd0.003870255688336928, 32'sd-0.05867315534325025, 32'sd1.0525572558162983e-124, 32'sd0.06526636070877785, 32'sd0.037708262418312155, 32'sd-0.05230622169760629, 32'sd0.03333975710199562, 32'sd0.017097019242178508, 32'sd-0.12414752551416053, 32'sd-0.10566655315507359, 32'sd0.053912234992433965, 32'sd-0.022224895946653157, 32'sd-0.056770491339996974, 32'sd-0.04666785853548648, 32'sd-0.09387308724149103, 32'sd0.01705235994805887, 32'sd0.07381195974462225, 32'sd-0.016983373032807482, 32'sd-0.08071839773459512, 32'sd-0.05728936585108071, 32'sd0.010628089630120297, 32'sd0.04001302201851729, 32'sd0.029121516601711188, 32'sd0.005248451519787345, 32'sd-0.034675167569315095, 32'sd-0.12523865928987216, 32'sd-0.11904808046407979, 32'sd-0.08339353454844993, 32'sd0.06444736210294769, 32'sd-0.027528850237376168, 32'sd-0.035999754062249124, 32'sd0.025929592678542612, 32'sd-0.016761970664275015, 32'sd-0.004486189009114177, 32'sd-0.001484259834461244, 32'sd0.017634019374709133, 32'sd-0.13012238823316294, 32'sd-0.15840933036139623, 32'sd-0.033209912907726444, 32'sd0.0289457710050634, 32'sd-0.13676228129085213, 32'sd-0.09152966028726743, 32'sd-0.06288355522242083, 32'sd0.1157358276398045, 32'sd0.05504718482849408, 32'sd-0.05690972829870862, 32'sd-0.16099457167978604, 32'sd0.00841111974812831, 32'sd0.04374751222647906, 32'sd0.023513051494314863, 32'sd0.04824658319949739, 32'sd-0.09679462932709311, 32'sd-0.15109597992567195, 32'sd-0.23685449636848527, 32'sd-0.1346457870628201, 32'sd-0.0019963963687040526, 32'sd0.005183629764722213, 32'sd0.05522192110169569, 32'sd0.05777747395166728, 32'sd-0.047277299114947935, 32'sd0.008840822224083916, 32'sd-0.05323026708302517, 32'sd0.06505896510632984, 32'sd-0.027094225090068935, 32'sd-0.08745844233098661, 32'sd-0.13768078987444815, 32'sd0.03829637237068502, 32'sd-0.048230334727928176, 32'sd-0.13942494908241748, 32'sd-0.13076949818641825, 32'sd-0.12386049903998494, 32'sd0.06899002045280003, 32'sd0.0613688461415468, 32'sd0.014898488355516755, 32'sd-0.03543153549727152, 32'sd-0.07488301174879325, 32'sd0.05679462410505542, 32'sd-0.04685276671225205, 32'sd-0.09032457595605448, 32'sd-0.09681808525905411, 32'sd-0.11820434961931402, 32'sd-0.08441408544477996, 32'sd-0.11622479860350744, 32'sd-0.026586969973377172, 32'sd0.07465276659014426, 32'sd0.05549478413722039, 32'sd3.709963481831336e-122, 32'sd-0.015312787632045487, 32'sd-0.06548949436510769, 32'sd0.07838716486201663, 32'sd0.2019684906088062, 32'sd0.07112356024572072, 32'sd-0.052511633005839164, 32'sd-0.09222700451747505, 32'sd0.004170822853859181, 32'sd-0.05508381512241742, 32'sd-0.13963669420858368, 32'sd-0.04790495728232718, 32'sd0.015692683594940467, 32'sd0.00982918932845471, 32'sd0.037529809185229766, 32'sd0.16685350039693825, 32'sd0.07179627404405511, 32'sd0.06712754308210739, 32'sd0.03356883078257237, 32'sd-0.05982368864530212, 32'sd-0.07598668461069065, 32'sd-0.0866028787607487, 32'sd-0.19407681813193356, 32'sd-0.11527114408572846, 32'sd0.013248440490990986, 32'sd0.03914775392963039, 32'sd0.01615540295339518, 32'sd-0.014563361391568382, 32'sd0.02580995118112919, 32'sd-0.01419231514944373, 32'sd0.055734813277690316, 32'sd-0.1540362439175559, 32'sd-0.02523126588157121, 32'sd0.002184037469599909, 32'sd0.0740900434849424, 32'sd-0.06596888680647776, 32'sd-0.0716738669229773, 32'sd0.09220887375311981, 32'sd0.014352059321664081, 32'sd0.06547526666245976, 32'sd0.056920397926997164, 32'sd0.06480853531099422, 32'sd0.017223720367056168, 32'sd0.07625058578790518, 32'sd0.1877318621358463, 32'sd0.12700116844885637, 32'sd0.014684023376395829, 32'sd0.023142926791369468, 32'sd0.09037268275913034, 32'sd-0.062475920567519085, 32'sd0.002434607232861874, 32'sd-0.05583844725599934, 32'sd-0.06807884966282886, 32'sd-0.0009081391618762182, 32'sd0.06593850441202687, 32'sd0.09480305570039461, 32'sd0.10363718814235429, 32'sd0.06715565919275662, 32'sd-0.05809581795046292, 32'sd-0.09629696931311106, 32'sd0.0190697924458556, 32'sd-0.05358451218656797, 32'sd-0.07858439018713825, 32'sd0.016941839806750375, 32'sd-0.09377896305303406, 32'sd0.026273998964473376, 32'sd-0.057114385362866324, 32'sd0.053118277352739135, 32'sd-0.012607811213418887, 32'sd0.04605419044949579, 32'sd0.01063637729150863, 32'sd0.007946407466005681, 32'sd0.1982751874155077, 32'sd-0.009740368984477756, 32'sd0.10208865168043489, 32'sd0.0283960804355046, 32'sd0.02985797564673567, 32'sd-0.06875647827772333, 32'sd-0.09631258314943568, 32'sd-0.020650633498863938, 32'sd0.06621014672719663, 32'sd-0.0514654809457874, 32'sd-0.007381532324248058, 32'sd0.08239450071753389, 32'sd-5.938399413668201e-122, 32'sd0.09614622237497612, 32'sd0.10086506780732106, 32'sd0.021900774104700024, 32'sd0.016493607987587172, 32'sd0.018808372187294628, 32'sd0.0517721569028295, 32'sd-0.09465819390040667, 32'sd-0.11033816825531352, 32'sd-0.014823186978207472, 32'sd-0.07433771552695138, 32'sd-0.22496419341896406, 32'sd-0.0008216017642381549, 32'sd-0.025662122149424964, 32'sd0.11318311942008472, 32'sd-0.012904282623773966, 32'sd0.019012813327659556, 32'sd0.024287099396097904, 32'sd0.017555804901851005, 32'sd0.029815435248778315, 32'sd0.07656684622174023, 32'sd-0.013664527781580255, 32'sd-0.10510488530426706, 32'sd-0.001115640842115657, 32'sd-0.06494169752806582, 32'sd0.017008249682532946, 32'sd-0.003275833107684725, 32'sd-9.024520229578544e-118, 32'sd1.6115866928791918e-127, 32'sd1.07049065987105e-124, 32'sd-0.031872556640553724, 32'sd0.016675740103226352, 32'sd0.060165988248505095, 32'sd0.11323694440740002, 32'sd0.05105200846242504, 32'sd-0.005042780979993035, 32'sd-0.010399734633867468, 32'sd-0.04502779933087905, 32'sd0.005941497562693645, 32'sd0.0014161903444864026, 32'sd-0.08009103314260133, 32'sd-0.021347523366609195, 32'sd-0.0437961396475381, 32'sd-0.010196569467494292, 32'sd-0.06849780346034394, 32'sd0.0594461157795195, 32'sd0.015009620126608602, 32'sd-0.03412144956554748, 32'sd-0.01602341696942844, 32'sd-0.05554253759572224, 32'sd-0.10888729490675736, 32'sd-0.010887624740805707, 32'sd0.024804775370612018, 32'sd0.0325849371312151, 32'sd-0.021994484460745943, 32'sd-7.892822707475099e-115, 32'sd-2.615360397056592e-120, 32'sd1.0454453325099694e-120, 32'sd0.0600947180297528, 32'sd0.14558735995898478, 32'sd-0.041870259674462076, 32'sd-0.07527943224172165, 32'sd0.10266737048996853, 32'sd0.0421018939651314, 32'sd-0.01758138121612645, 32'sd0.006041696374256918, 32'sd0.009017245342089752, 32'sd0.031234234816374492, 32'sd0.057432122571901834, 32'sd-0.007411942541215671, 32'sd0.047439373294279996, 32'sd-0.10974446326851812, 32'sd-0.0183879562015186, 32'sd0.1136165734897869, 32'sd0.05405643501326663, 32'sd-0.07732575384240382, 32'sd0.04938871017061973, 32'sd-0.057766704050867576, 32'sd0.07524957718735997, 32'sd0.009665444399875059, 32'sd-0.09387344322592456, 32'sd-0.07149125216640453, 32'sd0.03126407945660988, 32'sd1.4456603127940755e-120, 32'sd-9.26563869550175e-122, 32'sd-1.199300796373443e-121, 32'sd-3.960963761543877e-126, 32'sd0.14034983955604804, 32'sd-0.02305782141579001, 32'sd-0.09360490970553563, 32'sd0.03157734313494013, 32'sd-0.05552247400956251, 32'sd-0.0816275958621528, 32'sd0.1647897358840128, 32'sd0.011064427126398359, 32'sd0.08483823774804283, 32'sd0.0382022178381318, 32'sd0.11458772168150766, 32'sd-0.012264641640396071, 32'sd-0.06634915944877409, 32'sd0.03393308746735137, 32'sd0.042953199831205276, 32'sd-0.0005984884853045266, 32'sd0.08333536430887113, 32'sd-0.06701413191737571, 32'sd0.09467805309372587, 32'sd0.05361919235459927, 32'sd0.021880176169814067, 32'sd0.02590075675165748, 32'sd0.10731295429079539, 32'sd5.002571210233413e-115, 32'sd2.5976014282479808e-126, 32'sd1.8603930449033504e-117, 32'sd1.5352508936653614e-116, 32'sd3.6880872056031517e-125, 32'sd-1.98926393413611e-124, 32'sd0.15106867639065602, 32'sd0.08343620214260623, 32'sd0.07884403141126506, 32'sd0.06150149965660623, 32'sd0.10354061967073926, 32'sd-0.005078743098128188, 32'sd0.0041531533282174364, 32'sd0.08450474673559177, 32'sd0.005757436778140171, 32'sd-0.040873521692474435, 32'sd0.0337841167274075, 32'sd0.031395107828965714, 32'sd0.07389621969286082, 32'sd0.1026905804207456, 32'sd0.02090951041664565, 32'sd0.08081224266914695, 32'sd-0.025960597217125812, 32'sd0.10745399210726339, 32'sd0.09605137496554302, 32'sd0.0859545074759948, 32'sd-1.89591668628803e-125, 32'sd-5.032541517622797e-118, 32'sd6.0182261556459035e-123, 32'sd-1.0785830655729535e-124},
        '{32'sd1.2672163607471447e-121, 32'sd6.974238429150464e-115, 32'sd-5.806315212471822e-120, 32'sd-9.763359902851188e-120, 32'sd-9.548068103786497e-117, 32'sd-2.117653215629172e-117, 32'sd-6.672904812481742e-126, 32'sd1.767533898963246e-125, 32'sd2.2943405193438586e-123, 32'sd1.067728410860136e-124, 32'sd2.187591269986909e-126, 32'sd-1.8119948313364222e-126, 32'sd0.04988161622415852, 32'sd0.11565510173580343, 32'sd-0.024180204880180446, 32'sd0.1154993523905477, 32'sd7.705339040006766e-125, 32'sd-4.933674864110509e-125, 32'sd-2.8028453804522386e-125, 32'sd-8.138838066880214e-123, 32'sd1.22846541927465e-122, 32'sd-6.876712245524389e-124, 32'sd-3.0637849863674593e-121, 32'sd3.971246444218694e-124, 32'sd3.3008914371082404e-121, 32'sd6.728367600883163e-127, 32'sd1.8217058784109444e-123, 32'sd-1.1702286347074884e-119, 32'sd-1.0249044894924347e-125, 32'sd2.029094801221769e-117, 32'sd4.033210564948222e-122, 32'sd2.1622464114648235e-126, 32'sd0.020663986697537322, 32'sd-0.08787752214882517, 32'sd0.06289906029401876, 32'sd0.12505490328621005, 32'sd-0.010303415238000175, 32'sd0.025374284438280017, 32'sd0.10360893570597132, 32'sd0.008492562660914344, 32'sd0.06603660915465358, 32'sd-0.03474791056011041, 32'sd-0.09644069571374894, 32'sd0.01712291081226005, 32'sd0.041988769606888965, 32'sd0.06505165836855653, 32'sd0.06433989440430535, 32'sd0.009401978588920437, 32'sd0.06419203611461795, 32'sd0.0573048606452106, 32'sd0.07950063943835357, 32'sd-0.004324594528711608, 32'sd-2.155703071294719e-121, 32'sd1.0780640181918289e-117, 32'sd2.2895069171199546e-126, 32'sd-3.67139649583647e-129, 32'sd-8.719632850135296e-118, 32'sd1.3269362449731316e-126, 32'sd0.03250393824796849, 32'sd-0.0454287878527617, 32'sd0.02275639254810581, 32'sd0.030188771262463814, 32'sd0.08070199861939853, 32'sd0.03389714650731596, 32'sd0.12737429136630396, 32'sd0.03584243915484589, 32'sd-0.01464258643269353, 32'sd0.14337850217841622, 32'sd0.13141053178752043, 32'sd-0.00856534400264845, 32'sd-0.027741832855693028, 32'sd0.08175749996909469, 32'sd-0.0034830193670741935, 32'sd0.0898638856263074, 32'sd-0.011252096681438086, 32'sd0.00487208402442575, 32'sd-0.011986714904348912, 32'sd0.03850445923566379, 32'sd0.01648785191555459, 32'sd-0.032809852331784135, 32'sd0.05937360624594854, 32'sd0.10860210929089963, 32'sd7.765780901607565e-127, 32'sd-1.3155070736495076e-122, 32'sd-6.0588881464746334e-117, 32'sd3.859086430042983e-124, 32'sd0.04158938548124623, 32'sd0.07927742510479245, 32'sd0.10200819016049031, 32'sd0.11787095798799155, 32'sd0.1147156533596665, 32'sd0.12472637099550382, 32'sd0.033768245003815395, 32'sd-0.035419781131305415, 32'sd0.05880920059903524, 32'sd0.12302994400869503, 32'sd0.061566367051107844, 32'sd0.12321412274728953, 32'sd-0.008758810371086858, 32'sd-0.06201585274950294, 32'sd0.0382895511586919, 32'sd0.020429966726631364, 32'sd-0.09784333006716943, 32'sd-0.0591254250244342, 32'sd-0.04516649127978615, 32'sd0.06351334845448535, 32'sd0.04077515280719493, 32'sd0.09331214774663653, 32'sd0.09814957992564058, 32'sd0.010939168668113258, 32'sd0.09472120587735669, 32'sd2.5703215749801455e-115, 32'sd6.389359874156845e-116, 32'sd0.04403346274970991, 32'sd-0.00459046935865067, 32'sd0.0020456026747459966, 32'sd-0.012619789669227577, 32'sd0.07766274435967165, 32'sd0.10667147740341776, 32'sd0.047429315357339054, 32'sd0.034700045464679294, 32'sd-0.024289161289226844, 32'sd0.11172941473687938, 32'sd0.05793800124081187, 32'sd0.04639758007711169, 32'sd-0.043749194500998775, 32'sd0.04702094418978032, 32'sd0.008243521670807214, 32'sd0.0763738959526382, 32'sd0.04924917510944049, 32'sd0.03971892264702651, 32'sd0.03518016138127039, 32'sd0.03877989250555154, 32'sd-0.053966628388708825, 32'sd-0.04400298300081148, 32'sd0.007644438279443212, 32'sd0.02219092339127634, 32'sd-0.013284995150768756, 32'sd-0.02458900435882882, 32'sd0.0652869109165773, 32'sd4.4573595476421263e-122, 32'sd0.052005558954118326, 32'sd0.01019879189230713, 32'sd0.061308049129022185, 32'sd0.0417776772894085, 32'sd0.03155248168554654, 32'sd0.05103079092922112, 32'sd-0.10379917287016857, 32'sd-0.011096336881366296, 32'sd-0.07389529038618274, 32'sd-0.0023397633081017263, 32'sd-0.0016666111064323297, 32'sd-0.10373088236316642, 32'sd-0.10983066307899064, 32'sd-0.07747871809104682, 32'sd0.003722474809794882, 32'sd0.0130045811434353, 32'sd0.016599532538993714, 32'sd0.023680724807816314, 32'sd0.13363450187452805, 32'sd-0.006306478154044082, 32'sd-0.10824436914832068, 32'sd-0.08768776562550169, 32'sd-0.032075651300878194, 32'sd-0.0908575830977857, 32'sd-0.07299210563822162, 32'sd0.04178394540241206, 32'sd0.07747506587576618, 32'sd1.564976218038374e-120, 32'sd0.0065509331644906296, 32'sd0.015183084429226008, 32'sd0.0014990062965568817, 32'sd0.08083709047819361, 32'sd0.04290527786896577, 32'sd0.03361965471223882, 32'sd-0.055956318611071594, 32'sd-0.03521097744990667, 32'sd0.07243268689909539, 32'sd-0.0761623816137437, 32'sd0.021891287105697346, 32'sd-0.21576344808013084, 32'sd-0.16839747690305598, 32'sd-0.08617590981292478, 32'sd-0.05832631775656889, 32'sd0.058949873403565674, 32'sd0.09651487936826764, 32'sd0.10301476736040002, 32'sd0.11891913440565825, 32'sd-0.02048616048995704, 32'sd-0.05216985922201346, 32'sd-0.06283985904052702, 32'sd-0.1457224986821656, 32'sd-0.24313980817199005, 32'sd-0.09408237908044417, 32'sd0.0881044290898341, 32'sd-0.01666747005625082, 32'sd0.08303998487278709, 32'sd-0.014679062875358374, 32'sd0.0522928055971731, 32'sd0.07220492166703008, 32'sd-0.08704919451403323, 32'sd-0.03094848955368203, 32'sd-0.04729656701089399, 32'sd0.035446835394745295, 32'sd0.07118031539405187, 32'sd-0.009478957093657505, 32'sd-0.04161961140838335, 32'sd-0.14763548400925705, 32'sd-0.15694961486146697, 32'sd-0.12499169523583234, 32'sd0.07627955149020006, 32'sd-0.002772236378164128, 32'sd-0.13563493298839654, 32'sd0.02053274049898231, 32'sd0.08664126161813283, 32'sd0.07893003025268719, 32'sd-0.02320359643676857, 32'sd0.03368436777007086, 32'sd-0.0062637378046152175, 32'sd-0.03601778182369511, 32'sd0.01788405446599331, 32'sd-0.04509341376681437, 32'sd0.011523170360839172, 32'sd-0.00565337647018492, 32'sd0.05442098703040942, 32'sd0.06933497460678428, 32'sd0.0748895428181368, 32'sd-0.0007224522970353299, 32'sd-0.06472064008389086, 32'sd-0.06373838760180439, 32'sd0.02519915048551817, 32'sd-0.06819327494137821, 32'sd-0.06236225379398756, 32'sd-0.12061154584838964, 32'sd-0.0416566487844369, 32'sd-0.02837336854386333, 32'sd0.04160529369299231, 32'sd0.02273242528875743, 32'sd0.0779596336842944, 32'sd0.08674003210152358, 32'sd0.05296644735834919, 32'sd-0.03626699798700949, 32'sd-0.014695209938014894, 32'sd0.03692717277019852, 32'sd-0.028538298364159113, 32'sd-0.057282877764968286, 32'sd0.002994723869235633, 32'sd0.04154682898800855, 32'sd-0.03796293165372532, 32'sd-0.048275010360045625, 32'sd0.09813103197884072, 32'sd-0.01779130907762953, 32'sd0.044100518364160006, 32'sd-0.0907856593828218, 32'sd-0.005064038458452471, 32'sd-0.05746416094561289, 32'sd0.0465956887299281, 32'sd0.07093063098010188, 32'sd-0.008757570157134903, 32'sd-0.02775682973890054, 32'sd-0.06639743134510707, 32'sd-0.10214375945741695, 32'sd-0.12843584497415805, 32'sd-0.07615931718258627, 32'sd0.025378710275881997, 32'sd0.15791264777726058, 32'sd-0.007685598752668242, 32'sd-0.05643407298498545, 32'sd-0.09575549340140432, 32'sd-0.013424057161070205, 32'sd-0.05136678944742974, 32'sd-0.03517119860068613, 32'sd-0.0013414286981683306, 32'sd-0.06434019519303712, 32'sd0.08867613704432081, 32'sd0.08171131502736584, 32'sd0.0450756037190372, 32'sd-0.09635809380511684, 32'sd0.09346723872925886, 32'sd-0.03698772912548037, 32'sd-0.012433939073750346, 32'sd-0.012989353273308867, 32'sd0.02076680785828554, 32'sd-0.06244011147452994, 32'sd0.018613565447211305, 32'sd0.13379832169668943, 32'sd-0.01946182191355403, 32'sd-0.13932117565067914, 32'sd-0.07593486794899346, 32'sd-0.04685821565752817, 32'sd-0.10379526145495728, 32'sd-0.09662008020774154, 32'sd0.1429884114260973, 32'sd-0.016827638273109197, 32'sd-0.05240174940872271, 32'sd-0.11596274731184442, 32'sd-0.14619605234693703, 32'sd-0.10308601745288128, 32'sd-0.07099950477969234, 32'sd-0.07812484608265392, 32'sd-0.007156980070854175, 32'sd0.020770680444791675, 32'sd0.021251248999391573, 32'sd0.099252506556008, 32'sd-0.007887267911098542, 32'sd-0.04468173859547049, 32'sd0.0638945578667672, 32'sd0.018081607622018915, 32'sd-0.05576981955207603, 32'sd0.06382190761533972, 32'sd0.018510134420129797, 32'sd-0.07939223209588968, 32'sd-0.08772341762071727, 32'sd0.02350603207607581, 32'sd0.0011171012361965722, 32'sd-0.0438194820489346, 32'sd0.027674386792983327, 32'sd0.10691349113813328, 32'sd-0.12490669355829313, 32'sd0.07697681065161138, 32'sd-0.02172495425928618, 32'sd-0.05188566509869768, 32'sd-0.17028598791195462, 32'sd-0.24060965153421113, 32'sd-0.21517120336095044, 32'sd-0.06263316159162342, 32'sd-0.1094211257428457, 32'sd-0.10892103539602876, 32'sd0.11589912097911483, 32'sd0.06310651879948861, 32'sd0.08237329193573519, 32'sd-0.004620656418842819, 32'sd0.030689246509025075, 32'sd0.018648923965090526, 32'sd0.026748926901280723, 32'sd0.08255796914537453, 32'sd0.05892073127163767, 32'sd0.04785271588184123, 32'sd-0.07646078978492894, 32'sd-0.04515429559510491, 32'sd0.0771893791299261, 32'sd0.03676642313075326, 32'sd0.008665704616806668, 32'sd-0.028982464718831962, 32'sd-0.04037747377905905, 32'sd0.04919058847490068, 32'sd0.022272192219137933, 32'sd0.008476666164773607, 32'sd0.013663165195202475, 32'sd-0.04674295765395744, 32'sd-0.04479427990107792, 32'sd-0.01040674871875897, 32'sd0.00975923555707561, 32'sd0.05935886504022633, 32'sd0.10570793686921616, 32'sd-0.008196836416764134, 32'sd0.055589168113449584, 32'sd0.11501680079572323, 32'sd0.04326429207807178, 32'sd0.1240555130091401, 32'sd0.029888257927276108, 32'sd-0.005012885053991436, 32'sd-0.01926390005320586, 32'sd0.014987990300353705, 32'sd0.05427970588793793, 32'sd-0.05297897078887442, 32'sd-0.07581118247395328, 32'sd-0.05242111487301631, 32'sd0.045019214534137895, 32'sd0.07073323120674706, 32'sd-0.06276306359720948, 32'sd0.03343512180184366, 32'sd-0.032385653147555295, 32'sd0.10853619040673157, 32'sd-0.03806833179826962, 32'sd0.05499267421722002, 32'sd-0.09454644590313303, 32'sd-0.01048008450567694, 32'sd0.1223799257234378, 32'sd0.11126124395388483, 32'sd0.19636500697902123, 32'sd0.0334880219300684, 32'sd0.10007402072447158, 32'sd-0.007699682845887153, 32'sd0.07260394703403868, 32'sd0.0448837817973893, 32'sd0.16822239812150752, 32'sd0.0770857334667493, 32'sd-0.03001766316053083, 32'sd0.012772431364793224, 32'sd0.021672866843285232, 32'sd0.05785612976396351, 32'sd0.029427645826674873, 32'sd0.01991195906021909, 32'sd-0.020788574133580547, 32'sd-0.0946948406456589, 32'sd-0.0008366058330906977, 32'sd0.11021008161106005, 32'sd-0.006619798979206022, 32'sd0.0943072387556078, 32'sd0.056167252593519894, 32'sd0.09023692153369944, 32'sd0.08211740012292502, 32'sd-0.01310656367091266, 32'sd-0.08478791369548429, 32'sd-0.052525040074606795, 32'sd-0.026189153423295593, 32'sd0.2134963982874083, 32'sd0.1565263420545742, 32'sd0.0871263083352763, 32'sd-0.032434245218468154, 32'sd-0.0666288927401699, 32'sd-0.0181017147946213, 32'sd0.017841274417606686, 32'sd-0.007601657519840224, 32'sd0.06798532542617752, 32'sd-0.06554735134228194, 32'sd0.00028563642028734245, 32'sd0.001140741518313173, 32'sd0.07588857649164998, 32'sd-0.023873896637671997, 32'sd0.02409893237117763, 32'sd0.060301191594502035, 32'sd-0.09967999794325307, 32'sd-0.12287132819933258, 32'sd0.041603353498368925, 32'sd0.09068398888588236, 32'sd0.034666164000866966, 32'sd0.05652874626515269, 32'sd0.15459986169652912, 32'sd-0.008233077788055094, 32'sd-0.054930182981834996, 32'sd-0.0665824584806844, 32'sd-0.057153146018534245, 32'sd0.1206826232478222, 32'sd0.16451232533582694, 32'sd0.10472426902152603, 32'sd-0.05407885249825947, 32'sd0.0006130644545952584, 32'sd0.010485482515000337, 32'sd-0.013621838718835523, 32'sd0.05454233606687398, 32'sd-0.008023733398984705, 32'sd0.05980372270121914, 32'sd0.04627172434683864, 32'sd-0.06945614370277862, 32'sd0.05200824497180093, 32'sd0.029122716216450295, 32'sd0.03822126862806189, 32'sd0.10976171661253774, 32'sd0.05583937353770412, 32'sd-0.096854072304083, 32'sd-0.05092546117665958, 32'sd0.06509153108368033, 32'sd-0.028675724915830283, 32'sd-0.02315183299072334, 32'sd0.017553816705716135, 32'sd0.10713873602419424, 32'sd0.06838210536350427, 32'sd0.16157374062680904, 32'sd0.18450826562324235, 32'sd0.09697977767319295, 32'sd0.09214122261073973, 32'sd0.04254943982187564, 32'sd-0.03317178093423762, 32'sd-0.13309122792452352, 32'sd-0.05763154791498594, 32'sd-0.10748216572645894, 32'sd-0.06954782124042098, 32'sd-0.1287983064892454, 32'sd-0.12104538957038788, 32'sd-0.0037541150093133844, 32'sd-0.06510144659376299, 32'sd0.04104344742783776, 32'sd-0.02509370797604763, 32'sd-0.009837713919270453, 32'sd-3.1962276902538856e-119, 32'sd-0.0030848193111893906, 32'sd0.04397223835663814, 32'sd0.045239764186888284, 32'sd-0.0040283642969151275, 32'sd0.12091039410907924, 32'sd0.074490838604921, 32'sd-0.07208913038535752, 32'sd-0.037875455325829165, 32'sd-0.06773139037403632, 32'sd0.1052046469911344, 32'sd0.05415605935703057, 32'sd0.06225230100795032, 32'sd-0.03952832059512641, 32'sd-0.04373358574023463, 32'sd0.06659456449989654, 32'sd0.0012248533052638408, 32'sd-0.10650320047139802, 32'sd0.05145027070740227, 32'sd-0.051054982488050384, 32'sd-0.07057127125328705, 32'sd-0.004512435863004887, 32'sd-0.024778525825703626, 32'sd0.02992398549456501, 32'sd-0.0535073587920824, 32'sd0.09119316760255855, 32'sd-0.0675494112193576, 32'sd0.052810630100178564, 32'sd0.04502888018107247, 32'sd0.09453072325953871, 32'sd-0.036258920314595766, 32'sd0.0004819407298083077, 32'sd0.03213945873138667, 32'sd-0.0015664302851151472, 32'sd0.04157121886917788, 32'sd-0.003882688131845551, 32'sd0.017630813126722007, 32'sd0.04439933312998412, 32'sd0.12547581232175448, 32'sd0.12246470973758494, 32'sd0.03904621415938055, 32'sd0.06380097345909377, 32'sd-0.044483009168690926, 32'sd0.00968314036613046, 32'sd-0.05421528406396313, 32'sd0.009299270715179936, 32'sd0.07477850737058774, 32'sd0.0072738811218369245, 32'sd-0.012644251053454094, 32'sd-0.05052719984467101, 32'sd0.03790576061379027, 32'sd-0.014821123745746387, 32'sd-0.14489092386450184, 32'sd0.021626844258052464, 32'sd-0.08068690539353482, 32'sd-0.022835584445497624, 32'sd0.04898654664979376, 32'sd-0.048221028752009176, 32'sd0.03948359120530211, 32'sd0.03422681315197309, 32'sd-0.05768292858494514, 32'sd0.1114750850157035, 32'sd-0.045561444640503726, 32'sd0.028834822790388098, 32'sd-0.05052799210773685, 32'sd0.05575532214282125, 32'sd0.11103682869916258, 32'sd0.12172316545504448, 32'sd0.07980973765126566, 32'sd0.0012946909204200078, 32'sd-0.0068614545776308124, 32'sd0.015386089482611326, 32'sd0.01473658987781638, 32'sd0.06943170712974293, 32'sd0.09964923644825621, 32'sd0.05755518164449585, 32'sd0.024683917535939934, 32'sd0.01623273117686515, 32'sd-0.08553795882076268, 32'sd-0.062469848281738384, 32'sd0.0370365402571306, 32'sd-0.04330573889397944, 32'sd0.09781583917828793, 32'sd-0.039518715710401345, 32'sd-7.874177935543759e-125, 32'sd0.02008437450812766, 32'sd-0.0255678774129988, 32'sd0.0707284493803352, 32'sd-0.006774412156982895, 32'sd0.07106514989708397, 32'sd-0.012564945104637144, 32'sd0.027397020758814006, 32'sd-0.006226537253484705, 32'sd0.11345368098492895, 32'sd-0.008931817451781544, 32'sd0.0017633448086607148, 32'sd-0.021101505661524234, 32'sd0.07154104314693244, 32'sd0.11969915135635475, 32'sd0.1583593032106479, 32'sd0.0852849018011172, 32'sd0.06714115458111361, 32'sd0.17460892607781742, 32'sd0.10566534863324749, 32'sd0.013645049785288212, 32'sd-0.08282647870552665, 32'sd-0.1442771001935271, 32'sd-0.1922930397910367, 32'sd-0.049971926728097506, 32'sd-0.05234235009000447, 32'sd0.03959129762473179, 32'sd0.055191990073634685, 32'sd0.1036713878404114, 32'sd0.09596849497859235, 32'sd-0.01564965104664788, 32'sd0.034945178861997134, 32'sd0.08116635400392688, 32'sd-0.022965830460271862, 32'sd-0.07406381697350786, 32'sd-0.023659214129592463, 32'sd0.07265761625117034, 32'sd-0.024833454593045593, 32'sd0.011633852133354201, 32'sd-0.009106118324279657, 32'sd0.11547276963684651, 32'sd0.13207808185260514, 32'sd0.14603719033849186, 32'sd0.05176725760502996, 32'sd0.048101152156957074, 32'sd0.03244374572660591, 32'sd0.10133766485572021, 32'sd0.006051416572060814, 32'sd-0.08953127146104174, 32'sd-0.11970118049903308, 32'sd-0.09240709287572438, 32'sd-0.0982899856172353, 32'sd-0.08388888148120564, 32'sd0.0673642725647258, 32'sd0.011517709303602413, 32'sd0.03432107727039643, 32'sd0.10664790107344632, 32'sd0.08740579439663662, 32'sd0.04034512188487091, 32'sd-0.02069041887886098, 32'sd0.12555456963554418, 32'sd-0.039695192339143696, 32'sd-0.03637971467912504, 32'sd-0.06625593805974371, 32'sd-0.05315042050603456, 32'sd-0.007390802999217782, 32'sd0.0524485287378227, 32'sd-0.012917524902618552, 32'sd-0.07332663072792013, 32'sd-0.08646905511913205, 32'sd-0.03980013911525544, 32'sd0.18903289740661558, 32'sd-0.015013548625814117, 32'sd0.01653915419558102, 32'sd-0.10922595905477975, 32'sd-0.1088534949288226, 32'sd-0.09775696119035891, 32'sd-0.13807530950500066, 32'sd-0.17603695062572314, 32'sd-0.11574155507299452, 32'sd-0.05510693557063803, 32'sd0.02896285381313535, 32'sd0.007047549565350085, 32'sd-0.048242304156040576, 32'sd3.6039850274705273e-125, 32'sd0.04856774265842154, 32'sd0.057079873467855764, 32'sd-0.0723438374520285, 32'sd-0.035452052357043025, 32'sd-0.024348586616140946, 32'sd-0.03370010699088346, 32'sd0.015269138839754117, 32'sd-0.09178890010457634, 32'sd0.059480310457103766, 32'sd-0.034443062227499495, 32'sd-0.11481408063997738, 32'sd0.020100126404720867, 32'sd-0.003602608897571174, 32'sd0.008164004063740253, 32'sd0.08531106963452001, 32'sd0.061447526899241406, 32'sd0.007079153730645579, 32'sd-0.0328011059380885, 32'sd0.010856618593527559, 32'sd-0.008594971294024872, 32'sd-0.06969245672516719, 32'sd-0.01729716217358841, 32'sd-0.06963590752031772, 32'sd-0.04585803850204272, 32'sd-0.0298265548949731, 32'sd-0.02521036662198929, 32'sd4.922029784237379e-125, 32'sd-1.26017756494086e-118, 32'sd-7.128764596396422e-117, 32'sd0.017210681301572748, 32'sd-0.06419104274364788, 32'sd0.07950664076794822, 32'sd-0.0704709015059901, 32'sd-0.054361702123841386, 32'sd-0.08866973981425046, 32'sd0.07870531526760818, 32'sd0.021930577183613794, 32'sd-0.030786325810861433, 32'sd-0.10289997380210444, 32'sd0.059002814449322406, 32'sd-0.04579995102226349, 32'sd0.07511277373424743, 32'sd0.026217975517065173, 32'sd-0.0010388661276249165, 32'sd-0.02291127719179523, 32'sd-0.0010716629869790243, 32'sd-0.02275632590619274, 32'sd-0.104473663652808, 32'sd-0.11893020998375468, 32'sd-0.0708694365261461, 32'sd-0.0013859304123273767, 32'sd0.045350161444923966, 32'sd0.039106976625616435, 32'sd0.056844354458022155, 32'sd-7.476156556704429e-115, 32'sd-9.801791498031316e-121, 32'sd-3.2784022109018255e-119, 32'sd-0.023887330989003315, 32'sd-0.0019767419215269283, 32'sd0.030677596519953727, 32'sd-0.0713791204107965, 32'sd-0.025696246949588417, 32'sd0.04467189904463223, 32'sd-0.006754110282375107, 32'sd0.04222104870534489, 32'sd-0.05118920390382776, 32'sd-0.0068728530061712995, 32'sd-0.007978492571737925, 32'sd0.1349186326460021, 32'sd0.029023299464429154, 32'sd0.025763601417710384, 32'sd0.10718286147562477, 32'sd0.06244107092181048, 32'sd-0.0980412400919471, 32'sd-0.08276769601840009, 32'sd0.0854117045035778, 32'sd0.031846097725066226, 32'sd-0.04481793228407795, 32'sd-0.09127970945391636, 32'sd-0.047049052417017956, 32'sd0.055498889791000275, 32'sd0.018174742418754643, 32'sd1.039229238222253e-122, 32'sd5.34129169709051e-127, 32'sd3.177290353145635e-125, 32'sd3.592122446661085e-125, 32'sd0.05322579663886414, 32'sd-0.015040326089256031, 32'sd-0.011341757646307418, 32'sd-0.03176722233072796, 32'sd0.02484476147499135, 32'sd0.05880446173797711, 32'sd-0.030453827395862543, 32'sd-0.004188375349951818, 32'sd0.016424549799233492, 32'sd0.004963650965005806, 32'sd0.016593104830219422, 32'sd-0.03357960720591528, 32'sd0.03472601983781164, 32'sd0.10157129793255919, 32'sd-0.0043609839414536075, 32'sd-0.00288946072109519, 32'sd0.07454855771716362, 32'sd0.12974138133901625, 32'sd-0.004855799848662697, 32'sd-0.06564869197907436, 32'sd0.032057148323385, 32'sd0.05631319660491349, 32'sd-0.01319605936152251, 32'sd1.1237476310525099e-122, 32'sd-8.89852754048025e-126, 32'sd4.683622227494519e-118, 32'sd-1.3566808326383107e-125, 32'sd-4.8391784747833584e-122, 32'sd2.4014668879574025e-124, 32'sd0.11931582856904341, 32'sd0.00291379053139325, 32'sd0.04978692124626629, 32'sd0.08681564845329805, 32'sd-0.0126946060624361, 32'sd0.09221006206846837, 32'sd0.06172074159068016, 32'sd0.02418861768530603, 32'sd0.12196559552156933, 32'sd0.012885686581646719, 32'sd0.0805222245279683, 32'sd-0.07973400749945657, 32'sd0.020409942360629138, 32'sd0.023911546948086546, 32'sd0.04363991699407114, 32'sd0.05185273902269185, 32'sd0.04719815528834768, 32'sd0.08536831482574155, 32'sd-0.0741021826622971, 32'sd0.06703816750165072, 32'sd-1.6605681334503432e-126, 32'sd-4.598078429504248e-127, 32'sd1.9248114432654684e-122, 32'sd-1.8808901251818314e-121},
        '{32'sd1.2024271862189608e-118, 32'sd2.5635858656626357e-125, 32'sd-3.001092632268796e-126, 32'sd9.739599933096417e-123, 32'sd-3.7119166380370624e-119, 32'sd-1.4046118047712681e-118, 32'sd1.0758446826190912e-124, 32'sd-1.956927864461234e-127, 32'sd-1.037083786518362e-124, 32'sd4.6372920156504805e-118, 32'sd1.676679979733309e-125, 32'sd3.932960824159015e-124, 32'sd-0.010726276810626453, 32'sd-0.04017244415299454, 32'sd-0.025755413114465248, 32'sd-0.050590436550101564, 32'sd1.8168504089648902e-123, 32'sd3.8034182069942806e-122, 32'sd2.089790615094619e-124, 32'sd-2.1288900367335935e-127, 32'sd-7.883382814265542e-117, 32'sd2.166946221980668e-123, 32'sd-1.2439425788924615e-123, 32'sd-1.111309386786906e-121, 32'sd4.8780462528268475e-124, 32'sd7.550996107525166e-115, 32'sd-1.0912087367541485e-122, 32'sd2.270196975003319e-120, 32'sd1.1928532126459147e-118, 32'sd7.344304918376082e-123, 32'sd-7.400382000470731e-115, 32'sd-2.1637169182275484e-120, 32'sd0.005942514980607811, 32'sd-0.061500262666200414, 32'sd-0.043245037939780046, 32'sd-0.01446534714155823, 32'sd-0.06139875646832886, 32'sd-0.02939185182179157, 32'sd-0.01666521070422608, 32'sd0.04811551313880533, 32'sd0.007978661546259598, 32'sd-0.009986075950865548, 32'sd-0.05229311463416898, 32'sd-0.037054489611052115, 32'sd-0.10521583797784081, 32'sd-0.09731043273007177, 32'sd-0.0777570396365194, 32'sd-0.015637871516031982, 32'sd-0.08048686424345447, 32'sd-0.07490970778329638, 32'sd-0.05336681282350281, 32'sd-0.0137824118124733, 32'sd1.8687070686223342e-120, 32'sd2.1090580076235953e-127, 32'sd1.0552400001264685e-117, 32'sd1.9662222151084655e-119, 32'sd1.6534212545939188e-124, 32'sd2.872400062268916e-127, 32'sd-0.0411047713662934, 32'sd-0.06016031487078445, 32'sd0.07290750850156252, 32'sd0.01911053619407181, 32'sd-0.08417560747115486, 32'sd-0.00514233712426117, 32'sd0.006036091433001166, 32'sd-0.032921354093469676, 32'sd-0.005193903916427613, 32'sd-0.06560950926694017, 32'sd-0.11091824692050688, 32'sd-0.0792944086030377, 32'sd-0.09040146481813985, 32'sd-0.02165996997467454, 32'sd-0.01910531749368293, 32'sd-0.026471323278712492, 32'sd0.07499112829188344, 32'sd0.012958877852638166, 32'sd0.013834589196473809, 32'sd-0.050020133335537745, 32'sd-0.007632240912372328, 32'sd0.06495161682041456, 32'sd0.015797145611758382, 32'sd-0.04573252706570771, 32'sd1.1081527392373829e-126, 32'sd3.0701985009810268e-118, 32'sd-1.710205312294629e-125, 32'sd1.5748172768987753e-114, 32'sd-0.01849412103633957, 32'sd-0.06291093278016964, 32'sd0.026610831879319438, 32'sd0.03842996410436601, 32'sd-0.11068152040323377, 32'sd-0.08466572966858628, 32'sd-0.055405465949360695, 32'sd-0.01754217990412056, 32'sd-0.051337273494256354, 32'sd-0.09637996561186361, 32'sd-0.15568666314161975, 32'sd-0.1781616664296086, 32'sd-0.12168877592114102, 32'sd0.03070945722965946, 32'sd-0.0398095243150128, 32'sd-0.034078558250770705, 32'sd0.08732380027905014, 32'sd0.06353363418790232, 32'sd-0.024670286324723463, 32'sd0.0700291476170753, 32'sd0.07172695274486933, 32'sd-0.0627298515247909, 32'sd0.041592158547182484, 32'sd0.05955462888263786, 32'sd-0.010609343562186867, 32'sd2.1174414469258763e-117, 32'sd3.724252156123612e-129, 32'sd-0.03975984047928522, 32'sd0.020037602521158555, 32'sd-0.1428870309627374, 32'sd-0.026096452931776985, 32'sd-0.08016888077832182, 32'sd-0.005662686743609821, 32'sd-0.1152772485989604, 32'sd-0.06368477439059286, 32'sd-0.062034616791641205, 32'sd-0.05433490704184444, 32'sd-0.02729337473060009, 32'sd0.03436000763805148, 32'sd-0.09823736416093704, 32'sd-0.009882201445721196, 32'sd-0.02220199951002737, 32'sd0.09177750669464718, 32'sd0.05871069777813149, 32'sd0.03148777268301204, 32'sd-0.13000287431619706, 32'sd-0.08135887204665196, 32'sd0.002249384599343323, 32'sd0.0061183347565290855, 32'sd-0.030805985513230338, 32'sd0.07491202694849516, 32'sd0.029921547659522995, 32'sd0.06588930647345578, 32'sd-0.08734110451323257, 32'sd-2.142366588946486e-122, 32'sd0.005893113811973709, 32'sd-0.045363728499735856, 32'sd-0.04779313799082633, 32'sd-0.01868536081427627, 32'sd-0.03284612643935013, 32'sd-0.04591317314599578, 32'sd-0.09482734180421788, 32'sd-0.02084467733319828, 32'sd-0.06968388208460231, 32'sd-0.014579886592433262, 32'sd0.029557286887819053, 32'sd0.08762670069980055, 32'sd0.06538769682099986, 32'sd0.0963229682775849, 32'sd0.008025407122955965, 32'sd0.0538737667695397, 32'sd0.0064275680914839955, 32'sd-0.038185902392147086, 32'sd-0.10753613163487444, 32'sd-0.0818107322961941, 32'sd0.03412756580634495, 32'sd0.04523566580332717, 32'sd-0.08873766120139222, 32'sd-0.10162375691069221, 32'sd-0.0063613391034786386, 32'sd0.01604370159792837, 32'sd0.04668384084128069, 32'sd-1.4301481620743972e-122, 32'sd0.038272928341326125, 32'sd-0.08734087857805042, 32'sd0.051780346498302265, 32'sd-0.12078835289690089, 32'sd0.10333674595911832, 32'sd0.01661051381684402, 32'sd-0.07290721002183001, 32'sd-0.07242543015409612, 32'sd0.01894515110894892, 32'sd0.12486538930182225, 32'sd0.03650592247046482, 32'sd-0.03785285498789651, 32'sd-0.13694959131381193, 32'sd0.001084080827469148, 32'sd-0.1936296142412472, 32'sd-0.15161516314544377, 32'sd-0.184471918762144, 32'sd-0.006316871987904942, 32'sd-0.03301046735709057, 32'sd-0.012027386199884296, 32'sd-0.08976763565823503, 32'sd-0.04514743079538077, 32'sd0.07713278377856649, 32'sd-0.02184322699545087, 32'sd-0.024482805065707842, 32'sd-0.04701652521636627, 32'sd0.03618749520745177, 32'sd-0.052744228515861906, 32'sd0.06030709247268632, 32'sd-0.011922789597792784, 32'sd-0.07116367379813765, 32'sd-0.1259422673003795, 32'sd-0.0345010521476623, 32'sd-0.06289338430360529, 32'sd-0.09932034239558724, 32'sd0.011597886580965557, 32'sd0.02769510259807245, 32'sd0.09260479883174064, 32'sd-0.10833975552979869, 32'sd-0.13256572642002246, 32'sd-0.02942335486505301, 32'sd-0.15820102353277604, 32'sd-0.020120151752215393, 32'sd0.0014836043818308787, 32'sd-0.047826789418988276, 32'sd0.044135413205199814, 32'sd0.1311343119900567, 32'sd0.09270229571471658, 32'sd0.03305409515441685, 32'sd0.15755610988545862, 32'sd0.002366808410755327, 32'sd-0.01234481772240211, 32'sd0.024147067879981186, 32'sd0.0639609777531174, 32'sd-0.04089911949339387, 32'sd-0.022287080293051455, 32'sd0.015642545180244383, 32'sd0.039188753127787114, 32'sd-0.08060983715331484, 32'sd-0.07356155190077043, 32'sd-0.08615062474349137, 32'sd-0.015851615217188537, 32'sd0.030768563654589763, 32'sd0.14177671202416722, 32'sd0.009674049603459306, 32'sd-0.02872978846752045, 32'sd-0.07829281740554855, 32'sd-0.06180780139312209, 32'sd-0.05952151723549306, 32'sd0.12806498353457582, 32'sd0.057296657757477804, 32'sd0.0907789682853353, 32'sd0.07050838467757306, 32'sd0.06759863324492357, 32'sd0.03926425186042234, 32'sd0.15827428163447055, 32'sd0.1260602680095087, 32'sd0.05816411382273289, 32'sd0.022968795526415682, 32'sd0.05840303368624948, 32'sd-0.0979623700131387, 32'sd0.022899997468636586, 32'sd-0.08706327006427773, 32'sd-0.0609252397237765, 32'sd-0.003843847769191841, 32'sd-0.053453566584763385, 32'sd-0.09326839285171282, 32'sd-0.01521539644349153, 32'sd0.056362559319208194, 32'sd-0.03162764802378303, 32'sd0.043366092212256034, 32'sd0.0778974621718612, 32'sd0.051450631503298955, 32'sd-0.025659985359404936, 32'sd-0.05075764976121426, 32'sd0.04548104889784929, 32'sd0.07455896534233014, 32'sd0.03915033876520932, 32'sd0.13419667931914286, 32'sd0.1465349267461278, 32'sd0.017721361176204483, 32'sd0.013298294659104986, 32'sd0.05590246479748162, 32'sd-0.039639865656585026, 32'sd0.023609022366884554, 32'sd0.09845230784294001, 32'sd0.09002013015476519, 32'sd-0.0641183694476853, 32'sd-0.01740891116336049, 32'sd-0.025396952701422816, 32'sd-0.07813878927407798, 32'sd-0.05778909169588948, 32'sd-0.08041875142683251, 32'sd-0.08749054960869743, 32'sd-0.1356004417049009, 32'sd-0.006991889597176574, 32'sd0.018432635182582098, 32'sd-0.011628760908085683, 32'sd0.07207009942711139, 32'sd0.10619167123670224, 32'sd-0.016975578200968275, 32'sd0.030837624327551345, 32'sd-0.15998002909751388, 32'sd0.01686881313997137, 32'sd-0.10967332846918997, 32'sd-0.053593212913806344, 32'sd-0.017622019490721105, 32'sd-0.02717079512072764, 32'sd0.044911427648717785, 32'sd-0.023269598841358784, 32'sd0.020260989593132276, 32'sd-0.027509387617516267, 32'sd-0.05643302670010484, 32'sd0.10704020955717708, 32'sd0.019450575834603908, 32'sd0.06309422678033372, 32'sd0.11900881579642758, 32'sd0.004517254673717422, 32'sd0.06219503298094042, 32'sd-0.009895905564470661, 32'sd-0.007853239735251122, 32'sd-0.08290102877238385, 32'sd-0.1287630828910769, 32'sd-0.009031878069009057, 32'sd0.0715473334013071, 32'sd0.061524747592812956, 32'sd0.04440006895268442, 32'sd-0.03180247803862212, 32'sd0.22667933210218397, 32'sd0.18293790652352906, 32'sd-0.008835669322266522, 32'sd-0.07128142154416206, 32'sd-0.19437983866044228, 32'sd-0.17256645284651453, 32'sd-0.141179995312093, 32'sd-0.0012001890025773465, 32'sd0.0119907326943659, 32'sd-0.07679957259006419, 32'sd0.0035343673098376287, 32'sd-0.08786705669054197, 32'sd0.044148404983803284, 32'sd0.1308910088400602, 32'sd0.044735715636653225, 32'sd0.05121352746465537, 32'sd0.034755980184191446, 32'sd0.1748270445293527, 32'sd-0.033919532603458584, 32'sd0.027641492245997844, 32'sd0.04574837254128457, 32'sd-0.04269042279765971, 32'sd-0.0009360629285084362, 32'sd0.023465960835241467, 32'sd0.07647922268897804, 32'sd-0.021123947033971115, 32'sd0.10045017205819362, 32'sd0.21858773853646585, 32'sd0.3075315193346847, 32'sd0.20502741258752546, 32'sd0.14363512601979359, 32'sd-0.007928420704712572, 32'sd-0.06295147566311829, 32'sd-0.18666039842126914, 32'sd-0.1369956991676456, 32'sd-0.05286091192235094, 32'sd0.11632220185670997, 32'sd-0.04303952691158524, 32'sd0.007493136805486423, 32'sd-0.03129973972448689, 32'sd-0.01749858577006672, 32'sd0.051771586248381386, 32'sd0.17342586272256308, 32'sd0.06310622939903407, 32'sd0.043985186871810474, 32'sd0.10372156017414767, 32'sd0.051175371519917676, 32'sd-0.035760815628613524, 32'sd0.1192957716313632, 32'sd0.0632574233085588, 32'sd-0.11106292190441064, 32'sd-0.06261280768274785, 32'sd-0.1203988679538159, 32'sd-0.16735937804698903, 32'sd-0.04959577177255723, 32'sd0.05549990242180009, 32'sd0.2818732315265449, 32'sd0.1954418641483704, 32'sd0.18481903908201974, 32'sd0.12092051723840988, 32'sd0.20991785492102571, 32'sd0.08043414411972842, 32'sd0.024608342015483203, 32'sd0.07576229228449682, 32'sd-0.014969820212164408, 32'sd0.0076727225604474635, 32'sd-0.007798213261503131, 32'sd0.010016263239600542, 32'sd0.01707067017850066, 32'sd0.08369676502394784, 32'sd0.04732181330477087, 32'sd-0.07397134234247502, 32'sd0.06650803025738261, 32'sd0.03865899277865557, 32'sd0.03010703782037433, 32'sd-0.02171946208819889, 32'sd0.0568375014228201, 32'sd-0.05278216317143921, 32'sd-0.0007565259339997873, 32'sd-0.04790609715274307, 32'sd-0.02617653215608516, 32'sd-0.1561174459196492, 32'sd-0.13235960029657426, 32'sd-0.013206523497892635, 32'sd0.01431412330540497, 32'sd0.17873649401680203, 32'sd0.15461272682176652, 32'sd0.21615652092832555, 32'sd0.20129408474554367, 32'sd0.1042704467079225, 32'sd-0.13225813402722897, 32'sd-0.12310138021008799, 32'sd0.06322663572237651, 32'sd-0.09709518102799014, 32'sd-0.005251317683891432, 32'sd-0.005658673645668569, 32'sd0.033207407936956854, 32'sd-0.01053849290773915, 32'sd-0.04642405987458317, 32'sd-0.07697887540720288, 32'sd0.06850094612851185, 32'sd0.03152749299261275, 32'sd-0.055695018755046725, 32'sd0.08463772145041291, 32'sd-0.01682794021239947, 32'sd-0.08772661459196761, 32'sd0.061518330863158, 32'sd-0.07045404061748538, 32'sd-0.08530074922118182, 32'sd-0.22567123598276603, 32'sd-0.2768455377605991, 32'sd-0.21131408880243308, 32'sd-0.06201016914211979, 32'sd0.13120074837941795, 32'sd0.10792657650225643, 32'sd0.05864192602808004, 32'sd0.09272645666214153, 32'sd0.11889214236977935, 32'sd0.02047086138483574, 32'sd-0.012556132317902749, 32'sd-0.027262058059173373, 32'sd-0.023751380797031846, 32'sd-0.026763565692273363, 32'sd-0.07022480043552107, 32'sd-0.04998627261159785, 32'sd-0.19973419689936392, 32'sd-0.007353734719202257, 32'sd-0.22534364608348187, 32'sd-0.12078471058887477, 32'sd-0.16484325939359595, 32'sd-0.023514084255966343, 32'sd0.004966869447224065, 32'sd-0.08491695257018932, 32'sd-0.1492836699172751, 32'sd0.16358414292269338, 32'sd0.012178237527597186, 32'sd-0.15021520812126798, 32'sd-0.32825456022666466, 32'sd-0.26849916780265104, 32'sd-0.2741693040645489, 32'sd-0.13781812947043573, 32'sd-0.1575154967335126, 32'sd-0.19957018177579577, 32'sd-0.06716894598840235, 32'sd0.053617433417350466, 32'sd0.013362484998837626, 32'sd0.05411598887883462, 32'sd-0.05872166780911507, 32'sd-0.02351722434392285, 32'sd-0.11191548762828366, 32'sd-0.1507506424150598, 32'sd-0.18906673745505276, 32'sd-0.19289357323995177, 32'sd-0.09059825467091309, 32'sd-0.0745251067602474, 32'sd-0.20985016977007534, 32'sd-0.15364801660933786, 32'sd0.0235237056544169, 32'sd-0.0336516987605325, 32'sd-1.4475438073650263e-123, 32'sd0.038345645272450844, 32'sd-0.06964154263196257, 32'sd-0.008870976431394872, 32'sd0.07322430188826444, 32'sd-0.01670904345395626, 32'sd-0.09651202480482092, 32'sd-0.18049336527416823, 32'sd-0.3470673057402347, 32'sd-0.15693847682816292, 32'sd-0.3007027298355872, 32'sd-0.2130958305101632, 32'sd-0.12535615888811386, 32'sd0.08942347759206173, 32'sd-0.019830649432911688, 32'sd-0.06155354394389237, 32'sd-0.09676273016481958, 32'sd-0.04867587970023265, 32'sd0.009461434824650719, 32'sd-0.12584110289692024, 32'sd-0.05904804842907514, 32'sd-0.1689176609330484, 32'sd-0.13724677196580432, 32'sd-0.07931004307258784, 32'sd-0.1651805602424535, 32'sd0.029947970991240268, 32'sd0.05424960931491029, 32'sd0.0009337455404784568, 32'sd0.0007394173217453507, 32'sd0.050279609503098135, 32'sd0.007074898715219726, 32'sd-0.0004382879233318144, 32'sd0.11315957689719407, 32'sd0.1212525580265256, 32'sd-0.03253627819069515, 32'sd-0.08175666737655585, 32'sd-0.0512227880632284, 32'sd-0.17759092054742076, 32'sd-0.09206787090375264, 32'sd-0.08007546591600206, 32'sd-0.07821691542933933, 32'sd0.05282052937445287, 32'sd0.017461091204133555, 32'sd0.04776968284026189, 32'sd-0.07161622667146691, 32'sd-0.005241759131200777, 32'sd-0.0834300928146857, 32'sd-0.03625232429444446, 32'sd0.015750283999801305, 32'sd-0.048161113574725016, 32'sd-0.06895661198467003, 32'sd-0.0699322552067424, 32'sd-0.121540609165073, 32'sd0.05226406713199836, 32'sd0.05516877443755625, 32'sd-0.023115774099494286, 32'sd-0.039226684125877286, 32'sd-0.023206946762080603, 32'sd0.005398655865944257, 32'sd-0.0717313238789228, 32'sd-0.05079931436312626, 32'sd0.021229921626580158, 32'sd-0.050254448798567226, 32'sd0.07379710218719546, 32'sd0.1716870474117493, 32'sd-0.014644615774408249, 32'sd0.04853494040046639, 32'sd-0.16402679794751288, 32'sd-0.020764660833780597, 32'sd0.09179654627043389, 32'sd0.12184193883892079, 32'sd0.0396421210825696, 32'sd-0.011363479020416208, 32'sd-0.11076439126587652, 32'sd0.040219494112858016, 32'sd0.0077531852497499595, 32'sd0.06896951198033018, 32'sd-0.12357637060471965, 32'sd-0.011809396407667806, 32'sd-0.15882065757721595, 32'sd-0.051738945980246365, 32'sd0.02858927172094349, 32'sd-0.06919978754249334, 32'sd0.007765981743577993, 32'sd-1.3277709090278815e-118, 32'sd-0.005963105344787912, 32'sd0.0034223466142056284, 32'sd0.04502549890407938, 32'sd-0.11716391785318221, 32'sd-0.06631073650853386, 32'sd-0.04486613825056296, 32'sd0.1043138257537273, 32'sd0.07416169938604372, 32'sd0.11450268824046746, 32'sd0.019764730891348784, 32'sd-0.016250113825394652, 32'sd-0.049625006170924614, 32'sd0.05818542388507789, 32'sd-0.09063909644338393, 32'sd-0.014740133149441444, 32'sd-0.07913921680143789, 32'sd-0.03153859894153511, 32'sd0.0062587363338178085, 32'sd-0.01877619048242131, 32'sd0.02222484461130957, 32'sd-0.11622104949781191, 32'sd-0.03410319535111664, 32'sd-0.10038716796676513, 32'sd-0.06604851911474444, 32'sd-0.02762637615324933, 32'sd0.007418726073654017, 32'sd-0.0128384569195922, 32'sd-0.054068981467734936, 32'sd-0.08609175648538486, 32'sd-0.06763265406543245, 32'sd-0.11169271992250414, 32'sd-0.02113907324395849, 32'sd-0.003975611015102313, 32'sd-0.014914542346582576, 32'sd0.03597721102225168, 32'sd0.07054740125643102, 32'sd0.15972761559809656, 32'sd0.07317506295707131, 32'sd0.09974272172424534, 32'sd-0.009960619729291673, 32'sd0.03429314350039989, 32'sd-0.07049848526226803, 32'sd0.022763596960915386, 32'sd-0.028974560635426486, 32'sd0.060357204770668055, 32'sd0.10035948586554433, 32'sd-0.1253810583817266, 32'sd-0.024629166405236363, 32'sd-0.08429947557025974, 32'sd0.053447480770418485, 32'sd-0.08557573837845499, 32'sd-0.11971281843745732, 32'sd-0.06374550890312325, 32'sd-0.05548350491348612, 32'sd0.010714662880398938, 32'sd-0.030008419105359625, 32'sd0.017946307953835925, 32'sd-0.02048069694201388, 32'sd-0.052489520152193124, 32'sd-0.011379729101345453, 32'sd-0.10131933985873377, 32'sd-0.02261985566336023, 32'sd0.12064120894414927, 32'sd0.08583995431320927, 32'sd0.045202777602767225, 32'sd0.02773553807094775, 32'sd0.015963476086400072, 32'sd0.009638553847280134, 32'sd0.05413730939448451, 32'sd0.17297313967323139, 32'sd0.11666050168956399, 32'sd-0.004400051484346783, 32'sd0.13012719849811483, 32'sd-0.03478826617762021, 32'sd-0.052557311438152066, 32'sd-0.13709928465591512, 32'sd-0.07593409424723163, 32'sd-0.06485848386484483, 32'sd0.040664877151631154, 32'sd-0.04106683187714878, 32'sd-0.03394325598140771, 32'sd-0.016401158484649365, 32'sd-0.04474303421197765, 32'sd8.771943294126e-127, 32'sd-0.04683932552630277, 32'sd-0.02656257534373392, 32'sd-0.060271160980033656, 32'sd-0.03557995088367376, 32'sd0.07110842233473375, 32'sd-0.049311108787966525, 32'sd0.04648396346479112, 32'sd0.029661646931567552, 32'sd0.0044300131724828275, 32'sd-0.050556547590938944, 32'sd0.08926075055426289, 32'sd0.06940662817264968, 32'sd0.047182230191630946, 32'sd-0.007938586559648178, 32'sd0.07460667304789524, 32'sd0.005949977500705546, 32'sd0.1016548781601031, 32'sd-0.056924547896063674, 32'sd-0.06559462995820127, 32'sd0.0663176782650839, 32'sd-0.09139568500393419, 32'sd-0.0971288637388826, 32'sd0.07576313287530466, 32'sd0.028695340028892246, 32'sd-0.14926824329646177, 32'sd-0.07718599484178593, 32'sd1.0740339398877353e-124, 32'sd-1.2253985679038562e-124, 32'sd8.98506810652544e-124, 32'sd-0.0010706086139471518, 32'sd0.011747242499433461, 32'sd-0.05727714144435894, 32'sd-0.007328451310680922, 32'sd-0.05689827680817447, 32'sd0.011568626259090201, 32'sd-0.07449439859570638, 32'sd-0.18646812741997373, 32'sd-0.026764703428282296, 32'sd0.040111915206351045, 32'sd-0.05769578947187139, 32'sd0.07491192918179276, 32'sd0.005649920583940445, 32'sd0.035818480197730616, 32'sd-0.01776803573861819, 32'sd-0.07885433427311479, 32'sd0.12074712439949432, 32'sd0.13486035731594048, 32'sd0.005266932413707409, 32'sd-0.04753728292690804, 32'sd-0.10151173030131208, 32'sd0.07758890838567069, 32'sd-0.03552681974034954, 32'sd-0.06717692768206916, 32'sd-0.05816671333480321, 32'sd9.80141089975917e-121, 32'sd4.654703501749885e-124, 32'sd2.1691255264214623e-119, 32'sd-0.03145548242111715, 32'sd-0.01664724313205247, 32'sd-0.03103477081553522, 32'sd0.049237070094795644, 32'sd0.006739496270952938, 32'sd-0.04814024080652392, 32'sd-0.002043356988475783, 32'sd-0.08344631532023541, 32'sd-0.027831033859407325, 32'sd-0.022266500187410648, 32'sd-0.027501452789212663, 32'sd0.0554145001979538, 32'sd0.05370320882734871, 32'sd0.010752921392644919, 32'sd0.025608652615821074, 32'sd0.0698650479432235, 32'sd0.030329022493818147, 32'sd0.0953824322170912, 32'sd0.03527847042556826, 32'sd-0.024868795374781913, 32'sd0.021020188823614814, 32'sd-0.004365361007892017, 32'sd-0.048680844670430504, 32'sd0.010295529318017993, 32'sd-0.008088523878274044, 32'sd-1.5459714149579153e-115, 32'sd-8.214795405812229e-117, 32'sd2.1976374504653694e-121, 32'sd-7.287807214845328e-117, 32'sd-0.054207041319272044, 32'sd0.04446748980190533, 32'sd0.004745545717447567, 32'sd0.12192047478188288, 32'sd-0.0399777326442216, 32'sd0.14782088483227154, 32'sd-0.008096723565931873, 32'sd-0.006958381908788568, 32'sd-0.0034786754795052, 32'sd0.08716103238348025, 32'sd-0.0628826346870157, 32'sd0.13077118159332746, 32'sd0.11483112190824488, 32'sd0.07887851529936309, 32'sd0.047326015233075426, 32'sd0.07131043568340628, 32'sd-0.02349977080583824, 32'sd-0.07555149747260897, 32'sd0.028156358716476194, 32'sd-0.00610346072120717, 32'sd0.03697950971831654, 32'sd0.04743770759273323, 32'sd-0.04230026570438554, 32'sd3.6095450305577906e-123, 32'sd6.202897870782943e-121, 32'sd1.6489118310668164e-117, 32'sd-1.3653826847565915e-127, 32'sd5.2468674625105025e-127, 32'sd1.811272940078401e-123, 32'sd-0.0465728541677913, 32'sd-0.014398775960029815, 32'sd-0.10019297569447387, 32'sd0.061341747363059, 32'sd-0.02403059410900699, 32'sd0.01877960238871389, 32'sd0.03730859689140567, 32'sd-0.013580490656545686, 32'sd0.05970666294789586, 32'sd0.05947576929173156, 32'sd-0.04784226679525809, 32'sd0.033743557107153266, 32'sd0.005383353972521746, 32'sd0.01939641330588331, 32'sd0.0312956936298288, 32'sd0.02996469244178269, 32'sd0.0328453038401803, 32'sd-0.011975048227310324, 32'sd-0.03622632217689142, 32'sd-0.015827331882106513, 32'sd-1.4755543288331494e-123, 32'sd1.0903588055193332e-117, 32'sd2.066839044361438e-121, 32'sd-2.612429062769762e-126},
        '{32'sd-4.664073029053191e-127, 32'sd5.260194921617317e-115, 32'sd-1.729699634665817e-125, 32'sd3.1829303510497043e-121, 32'sd-1.4136296807130703e-120, 32'sd-1.8980233959647304e-115, 32'sd-8.882344547914429e-127, 32'sd-1.0768132092775554e-124, 32'sd-5.847006256282128e-119, 32'sd2.0197787220333276e-121, 32'sd-9.529315368693283e-115, 32'sd1.04939093996423e-120, 32'sd-0.057072125285707105, 32'sd-0.008041259576734591, 32'sd-0.035034067002471685, 32'sd-0.07166707887704486, 32'sd3.06385698933612e-120, 32'sd-1.3185186091208987e-127, 32'sd-1.4362797263424183e-118, 32'sd6.887448141601451e-124, 32'sd-4.698290110058851e-122, 32'sd9.174253629180257e-115, 32'sd7.842105218963489e-117, 32'sd1.0916959770003496e-119, 32'sd-5.929385934238716e-117, 32'sd-2.944821577282262e-129, 32'sd2.712103491964215e-124, 32'sd4.830994668504382e-124, 32'sd3.87392403457294e-123, 32'sd-2.8288182778654944e-121, 32'sd2.3945279159386954e-119, 32'sd-2.107988777125543e-117, 32'sd-0.08164887958329503, 32'sd-0.05517765363865604, 32'sd-0.05885764998711414, 32'sd-0.08346080581863793, 32'sd-0.09498310490778462, 32'sd-0.13010665416299838, 32'sd-0.06734176782629751, 32'sd0.017477904990854814, 32'sd-0.06850553868448786, 32'sd-0.036681463056240905, 32'sd-0.07919567533002107, 32'sd-0.10902604567254853, 32'sd-0.05173462110831301, 32'sd-0.11552338211197297, 32'sd-0.12185668774474501, 32'sd-0.11810398149919661, 32'sd-0.08404618095320628, 32'sd-0.04267194783316555, 32'sd0.01274063373561711, 32'sd0.0386903496056025, 32'sd8.774458726011938e-122, 32'sd3.1963923118072787e-127, 32'sd-4.102180215775352e-121, 32'sd8.594347549307736e-117, 32'sd-1.5052501019228714e-128, 32'sd-6.55306455623018e-117, 32'sd-0.07268348135798777, 32'sd-0.05792353557134223, 32'sd-0.09137984128561594, 32'sd0.05458854972485842, 32'sd0.09861980577959911, 32'sd-0.015326082237984266, 32'sd0.049522717024283354, 32'sd-0.10609749984274017, 32'sd-0.015672191637537507, 32'sd-0.051992767850543915, 32'sd-0.03657145721350835, 32'sd-0.08243638083926072, 32'sd-0.03372536034901685, 32'sd-0.04367633691447883, 32'sd-0.050838935779709486, 32'sd-0.09546161883442916, 32'sd-0.06477048834691025, 32'sd-0.10852328977287092, 32'sd-0.1310562619123554, 32'sd-0.12481351147677595, 32'sd-0.04263364643482031, 32'sd0.03224923037914305, 32'sd-0.023364558553281893, 32'sd-0.10626819400785657, 32'sd-3.323207015978805e-126, 32'sd-3.0973224133607595e-118, 32'sd6.770824984049458e-127, 32'sd-2.012168518280704e-119, 32'sd-0.09127565252952952, 32'sd-0.02346874919809765, 32'sd-0.08265127375726881, 32'sd-0.05887821115066422, 32'sd-0.03249303548471817, 32'sd0.10592558362804083, 32'sd0.008048643408678651, 32'sd-0.07357035296162316, 32'sd-0.0045922339314661215, 32'sd-0.05695590151465319, 32'sd-0.03717200129651047, 32'sd0.08102519656129906, 32'sd0.20141219750063652, 32'sd-0.0158314815735828, 32'sd0.006283369376856592, 32'sd-0.028550267150644803, 32'sd-0.048961930896706245, 32'sd-0.2472914167644662, 32'sd-0.13317171895617386, 32'sd-0.0029670925802385215, 32'sd0.03782516574206776, 32'sd0.05238793396403861, 32'sd-0.04291470843243117, 32'sd-0.058156731331657024, 32'sd-0.08739638825829063, 32'sd-1.3810261743326643e-117, 32'sd1.8554663227031366e-116, 32'sd0.02021573263480427, 32'sd-0.013454061823252402, 32'sd-0.026301764627895147, 32'sd0.11189590313752945, 32'sd0.0853599015996227, 32'sd0.09951828015892095, 32'sd0.009716674204389002, 32'sd0.024829263973554897, 32'sd-0.07328145619760569, 32'sd-0.004101636868285649, 32'sd-0.03661716459517292, 32'sd0.13166122204177255, 32'sd0.1828418378820861, 32'sd0.006637730029658227, 32'sd0.029494341552315482, 32'sd-0.045081625957699385, 32'sd0.07527801927199876, 32'sd-0.07846033869924397, 32'sd-0.10398857305310213, 32'sd-0.17781958112871113, 32'sd-0.14098537986570125, 32'sd0.053673580463385356, 32'sd-0.0746823325650488, 32'sd0.014979199684190588, 32'sd-0.01637559443886147, 32'sd-0.04415430352604335, 32'sd-0.043389478789926175, 32'sd-3.6986716479552893e-128, 32'sd-0.06576753414685252, 32'sd0.027289322025712624, 32'sd-0.11173991202353267, 32'sd-0.028006439760509424, 32'sd0.023278199966421186, 32'sd-0.051126173384969525, 32'sd-0.13234063872793972, 32'sd-0.13341022600572358, 32'sd-0.11456427904484108, 32'sd-0.06557850392243675, 32'sd0.011592206747101185, 32'sd0.08181529424059482, 32'sd0.012793261268454797, 32'sd0.06049843689562683, 32'sd0.21444890389160065, 32'sd0.2225186380003028, 32'sd0.014516672404712579, 32'sd0.08020230355978991, 32'sd0.14901938177956783, 32'sd-0.12196212338730365, 32'sd-0.09635103829128829, 32'sd-0.04844195094912971, 32'sd0.0535336726688189, 32'sd0.022478754955908096, 32'sd0.04107519977328002, 32'sd0.05342928404708627, 32'sd-0.0974717440334194, 32'sd-1.3838579929994695e-125, 32'sd0.052380142648726175, 32'sd0.010554268609252654, 32'sd-0.06575514614801954, 32'sd-0.043722579914228024, 32'sd-0.03409931826871998, 32'sd-0.05603369884963577, 32'sd-0.129632027663737, 32'sd-0.036707229425344004, 32'sd0.06654908921115314, 32'sd0.05438704123565271, 32'sd0.0518425448274049, 32'sd0.11110275329304053, 32'sd0.12432050093181533, 32'sd0.18475013271514873, 32'sd0.16801596470315827, 32'sd0.08554700660170726, 32'sd0.13757085206767738, 32'sd0.07131973845810972, 32'sd-0.06017631357118597, 32'sd-0.05545145616579816, 32'sd-0.05761969656199315, 32'sd0.09616880007818855, 32'sd0.02110664853866833, 32'sd0.06228175553683016, 32'sd-0.05824278404948259, 32'sd0.06656071964763204, 32'sd0.03624802233549093, 32'sd-0.025700656934936995, 32'sd-0.051570643664360004, 32'sd-0.06765550628320945, 32'sd-0.0004958670933625496, 32'sd-0.11815229464238206, 32'sd0.05594842133181035, 32'sd-0.01518402837548293, 32'sd0.01526081580604246, 32'sd-0.0800388628289983, 32'sd0.06178332761859092, 32'sd0.11762047898122513, 32'sd0.0664438804595347, 32'sd0.12618302547026825, 32'sd-0.003616366248134377, 32'sd-0.04836912132794809, 32'sd-0.0735232664297142, 32'sd-0.030851707367458972, 32'sd0.02371917867621073, 32'sd-0.059774345153851806, 32'sd-0.04876271934437402, 32'sd-0.1069721677690082, 32'sd-0.16559474992272782, 32'sd0.003055550094683033, 32'sd0.009615209475249634, 32'sd0.04242045162640964, 32'sd-0.10978306087250464, 32'sd-0.053531296706656586, 32'sd-0.0419265739295542, 32'sd-0.09289416899228083, 32'sd-0.07153212258602847, 32'sd0.04164561213938393, 32'sd0.06114312112821136, 32'sd0.028769672403550762, 32'sd0.013362272782037752, 32'sd0.04963516203405486, 32'sd0.029418435781886763, 32'sd0.14422676869652074, 32'sd0.17698033391280496, 32'sd0.013765193179389585, 32'sd0.02694364300549379, 32'sd-0.020068687437974447, 32'sd-0.20791832300229962, 32'sd-0.1321620363149425, 32'sd-0.06169077264580975, 32'sd0.02332854275602329, 32'sd0.0942871375636086, 32'sd0.20977199572764763, 32'sd0.08672587634716683, 32'sd-0.03488669252934384, 32'sd-0.044939787463623294, 32'sd-0.0081209117077326, 32'sd0.014449631161524255, 32'sd-0.03990268284030244, 32'sd0.025778983918588582, 32'sd-0.01820014856224502, 32'sd0.008908181678282275, 32'sd-0.02799204419485772, 32'sd-0.13213342723650717, 32'sd-0.019476241648409613, 32'sd-0.029256269242485575, 32'sd0.02699846133633227, 32'sd-0.002293828706244392, 32'sd0.07653796049584727, 32'sd0.10953819685269307, 32'sd0.16636662588784681, 32'sd0.07443961536679992, 32'sd0.05669176295276367, 32'sd-0.03645595680740777, 32'sd-0.2032017769363784, 32'sd-0.15173677660311113, 32'sd-0.23001454682361333, 32'sd0.0542187288310777, 32'sd0.16336667833578908, 32'sd0.3417398543520479, 32'sd0.186396193757407, 32'sd0.19450447689600392, 32'sd0.061512467431685286, 32'sd0.0370218260707685, 32'sd-0.012134225306943596, 32'sd-0.06180445580210505, 32'sd-0.198845983256508, 32'sd-0.05391841069267904, 32'sd0.025874597963769275, 32'sd0.0629396555276281, 32'sd-0.06086311416919957, 32'sd-0.0263928487932905, 32'sd-0.05602924270824109, 32'sd0.06738946464805524, 32'sd-0.02920571839981131, 32'sd0.08279697942445637, 32'sd-0.03054310150949548, 32'sd0.039697649846450495, 32'sd-0.0020471027856006994, 32'sd0.05007422306962767, 32'sd-0.13944689232738325, 32'sd-0.11421609565790031, 32'sd-0.29785011620025986, 32'sd-0.23750382969806907, 32'sd-0.1119236530651973, 32'sd0.009824235279389843, 32'sd0.17452041977427013, 32'sd0.20383614330804764, 32'sd0.10226921137910679, 32'sd0.20321152557066866, 32'sd0.11919187852655547, 32'sd0.05293862138173949, 32'sd0.06717556532659183, 32'sd-0.09836707821650269, 32'sd-0.1749144776885377, 32'sd0.04327946799459845, 32'sd-0.013955056615945056, 32'sd0.0636139068680826, 32'sd-0.061512896157288985, 32'sd-0.12516359639541186, 32'sd-0.0013410131371386388, 32'sd-0.06614235069838127, 32'sd-0.012096173027170325, 32'sd0.06997255548809797, 32'sd-0.04362984841954173, 32'sd-0.013250182026528815, 32'sd0.05375037226859437, 32'sd-0.010544436211023382, 32'sd-0.03340693037494906, 32'sd-0.24356772274146968, 32'sd-0.1993258311062432, 32'sd-0.103747483451958, 32'sd0.07155707384991679, 32'sd0.11409381844295105, 32'sd0.1279353024942931, 32'sd0.15113414679528017, 32'sd0.15618319773763098, 32'sd0.22085755688313452, 32'sd0.14811259004575372, 32'sd-0.009881643904521143, 32'sd0.05380772050652741, 32'sd0.03149034456749971, 32'sd-0.17191475341047796, 32'sd-0.1002752299393096, 32'sd-0.06970309627363512, 32'sd-0.10262563998983977, 32'sd-0.06648484609932975, 32'sd-0.03416364306170272, 32'sd0.0485206653481631, 32'sd-0.058289259904094934, 32'sd0.04383082533093676, 32'sd0.03980809235531378, 32'sd-0.11022942682588363, 32'sd0.017100786307030283, 32'sd-0.01692499814514293, 32'sd-0.02884987642654205, 32'sd-0.05427346447627876, 32'sd-0.07589093116144405, 32'sd-0.023096352063172586, 32'sd0.0159937518677541, 32'sd0.03701586605582643, 32'sd0.04668397746430908, 32'sd-0.005192735041181461, 32'sd-0.06316856055748778, 32'sd0.11933574307628074, 32'sd0.04794233341655642, 32'sd0.03118731997409257, 32'sd0.07576912656093149, 32'sd0.024731031354946986, 32'sd0.11673410811406325, 32'sd-0.08236370593580704, 32'sd-0.11478150925379652, 32'sd0.12896648885558726, 32'sd-0.019212112989555778, 32'sd-0.05565546170016213, 32'sd-0.10995068842448025, 32'sd-0.06307260137078555, 32'sd0.08621662345301194, 32'sd0.011170444722383053, 32'sd0.017357258863508248, 32'sd-0.09330214648245858, 32'sd-0.03830414744873933, 32'sd-0.03400358942459837, 32'sd-0.13925151487967566, 32'sd-0.04761548694262176, 32'sd0.017101394861126978, 32'sd0.10287807571111222, 32'sd0.1349241885845651, 32'sd0.00718281643899851, 32'sd0.032379180393576075, 32'sd0.02407779708572036, 32'sd-0.06471998192956864, 32'sd0.11816393364506292, 32'sd0.09684960081207876, 32'sd0.11254085121849557, 32'sd0.1306167526341015, 32'sd0.06491719533037721, 32'sd0.05894879061684683, 32'sd-0.02580041238234817, 32'sd0.06136071346032056, 32'sd0.06499387822229692, 32'sd-0.09976827812684287, 32'sd-0.033639691101519285, 32'sd-0.08303091812309027, 32'sd0.01234790477156906, 32'sd-0.031273149558645, 32'sd-0.055350538077137156, 32'sd-0.08346562054753688, 32'sd-0.1598550832867787, 32'sd-0.041942340760762364, 32'sd0.06135749442949583, 32'sd0.027243918281212434, 32'sd0.08713756731791107, 32'sd-0.03894799183085737, 32'sd0.08972044108480297, 32'sd-0.03211596146947191, 32'sd0.03449330091995451, 32'sd-0.09029455387163812, 32'sd-0.013006434043310424, 32'sd0.1198098718232106, 32'sd-0.007132406202413562, 32'sd0.08025293863332685, 32'sd0.18975229471169983, 32'sd0.34008033661182435, 32'sd0.1329436325482191, 32'sd0.0019935167018224286, 32'sd-0.06792577153684538, 32'sd0.05103851396232588, 32'sd-0.00024287868059552422, 32'sd-0.060126581755904455, 32'sd-0.02621736380738257, 32'sd0.05904461406079692, 32'sd-0.00890933230422941, 32'sd-0.009740174466366547, 32'sd-0.041087050323840024, 32'sd0.05082403442889693, 32'sd-0.04512601961439792, 32'sd0.0015116784605508525, 32'sd0.026961481368529674, 32'sd-0.005130037745567505, 32'sd-0.01828291300477719, 32'sd0.060487991725712155, 32'sd0.052537118792478875, 32'sd-0.05204947410344765, 32'sd-0.07763791254461742, 32'sd-0.15615478848468928, 32'sd-0.10131885191427126, 32'sd0.06336420096313383, 32'sd-0.08047501639174533, 32'sd0.14084513532157752, 32'sd0.12453863055397643, 32'sd0.19596584461142005, 32'sd0.0319275720452302, 32'sd-0.06441156645933899, 32'sd-0.14605942083040926, 32'sd0.040676677035745804, 32'sd0.012300395434625511, 32'sd-0.07794964147271939, 32'sd0.015865503173336053, 32'sd0.061091235247493894, 32'sd0.007259478891535545, 32'sd-0.061177300756360097, 32'sd0.0032225168222011977, 32'sd0.09296911696480782, 32'sd-0.13375490121141653, 32'sd-0.03606643376188722, 32'sd-0.22125104880341648, 32'sd-0.07176679973242814, 32'sd0.08272821579037085, 32'sd0.07617571257666336, 32'sd0.09873580640501861, 32'sd0.002938700768548109, 32'sd-0.01258476512087425, 32'sd-0.21404631800162272, 32'sd0.0002879532486139067, 32'sd0.11110223903437294, 32'sd-0.03967761349296725, 32'sd0.13419874800929563, 32'sd0.1371022577200639, 32'sd0.03165221417571691, 32'sd0.006486287948567787, 32'sd-0.08124113581242676, 32'sd-0.0024038640644936794, 32'sd-0.02082020347941774, 32'sd0.09214774451826784, 32'sd-0.08251797973565703, 32'sd7.624865376059979e-127, 32'sd-0.06881570781968516, 32'sd-0.018714614131671907, 32'sd-0.015225271909908787, 32'sd0.039789811415734164, 32'sd0.04724472249454743, 32'sd-0.17866675973859997, 32'sd-0.1767840847666214, 32'sd-0.15423734223888289, 32'sd0.034695050141432135, 32'sd0.11529879474488389, 32'sd-0.1164824012125907, 32'sd-0.08251936783013226, 32'sd0.041144249104836085, 32'sd-0.0037477939345686973, 32'sd-0.032494775818301555, 32'sd0.1033398834230661, 32'sd0.09759414404434452, 32'sd0.05372262308364537, 32'sd0.025712321079531992, 32'sd-0.07107402730643106, 32'sd-0.029072082055660874, 32'sd-0.10873823694427213, 32'sd-0.15329944135435083, 32'sd-0.014267963321420968, 32'sd-0.01810496580969566, 32'sd-0.06718131930585146, 32'sd-0.09706010452686326, 32'sd-0.0759959109588607, 32'sd0.04290610189355551, 32'sd0.11559631634600155, 32'sd0.04177385404435835, 32'sd-0.1369787656638851, 32'sd0.11820992484626786, 32'sd-0.006571502121928871, 32'sd-0.17374872138777903, 32'sd-0.008617667352874999, 32'sd-0.06680275250817673, 32'sd-0.013688828669407209, 32'sd0.008782576378415225, 32'sd-0.04703398886473817, 32'sd-0.1179683928660593, 32'sd-0.05770838037889559, 32'sd0.0791609227314155, 32'sd0.12694536757909072, 32'sd0.11758491578801988, 32'sd0.015950517544300512, 32'sd0.08436155041413108, 32'sd-0.07617914936947182, 32'sd0.022848447026046298, 32'sd0.0014959738475557702, 32'sd-0.026624676474316603, 32'sd-0.08261026532782928, 32'sd0.01425191234476842, 32'sd-0.08745007234828088, 32'sd-0.10233578192440605, 32'sd0.04256872123232506, 32'sd-0.050044132488645254, 32'sd-0.008589287241601929, 32'sd0.09414445807552614, 32'sd-0.07162384608495183, 32'sd0.12921199975400205, 32'sd0.01742943649182976, 32'sd0.06653362863750123, 32'sd0.025497588719212604, 32'sd0.07161617076726791, 32'sd-0.02997484669163039, 32'sd-0.07301154634390158, 32'sd-0.05382891968547252, 32'sd-0.13875749572959464, 32'sd0.015672295948390664, 32'sd0.15180940941365922, 32'sd0.11726500989751551, 32'sd-0.10877901132632378, 32'sd0.08351407607232537, 32'sd-0.0429231738009906, 32'sd-0.08936907871370808, 32'sd-0.04898688702389023, 32'sd-0.09778204312575048, 32'sd-0.04977536354247995, 32'sd-0.06956824506788732, 32'sd0.0733010501378795, 32'sd0.009276312567944459, 32'sd-0.03885823117350079, 32'sd-1.2863822033723277e-128, 32'sd0.01864262447072096, 32'sd0.06555430542995369, 32'sd0.035548542318493984, 32'sd-0.02498439372951644, 32'sd0.08561696961752281, 32'sd-0.027410137038070475, 32'sd0.02945064651738462, 32'sd0.03058645635532239, 32'sd0.0007921020405861234, 32'sd-0.02835156424415429, 32'sd-0.07547624343312376, 32'sd0.0678849373315767, 32'sd-0.10655680384628688, 32'sd-0.032200613932651896, 32'sd0.026153794971239347, 32'sd0.02041817285832516, 32'sd0.08978619328710852, 32'sd-0.02569551051762529, 32'sd-0.02389323453423898, 32'sd0.034081241884890395, 32'sd-0.027246213159497535, 32'sd-0.08603010961362378, 32'sd-0.007690081649157198, 32'sd-0.06667132312485588, 32'sd-0.012084906541847623, 32'sd-0.012223315746240611, 32'sd-0.09611634400965598, 32'sd-0.06958961664732664, 32'sd-0.0364466989782107, 32'sd0.023840111638826513, 32'sd0.036444683898639654, 32'sd-0.0789122642997939, 32'sd-0.021024723105818734, 32'sd0.0660131747163653, 32'sd-0.010448298398874062, 32'sd-0.12054851214434532, 32'sd-0.05315608533202723, 32'sd-0.02783406355303566, 32'sd-0.07377897288868975, 32'sd0.044425740011197215, 32'sd0.11314724470097284, 32'sd0.04450987641790167, 32'sd0.06206400657263311, 32'sd-0.05913825404697863, 32'sd-0.07363385193203396, 32'sd-0.10132138579146024, 32'sd0.07168575229039505, 32'sd0.03715597088163866, 32'sd-0.017526128622094357, 32'sd-0.1564515161731509, 32'sd-0.06633214674727081, 32'sd-0.06956343743505375, 32'sd0.02314917391246495, 32'sd0.13437024150257484, 32'sd-0.07825545099991497, 32'sd-0.05782567721294592, 32'sd0.059965785313113, 32'sd0.07997616677293232, 32'sd0.04350418598822674, 32'sd-0.08954207422561075, 32'sd0.03182394417511194, 32'sd-0.0412393990781192, 32'sd-0.04693403075918776, 32'sd0.022061941509847003, 32'sd-0.0178183807051885, 32'sd0.09438064901667124, 32'sd-0.03914698312080884, 32'sd0.04767352535381318, 32'sd0.13381944978725605, 32'sd0.06498655078234883, 32'sd0.048902812602829644, 32'sd-0.09782799365077186, 32'sd-0.10813004293450619, 32'sd-0.07309898682155941, 32'sd-0.049102697045244795, 32'sd0.03340902948086188, 32'sd-0.018925285672779305, 32'sd-0.028082737738351935, 32'sd-0.1488930382524532, 32'sd-0.09591242010530414, 32'sd0.08171950522658077, 32'sd0.1126969659546926, 32'sd-0.02456039245035545, 32'sd-1.7062692811027293e-120, 32'sd-0.06035461602086657, 32'sd0.01868391666462675, 32'sd-0.036006745621944815, 32'sd-0.015204634441837794, 32'sd-0.04622119827514127, 32'sd-0.021659184518226304, 32'sd0.05132568145579952, 32'sd-0.009876196745365128, 32'sd-0.026594635461356122, 32'sd0.034480399328873174, 32'sd0.12773883299315456, 32'sd0.0964735163560131, 32'sd0.07285458971860088, 32'sd-0.057219034018531206, 32'sd-0.10706039318721597, 32'sd-0.09781242946821156, 32'sd-0.029182076526232753, 32'sd0.023999931494596144, 32'sd0.046009913376283115, 32'sd0.06997648901405214, 32'sd-0.0340971301812449, 32'sd-0.007570639937884, 32'sd0.004267014377707582, 32'sd-0.09406704507529018, 32'sd0.07072855929522345, 32'sd-0.0073054006526956485, 32'sd-4.561229231443897e-121, 32'sd-3.2104210698039924e-116, 32'sd1.9162502289927136e-120, 32'sd0.07260562597517775, 32'sd-0.017071929155836423, 32'sd-0.02049945024985712, 32'sd-0.013410769802922072, 32'sd-0.08379045315326326, 32'sd0.016353590825486305, 32'sd0.03582976142877997, 32'sd-0.08536849160481082, 32'sd0.007830212731883985, 32'sd-0.018664881693231123, 32'sd0.00457041624163964, 32'sd0.017197324820426456, 32'sd-0.05148205733433323, 32'sd-0.02950472203878719, 32'sd0.02833074486268804, 32'sd-0.019827785530365526, 32'sd-0.14485611749679428, 32'sd0.018365840288673038, 32'sd0.11325257507895035, 32'sd0.15602005037762692, 32'sd-0.028401226579176573, 32'sd-0.05458973985132996, 32'sd-0.005549683716397921, 32'sd0.06074636477972705, 32'sd-0.06282594705546787, 32'sd-2.912609936453799e-119, 32'sd-4.950043002167074e-120, 32'sd-2.2891972975730553e-121, 32'sd-0.07597987711974225, 32'sd-0.05684408294511658, 32'sd-0.058373771084971646, 32'sd-0.07887876061923013, 32'sd-0.12267243259032284, 32'sd-0.09671445007032439, 32'sd0.005847710961200395, 32'sd0.02794980195392625, 32'sd0.06899589548445398, 32'sd0.014799944679178667, 32'sd0.0006162491016903703, 32'sd0.10445245887168751, 32'sd0.0273656420302173, 32'sd-0.01104733325818578, 32'sd-0.05848018827562798, 32'sd-0.03347211185983056, 32'sd-0.23073503660702926, 32'sd0.018590703702418627, 32'sd0.05388831743724801, 32'sd0.1295066325342325, 32'sd0.008457518167605942, 32'sd-0.018566719706062506, 32'sd0.09246879871878573, 32'sd-0.09418791316140825, 32'sd-0.006351023737453631, 32'sd1.6430621345655413e-127, 32'sd1.0355889377761584e-124, 32'sd1.000383152495513e-120, 32'sd-1.190355259813687e-117, 32'sd-0.00651623823403769, 32'sd0.001338392847364161, 32'sd-0.16443810185423902, 32'sd-0.0982695313399051, 32'sd-0.11535056246575535, 32'sd0.1261602690246752, 32'sd-0.016552115294437963, 32'sd0.07097006593095173, 32'sd-0.032626312789061515, 32'sd-0.1308660846638633, 32'sd-0.12510390018370204, 32'sd0.003973913254241298, 32'sd-0.11744371634937133, 32'sd-0.03520825626367104, 32'sd-0.027087577224886694, 32'sd-0.01511494946378483, 32'sd-0.11805864952937717, 32'sd-0.0749706304432751, 32'sd-0.011623374474269402, 32'sd0.06467767008555292, 32'sd0.09986520712473963, 32'sd0.024709091926007752, 32'sd-0.030516478383803336, 32'sd1.5214859669905388e-125, 32'sd-2.6220168801005922e-124, 32'sd3.7855977612015953e-116, 32'sd3.4260798061207525e-126, 32'sd-1.1531871613675568e-125, 32'sd-1.0345874945173118e-120, 32'sd-0.09567811319078257, 32'sd0.03533330719045764, 32'sd-0.009872106995543818, 32'sd-0.0762266016116265, 32'sd-0.009743250639464357, 32'sd-0.005637574421010219, 32'sd-0.14871874367778523, 32'sd-0.05649460625139312, 32'sd-0.08355518564089538, 32'sd-0.09292489005571515, 32'sd-0.1352589666560656, 32'sd-0.131326275262266, 32'sd-0.07704047486239783, 32'sd-0.08472858518976563, 32'sd-0.06293873734143585, 32'sd-0.03253371407879957, 32'sd0.0020052329323635484, 32'sd0.09639204010417589, 32'sd-0.02930105159884817, 32'sd0.08561281343808845, 32'sd-2.5077053517986403e-126, 32'sd8.528982800556768e-121, 32'sd-1.6725854729629784e-117, 32'sd-3.457049845391082e-122},
        '{32'sd-1.1317428282312199e-126, 32'sd2.1303028154421862e-125, 32'sd-7.525490279233655e-115, 32'sd-4.880330166174032e-126, 32'sd-1.9642080684713097e-125, 32'sd-9.41593782215934e-123, 32'sd7.566223004201544e-115, 32'sd-5.817900063036632e-126, 32'sd-3.331523999426374e-121, 32'sd6.57633123593295e-117, 32'sd5.772520358704667e-121, 32'sd-1.296477809835835e-118, 32'sd-0.05309240869890956, 32'sd0.041976891253649055, 32'sd0.06449919018146844, 32'sd0.05296041588273043, 32'sd7.84576223954554e-127, 32'sd3.093630280641874e-118, 32'sd1.4217022941311293e-118, 32'sd1.2050167703749482e-116, 32'sd-7.529021998684318e-115, 32'sd-7.644761719771832e-126, 32'sd2.966731035534611e-127, 32'sd4.057330310916482e-115, 32'sd1.7886587774948575e-128, 32'sd-3.0808429919322537e-125, 32'sd-1.8491208117765885e-123, 32'sd-6.166238457210224e-122, 32'sd-1.21394054662775e-116, 32'sd-9.035114111515205e-119, 32'sd6.740035383938693e-115, 32'sd4.711790689296628e-115, 32'sd0.013115416809189043, 32'sd0.09225979222554659, 32'sd0.005581341510098351, 32'sd-0.10786564994636119, 32'sd-0.0016798252858599735, 32'sd-0.10156276552261058, 32'sd-0.10156123227562219, 32'sd0.010807489932540744, 32'sd0.052621161618082606, 32'sd-0.049468971274777306, 32'sd0.04560078391847434, 32'sd-0.006412737300019504, 32'sd0.14152916484565384, 32'sd0.08336639943727427, 32'sd0.08391027280217347, 32'sd0.002361197737098404, 32'sd0.028185588219800675, 32'sd0.10474032027422964, 32'sd0.10350972283802724, 32'sd0.012526011756974261, 32'sd-2.4316188908794805e-118, 32'sd-3.9662350386709104e-119, 32'sd-2.326124019250897e-120, 32'sd-2.7706459285244137e-118, 32'sd-1.925696931794575e-114, 32'sd-3.20100797397463e-119, 32'sd0.02119269749697674, 32'sd0.05589015310229857, 32'sd0.024557857019268315, 32'sd0.030382147991574068, 32'sd0.009668382129943254, 32'sd0.1092815345282914, 32'sd0.02086482533631808, 32'sd-0.1412921238500624, 32'sd-0.15034134535270852, 32'sd-0.14024358856598684, 32'sd-0.008989079151926184, 32'sd-0.08849856239802947, 32'sd0.05800814932931406, 32'sd0.027824623469052647, 32'sd0.06531210334456268, 32'sd0.1535046440315293, 32'sd0.030785872497954725, 32'sd0.12571191032145193, 32'sd0.11922787499510244, 32'sd-0.033985494004023405, 32'sd0.037176539900644956, 32'sd0.006591232852799458, 32'sd-0.017219034730825058, 32'sd-0.012953999278851406, 32'sd-9.189386417369735e-125, 32'sd6.19475001137563e-122, 32'sd9.253195960865798e-123, 32'sd-1.9570154323721525e-124, 32'sd0.0035983978866459686, 32'sd0.07942908036569772, 32'sd0.05242651836373312, 32'sd-0.0693181493346584, 32'sd0.008657995054613286, 32'sd-0.01050204606609146, 32'sd-0.015688344434973963, 32'sd0.005899217561488869, 32'sd-0.07735442629004789, 32'sd0.019216332103259744, 32'sd0.11548796931796304, 32'sd0.11670719209004488, 32'sd0.009201239087933091, 32'sd0.06556621869134734, 32'sd0.05002393738205408, 32'sd-0.04423219885873129, 32'sd-0.03893782868930147, 32'sd-0.158356173346546, 32'sd-0.02635159093521016, 32'sd0.012109896900355513, 32'sd-0.06941588401014692, 32'sd0.01610815976611428, 32'sd-0.055876887577133334, 32'sd-0.059537677526299175, 32'sd0.007909248568512968, 32'sd-4.3410689780799416e-122, 32'sd1.4827282746981978e-122, 32'sd0.016820298925755296, 32'sd0.059790208015586266, 32'sd0.023325749730476526, 32'sd0.041605424401274356, 32'sd0.015919502486738298, 32'sd-0.03506152845181866, 32'sd-0.11564422679631664, 32'sd0.021851372721705935, 32'sd0.06982269488187247, 32'sd0.10554048610156866, 32'sd-0.06771876752498844, 32'sd-0.0789786254960309, 32'sd0.04645257471529087, 32'sd0.11115726507194257, 32'sd-0.05139139645418795, 32'sd0.06265858505485544, 32'sd0.006077504189228962, 32'sd-0.09031249035555235, 32'sd-0.05030087014090007, 32'sd-0.15169231783257842, 32'sd-0.11417787636430467, 32'sd-0.0024019201394737807, 32'sd-0.11493811749201144, 32'sd-0.08691864651905702, 32'sd-0.0423616235819676, 32'sd0.03632970257856513, 32'sd0.02534404866789344, 32'sd-9.263283656899897e-128, 32'sd0.007624736001529247, 32'sd0.06582739229823292, 32'sd0.04613909348646271, 32'sd0.04129345198708986, 32'sd0.07638553047677325, 32'sd0.04504852032178454, 32'sd0.00303431423408055, 32'sd-0.04766648226877826, 32'sd0.008798368773110625, 32'sd-0.07250445622742266, 32'sd-0.005280699857693438, 32'sd0.022077776510281148, 32'sd-0.08229980507892153, 32'sd0.06698398122577018, 32'sd0.020116221519766445, 32'sd0.011295568783514663, 32'sd-0.04468422436827567, 32'sd-0.16488122574868072, 32'sd0.0077502147557927635, 32'sd0.022360204181277106, 32'sd-0.043515942972330184, 32'sd-0.07159797674307454, 32'sd-0.09963198690951822, 32'sd-0.0009344028789570412, 32'sd0.004992651082396918, 32'sd-0.11208721966019249, 32'sd0.05461528449180517, 32'sd1.586121896446269e-123, 32'sd-0.01257075206726785, 32'sd0.0007710015102469287, 32'sd0.0829925803297286, 32'sd-0.09426727730503916, 32'sd0.05119740473349717, 32'sd0.10747706418590686, 32'sd0.05750198589384588, 32'sd0.04065382650626495, 32'sd-0.09460766730510085, 32'sd-0.17527491335104647, 32'sd-0.03609802296512066, 32'sd0.021508400800798112, 32'sd-0.06387818983107, 32'sd0.0035751457621438346, 32'sd-0.10786239978159962, 32'sd-0.034275490305373926, 32'sd-0.16117923899307446, 32'sd-0.08468211385684198, 32'sd-0.02891511831854712, 32'sd-0.06740544972846783, 32'sd-0.07375149769405641, 32'sd-0.1017605529443845, 32'sd0.019477761402398597, 32'sd0.05267325483626128, 32'sd0.08161487610326505, 32'sd-0.06748506292164554, 32'sd-0.058418682215057305, 32'sd-0.007455265782048868, 32'sd0.03222864119873557, 32'sd0.0006538424605263085, 32'sd0.01437966791326098, 32'sd-0.030294107473913066, 32'sd-0.00029999038445663177, 32'sd-0.043705940945679714, 32'sd-0.03011132070225014, 32'sd0.033201258782713045, 32'sd-0.02002231382914644, 32'sd-0.05285441447019318, 32'sd0.08879719978248422, 32'sd-0.015997081341303634, 32'sd-0.11319936220304191, 32'sd-0.1527728688711003, 32'sd-0.1352070439719696, 32'sd-0.17328137708902017, 32'sd-0.06906107578656759, 32'sd-0.170959235316143, 32'sd-0.07546777550671747, 32'sd-0.06457112220217902, 32'sd0.024747699596226587, 32'sd-0.01613846105096916, 32'sd-0.14321069011566906, 32'sd-0.022847428931120985, 32'sd0.019791732357614247, 32'sd-0.10534904643374317, 32'sd0.05438066622378255, 32'sd0.037633349640026785, 32'sd0.07129426138922364, 32'sd-0.013412044297096117, 32'sd-0.003661899837622629, 32'sd-0.04197267609414622, 32'sd0.05261358059985947, 32'sd0.0012022978250845842, 32'sd-0.0015901903510481662, 32'sd0.03560719791107139, 32'sd-0.024275968174569198, 32'sd0.1034399668182821, 32'sd0.046759811962238516, 32'sd-0.019706469711720125, 32'sd-0.12603917207443, 32'sd-0.22417638557052127, 32'sd-0.22517793822970453, 32'sd-0.20175413845790283, 32'sd-0.14526850548711673, 32'sd-0.20407934525501434, 32'sd-0.12242744599329376, 32'sd0.029166071318245633, 32'sd0.012560114352392005, 32'sd-0.13312055629888517, 32'sd-0.008382751256010686, 32'sd-0.06620575222596496, 32'sd0.026666418472021242, 32'sd0.022227879899195245, 32'sd-0.06503325880896128, 32'sd-0.03908901130349219, 32'sd-0.078151342201218, 32'sd0.06781744005268941, 32'sd-0.12011489803464552, 32'sd-0.07017461691648542, 32'sd-0.08392490188399192, 32'sd-0.04363627378101705, 32'sd0.08766783335480319, 32'sd-0.04826211078528554, 32'sd0.03124748303947218, 32'sd-0.012283108899934265, 32'sd0.0606441532054282, 32'sd0.016002211531494434, 32'sd-0.099031437517134, 32'sd-0.12063667128510835, 32'sd-0.12469426551800353, 32'sd0.012549638085677342, 32'sd-0.06407859616784387, 32'sd-0.12207632532368072, 32'sd0.004767951024301559, 32'sd0.0586216328544751, 32'sd0.05435994330312278, 32'sd-0.02688516197593758, 32'sd-0.08230168643877456, 32'sd0.03662067338437129, 32'sd-0.10472801149897396, 32'sd0.007917923426740761, 32'sd0.004751522853375823, 32'sd0.01076050404098976, 32'sd0.047403866161353246, 32'sd0.04701027132303242, 32'sd-0.13632899001000318, 32'sd-0.11544033712256534, 32'sd-0.005941335923269738, 32'sd0.0666410474326657, 32'sd-0.002054521165119791, 32'sd0.07003577142473229, 32'sd0.014342069963603167, 32'sd0.020249427297662263, 32'sd0.07840105676183722, 32'sd0.1313965408703833, 32'sd-0.08385624336053278, 32'sd-0.07100368738036386, 32'sd0.019115641750837027, 32'sd0.13343410594171365, 32'sd0.079922150415864, 32'sd-0.04587149234599337, 32'sd0.07377845724095033, 32'sd0.009439005859331981, 32'sd0.0007703578671026563, 32'sd-0.040842300463354464, 32'sd-0.018436882567297457, 32'sd0.12905499405301707, 32'sd-0.016334858031351786, 32'sd0.004806462554573121, 32'sd0.02507430677675895, 32'sd-0.05386811597031422, 32'sd0.13063861765108278, 32'sd-0.10622413099248444, 32'sd-0.16247111100515316, 32'sd-0.10950296035871677, 32'sd-0.01600444505333894, 32'sd0.052285451773158804, 32'sd-0.04770575518388474, 32'sd0.0670844288048122, 32'sd0.10153297559917467, 32'sd-0.06489779890830678, 32'sd-0.06505358623848483, 32'sd-0.07809402251206085, 32'sd-0.07860816944847764, 32'sd-0.09598275483246657, 32'sd0.06400450301901728, 32'sd0.08769745001103951, 32'sd0.00435232103886968, 32'sd0.09032287845583369, 32'sd0.026785046560378566, 32'sd0.08672548690833107, 32'sd0.09546273054876597, 32'sd-0.03527098124728495, 32'sd0.028851018067744396, 32'sd0.03926209384851739, 32'sd0.065503396843692, 32'sd-0.02957916979134009, 32'sd-0.11154359910352224, 32'sd0.0258076828179039, 32'sd0.04152178502028945, 32'sd-0.151629325216909, 32'sd-0.0707000640998764, 32'sd0.05886381783831685, 32'sd0.07165411484834429, 32'sd0.02856400141579827, 32'sd-0.03988984182252566, 32'sd0.04474027449900726, 32'sd0.024746789361749035, 32'sd-0.017239911604357346, 32'sd0.042701700755703176, 32'sd-0.1317243769207997, 32'sd0.012465142588406652, 32'sd0.0371843583585755, 32'sd-0.025137543521535723, 32'sd0.08898450004212377, 32'sd-0.07768770833137006, 32'sd-0.023289905261205356, 32'sd-0.07395326566532755, 32'sd0.11973655238594445, 32'sd0.05121384655259062, 32'sd0.034263259435462066, 32'sd0.005270683173140893, 32'sd-0.014909412643086473, 32'sd0.0357801200987774, 32'sd-0.009970374967212205, 32'sd-0.07795061446650804, 32'sd0.00033349634731805704, 32'sd-0.0266192987886748, 32'sd-0.11035896985299135, 32'sd-0.14295623274535857, 32'sd-0.07365296697158787, 32'sd-0.0030340430722897794, 32'sd-0.09105519070549847, 32'sd-0.1259734959883026, 32'sd-0.11509465478311928, 32'sd-0.06307181691367235, 32'sd-0.10119465374580065, 32'sd-0.12436750582010259, 32'sd-0.03872841825291198, 32'sd0.006752465966384623, 32'sd0.020744561444937373, 32'sd-0.03153311823276503, 32'sd0.0012570539352180087, 32'sd-0.09652863336213012, 32'sd0.04701782031386192, 32'sd-0.008384992615709705, 32'sd0.0544690624787337, 32'sd0.1684895935281223, 32'sd0.10157378981341839, 32'sd0.07768885412172008, 32'sd-0.08748711418719107, 32'sd-0.08102789809097127, 32'sd0.04446770871462696, 32'sd-0.022066902759702255, 32'sd-0.031083138174599144, 32'sd-0.041742794892347175, 32'sd-0.05656839028361474, 32'sd0.0189016664734436, 32'sd-0.14736919224594733, 32'sd0.008928875946221628, 32'sd-0.011832186307387001, 32'sd-0.1331977787550901, 32'sd-0.02979137253917309, 32'sd-0.08448929207601313, 32'sd-0.018966462403451297, 32'sd-0.017991390116920025, 32'sd0.02596648670228643, 32'sd0.15107366694471067, 32'sd0.19703302622280583, 32'sd0.09752663358855461, 32'sd0.008154272431558073, 32'sd-0.10656710184800175, 32'sd-0.11761707597413838, 32'sd0.051476949691007357, 32'sd0.052563274278945644, 32'sd0.03181590107496019, 32'sd0.04704592865952337, 32'sd-0.03948072316837086, 32'sd-0.013748913205250408, 32'sd0.07033416949557715, 32'sd-0.016004818995939904, 32'sd-0.002116719306763419, 32'sd0.058165347669319654, 32'sd0.05746564108339029, 32'sd-0.057998644177614175, 32'sd0.04362216307601951, 32'sd0.018747543737748867, 32'sd0.04776975734014054, 32'sd0.029155615982317324, 32'sd-0.010991201406982095, 32'sd-0.04242138184315809, 32'sd-0.049693198062831484, 32'sd-0.12207234476060128, 32'sd-0.13945695896476037, 32'sd0.021928801200798344, 32'sd0.26712399843891166, 32'sd0.19300357994303474, 32'sd0.13406290136954135, 32'sd0.015760533696030764, 32'sd-0.15269939876801733, 32'sd-0.07130298378443828, 32'sd0.0010391278855417445, 32'sd0.028566345316435662, 32'sd0.030892729936385917, 32'sd0.03181183196967939, 32'sd-0.0020009931020587247, 32'sd0.014324857331163527, 32'sd0.04224310774534554, 32'sd0.04171933176332102, 32'sd0.057048763903792224, 32'sd-0.003180648860026318, 32'sd-0.03364619140095638, 32'sd-0.051087989980929366, 32'sd0.009042458493056653, 32'sd0.02098477107822756, 32'sd0.022526821603972357, 32'sd-0.0704295955860978, 32'sd-0.09837434877737211, 32'sd-0.0541964994707141, 32'sd-0.06879905560765093, 32'sd-0.06815595147129705, 32'sd0.06077342157298999, 32'sd0.06726261930664403, 32'sd0.03473029952781321, 32'sd0.17052417533493253, 32'sd0.24743207362171343, 32'sd0.013817710724891956, 32'sd0.06669957035208841, 32'sd0.044887485540073095, 32'sd0.05419874892928954, 32'sd0.03760384043215471, 32'sd0.019106321767475867, 32'sd-0.012823323395256504, 32'sd0.01148048535018039, 32'sd-0.12012265720398631, 32'sd0.02762943597171175, 32'sd0.029213389369447486, 32'sd-0.019590162395239783, 32'sd1.2426094561227862e-125, 32'sd0.018067388975948655, 32'sd-0.0541748151878438, 32'sd0.0556004399039504, 32'sd0.024246933832576433, 32'sd-0.11008538892902738, 32'sd-0.07187539996364983, 32'sd-0.2509262229759039, 32'sd-0.1062523752402663, 32'sd-0.05466853844902781, 32'sd-0.025876104866483566, 32'sd0.0028000487874341308, 32'sd0.10181577790585203, 32'sd-0.06811276751868621, 32'sd0.047788348358256724, 32'sd0.19772519635116367, 32'sd0.10087082705094122, 32'sd0.0971442414334256, 32'sd0.14553097450686137, 32'sd0.05646849709449323, 32'sd0.062167993412073526, 32'sd-0.05859915172009893, 32'sd0.06569818307905433, 32'sd0.016030225394734716, 32'sd0.10564395391366507, 32'sd0.05703384274828078, 32'sd-0.03828468242870991, 32'sd0.022403920854785302, 32'sd0.0748406685955546, 32'sd-0.0031018709174124204, 32'sd0.08305196692121614, 32'sd0.016432911997359325, 32'sd-0.05835245374783426, 32'sd-0.11952565835101714, 32'sd-0.1578635989202131, 32'sd-0.02018587261072022, 32'sd0.09381310040387376, 32'sd0.07551604858962364, 32'sd0.01974934358689954, 32'sd-0.08383848393664772, 32'sd0.06296345517559093, 32'sd-0.09372113157359843, 32'sd0.1646226564356855, 32'sd0.11972896018592119, 32'sd-0.004802990237202882, 32'sd-0.0244344763247968, 32'sd0.050125991923614006, 32'sd-0.05425605467246668, 32'sd-0.08501561181665315, 32'sd0.06624354783248289, 32'sd-0.009194474867027833, 32'sd0.07649157257359183, 32'sd0.1022843027355042, 32'sd0.11434539182217661, 32'sd-0.09414955203907473, 32'sd0.0005044999137317057, 32'sd0.02667884200347484, 32'sd-0.028985251832003133, 32'sd0.021417219068059653, 32'sd0.08891764458074135, 32'sd-0.07705653113711304, 32'sd-0.13058227421474886, 32'sd-0.183410269321255, 32'sd0.038916917355069136, 32'sd0.11218410937839228, 32'sd0.09659099052445588, 32'sd0.17155474217043143, 32'sd0.08297369598048115, 32'sd-0.07966099513749277, 32'sd-0.03253584414513033, 32'sd-0.014762515924384554, 32'sd0.11295430579630836, 32'sd0.0786413418465531, 32'sd0.08363689465698657, 32'sd0.08184348242134779, 32'sd-0.04686622749802849, 32'sd0.054460879220293114, 32'sd0.07686332850429455, 32'sd-0.030817408284240518, 32'sd0.11078071017747249, 32'sd0.06472317748162998, 32'sd-0.00015803527877730525, 32'sd0.020232308276071035, 32'sd0.12189336218186743, 32'sd-4.50161369538622e-121, 32'sd-0.09495549183746708, 32'sd0.059696441397826774, 32'sd0.027553451967730153, 32'sd-0.12217699412969243, 32'sd-0.2157972812137283, 32'sd-0.08390362715333904, 32'sd-0.009662372927617837, 32'sd-0.04758522229338928, 32'sd0.04712363303009126, 32'sd0.1897082592531943, 32'sd0.18482778756507035, 32'sd0.006472125170381996, 32'sd0.006784542255983101, 32'sd-0.04019989227993777, 32'sd0.04519922033466415, 32'sd0.03196598167309437, 32'sd0.002164075636122362, 32'sd0.17242124071875745, 32'sd0.12359250303235095, 32'sd0.15314277656481276, 32'sd-0.0017966690406971578, 32'sd-0.008683910700968312, 32'sd-0.024531714428711163, 32'sd0.10995681465749299, 32'sd-0.015613768378859262, 32'sd-0.05882538299177142, 32'sd0.028130245257212697, 32'sd-0.00046941912987271284, 32'sd0.02413657068654108, 32'sd0.01637521155062697, 32'sd0.049435056951983476, 32'sd0.013681168867869917, 32'sd-0.10315683740506447, 32'sd-0.0715206939029274, 32'sd-0.058885727443700756, 32'sd0.10897709987065451, 32'sd0.13690065959480321, 32'sd0.11995498356721272, 32'sd-0.05871057220149455, 32'sd-0.08649667660100988, 32'sd0.1046749524495778, 32'sd0.0828565861729324, 32'sd-0.028206525818248607, 32'sd0.04661323167187191, 32'sd0.15618514197661038, 32'sd0.053580183361899784, 32'sd0.01829668173202994, 32'sd0.04423414637737677, 32'sd-0.022777800466852308, 32'sd-0.12632208618143023, 32'sd-0.13832594311423832, 32'sd0.011544805280207184, 32'sd0.04653040826165498, 32'sd-0.11249148762183762, 32'sd0.03586459732290628, 32'sd-0.0007671082054833042, 32'sd0.01090954386405747, 32'sd-0.04282962316345713, 32'sd-0.054052084191167596, 32'sd0.03538279408042953, 32'sd0.030191062521482924, 32'sd-0.07321461894408703, 32'sd-0.1513498147272184, 32'sd0.006891643370743431, 32'sd-0.07944701279416358, 32'sd-0.01740409730305651, 32'sd-0.0808752296518828, 32'sd-0.0380737502182542, 32'sd0.03532819792981777, 32'sd0.01938798609316261, 32'sd-0.13665019017618002, 32'sd-0.04751937564735695, 32'sd-0.01854717729921516, 32'sd-0.07085278477931993, 32'sd-0.07850432732961374, 32'sd-0.10269557461347922, 32'sd-0.043145560377250244, 32'sd-0.004747640792193423, 32'sd-0.06780654274243159, 32'sd-0.10959438433696239, 32'sd0.08895640001620128, 32'sd-0.07911188847964597, 32'sd0.05823666880921876, 32'sd-2.173077414443189e-122, 32'sd0.028598583353437693, 32'sd-0.0946840901976716, 32'sd-0.047393371749996895, 32'sd-0.028912010230350702, 32'sd-0.03965748726935757, 32'sd-0.08321139112446449, 32'sd-0.12298875170250154, 32'sd-0.0573951317524405, 32'sd-0.06240466773657055, 32'sd-0.07311151379576193, 32'sd-0.11058850091531561, 32'sd0.034260349440934826, 32'sd0.10492212031249887, 32'sd-0.06218272658037337, 32'sd-0.05144280108562079, 32'sd-0.11978357489901005, 32'sd-0.07042452179556757, 32'sd-0.2009548724550815, 32'sd-0.18637536419009426, 32'sd0.04179333175221233, 32'sd0.020534716004694593, 32'sd-0.03665392005189501, 32'sd-0.09545239434675278, 32'sd-0.04389518316471537, 32'sd0.03768088202759237, 32'sd0.02256342692431577, 32'sd-1.1144373958688701e-119, 32'sd1.5643110344271939e-115, 32'sd-3.1684985708719718e-114, 32'sd0.009109662372999186, 32'sd-0.02231685550224128, 32'sd0.10705571787565352, 32'sd-0.06857616558936301, 32'sd-0.01460988766588655, 32'sd-0.12254824069862368, 32'sd-0.056913789743398814, 32'sd0.04856600914392876, 32'sd-0.01720164321979959, 32'sd-0.10258240235006376, 32'sd-0.1608488086982794, 32'sd-0.13430939002510747, 32'sd-0.025366754314988478, 32'sd-0.08646810281546422, 32'sd-0.06989373991829094, 32'sd-0.09124373589800956, 32'sd-0.12762277414924647, 32'sd-0.14797301116175363, 32'sd-0.12057681828875508, 32'sd0.007160828444437699, 32'sd-0.11273979674306081, 32'sd-0.12313188114066159, 32'sd-0.004755108153224189, 32'sd-0.018585086206166276, 32'sd-0.012134147713409454, 32'sd1.6311848164649468e-121, 32'sd7.542922815559836e-118, 32'sd-1.0240434393353163e-121, 32'sd0.02555020185598146, 32'sd0.04420123991847769, 32'sd-0.06430666419977625, 32'sd-0.08075847863453785, 32'sd-0.0018654250888824613, 32'sd0.037491231135100535, 32'sd-0.0043531725401520106, 32'sd-0.028400799886748616, 32'sd-0.03960461440890472, 32'sd-0.041227167149241205, 32'sd-0.08614386459236012, 32'sd-0.22099922150365517, 32'sd-0.034799308651377224, 32'sd-0.09652782316007393, 32'sd-0.12352984720862428, 32'sd-0.1938812620543497, 32'sd-0.11369040023262858, 32'sd0.009660819670132942, 32'sd-0.024172566820862607, 32'sd-0.05419622369131614, 32'sd-0.08080810394025317, 32'sd0.02639341068859196, 32'sd-0.05697726224398211, 32'sd0.014723932920511858, 32'sd0.03282015988444786, 32'sd-1.2391116162579486e-126, 32'sd-2.299370943341399e-124, 32'sd4.06345885675668e-123, 32'sd8.936728831190897e-123, 32'sd-0.006928816535009397, 32'sd-0.0698430565831998, 32'sd0.03623340604590886, 32'sd-0.03637850553890008, 32'sd0.07564303667809961, 32'sd-0.08684437898524879, 32'sd0.03915002454737993, 32'sd-0.09053698946712396, 32'sd0.004366554136111886, 32'sd-0.0241656532767094, 32'sd-0.08084369938298888, 32'sd-0.1806686164745172, 32'sd-0.07946244318802043, 32'sd0.11803754480421139, 32'sd0.08282495631407752, 32'sd-0.0758619777796539, 32'sd-0.04739998198805491, 32'sd-0.0769249442668074, 32'sd-0.07703883178605236, 32'sd-0.06104147439145819, 32'sd-0.0021083672071202666, 32'sd0.014417385563567423, 32'sd0.0021506482469460194, 32'sd-6.25698872869844e-124, 32'sd8.624117811787232e-117, 32'sd-1.3228275758770654e-122, 32'sd3.233125027793071e-123, 32'sd-4.721374435384015e-124, 32'sd-1.6316354872248826e-126, 32'sd0.04494873730303353, 32'sd-0.013129457254853705, 32'sd0.040929854391494144, 32'sd0.021900084908488895, 32'sd0.021011069807560002, 32'sd-0.04513190574547683, 32'sd0.026960100543224643, 32'sd-0.0008510578669297719, 32'sd-0.023612888440959514, 32'sd0.05343071145163556, 32'sd0.045611170703442575, 32'sd0.09885660064566335, 32'sd0.05495983953602206, 32'sd0.06152598346758133, 32'sd0.02688486212277302, 32'sd0.023552583101304727, 32'sd0.0045944406936588725, 32'sd-0.036823027921469964, 32'sd-0.0015522919146586133, 32'sd-0.025972644572806902, 32'sd1.2559547606815866e-125, 32'sd9.444911089204732e-122, 32'sd1.6526012020180413e-124, 32'sd8.597481410069199e-117},
        '{32'sd-2.471987211232893e-119, 32'sd-1.2839122961057626e-119, 32'sd2.979445797349639e-120, 32'sd6.703898746252551e-124, 32'sd-6.739965611882024e-123, 32'sd6.88204236997238e-126, 32'sd-2.682127442324296e-124, 32'sd3.863255597718587e-119, 32'sd1.0375571700543838e-120, 32'sd-2.283877162108609e-123, 32'sd-1.2881047543704808e-123, 32'sd1.785611227597389e-121, 32'sd0.010324233959586088, 32'sd-0.04846144121698561, 32'sd0.032851526055508486, 32'sd-0.030307495531758863, 32'sd8.668944181066622e-120, 32'sd6.864487980729378e-126, 32'sd-2.9698676251597006e-124, 32'sd-8.164136160222177e-121, 32'sd-1.5001702345119276e-115, 32'sd3.5011236558751344e-123, 32'sd-8.927437190355137e-124, 32'sd3.185336396427675e-119, 32'sd-4.378855515672406e-118, 32'sd8.745715623084342e-120, 32'sd5.731600738294518e-120, 32'sd1.3416176305290805e-120, 32'sd2.529871539485218e-126, 32'sd-2.5866361377415657e-124, 32'sd-8.681230050224724e-119, 32'sd1.2759462571591991e-122, 32'sd0.06289387603494051, 32'sd-0.006057646591552921, 32'sd-0.003086914326067879, 32'sd0.015861839895297308, 32'sd0.00840652258582209, 32'sd0.03646442446522706, 32'sd0.02811928562702369, 32'sd0.015498603055809848, 32'sd0.06968774843195659, 32'sd-0.08387949783396473, 32'sd-0.010230167293764428, 32'sd0.02334391387195249, 32'sd0.09440515243063863, 32'sd-0.024972791593344455, 32'sd0.056733765228187405, 32'sd0.011664936181501068, 32'sd0.022204579124078572, 32'sd-0.010610622686720729, 32'sd-0.01976519372139952, 32'sd0.03447700992083084, 32'sd6.953509461490014e-124, 32'sd2.2629387405227467e-114, 32'sd-1.7557983846325223e-116, 32'sd2.822141206612364e-121, 32'sd9.429894824094147e-120, 32'sd-3.441351857838139e-127, 32'sd0.04099063793663813, 32'sd-0.016586972897598237, 32'sd0.058392435061011036, 32'sd0.04418771241300999, 32'sd-0.08991791336696195, 32'sd-0.06651099671398457, 32'sd-0.065669884595103, 32'sd-0.020009856133062193, 32'sd-0.07948764860980907, 32'sd0.048392285920011796, 32'sd0.04796824817593705, 32'sd0.006762570380322444, 32'sd0.07573487890475797, 32'sd-0.06975645002593217, 32'sd-0.04388172617704322, 32'sd0.038241009084393075, 32'sd-0.05596537841824699, 32'sd0.03944004257611372, 32'sd0.08499351958514474, 32'sd0.03516322837771581, 32'sd0.008697877347011098, 32'sd0.060654675323939554, 32'sd-0.016245204983316733, 32'sd0.06100321059829698, 32'sd-5.5113583969835215e-121, 32'sd6.97765658473592e-123, 32'sd6.498868381913645e-126, 32'sd4.7436055836262e-124, 32'sd0.06492743914779811, 32'sd0.025067439704877667, 32'sd0.0004258961588633746, 32'sd-0.032066058190346594, 32'sd-0.014496959390796194, 32'sd-0.03153924002288326, 32'sd-0.006631542959622328, 32'sd0.008478860356009742, 32'sd0.09751024817902675, 32'sd0.05777767932067619, 32'sd0.0013516450430515069, 32'sd0.03155889339295201, 32'sd0.00585381153462516, 32'sd0.03819128647660243, 32'sd-0.062059189277865225, 32'sd0.06837708738450017, 32'sd0.043466616743564064, 32'sd0.04608279672085311, 32'sd-0.04769474447011051, 32'sd-0.12639264485175042, 32'sd-0.07676369497841098, 32'sd-0.06557675250336165, 32'sd-0.0540418047653397, 32'sd-0.020473980029848564, 32'sd0.01795107303765671, 32'sd4.882696203310981e-124, 32'sd-1.5093095090446394e-127, 32'sd0.047133900992988094, 32'sd-0.0048130052035042495, 32'sd0.06646672263468328, 32'sd-0.04664641761705618, 32'sd0.038089410295763765, 32'sd-0.05786079170337296, 32'sd-0.046505507435634315, 32'sd-0.09727289414053818, 32'sd0.035225505466440286, 32'sd0.05259233430537621, 32'sd-0.014490109994666015, 32'sd0.057132854920091465, 32'sd-0.01330180862348458, 32'sd0.07850067737377711, 32'sd0.054470243286421936, 32'sd0.03145777776136484, 32'sd-0.049684903315177754, 32'sd0.024379458637916008, 32'sd0.025500500398104572, 32'sd-0.09800376931258321, 32'sd0.008867645761588692, 32'sd0.08299233619377007, 32'sd0.0013165902384575333, 32'sd-0.06107786839043562, 32'sd-0.13757422560343624, 32'sd-0.0708182115194487, 32'sd0.012574036538874412, 32'sd-1.281669237606699e-123, 32'sd-0.010783882324691399, 32'sd-0.07034461419586897, 32'sd-0.05569043821785993, 32'sd0.018783095076975197, 32'sd0.05846469782485462, 32'sd-0.12410231545305238, 32'sd-0.19016082416631988, 32'sd-0.07217446110530719, 32'sd-0.04547437623378762, 32'sd-0.06560205266791133, 32'sd0.07034225228341295, 32'sd-0.040494723398543264, 32'sd-0.12279556373821418, 32'sd-0.12399758976075859, 32'sd-0.05937896288314729, 32'sd-0.10566978420187448, 32'sd-0.02701398226739901, 32'sd-0.09717474377561226, 32'sd0.030748025495000053, 32'sd-0.08553766244871029, 32'sd-0.04372788405148935, 32'sd0.062320120686769835, 32'sd-0.058462052191888825, 32'sd-0.07757074079701175, 32'sd-0.06802076630133755, 32'sd-0.09620178802289403, 32'sd0.002658062410443275, 32'sd-7.059620418801569e-127, 32'sd0.014922469437797651, 32'sd-0.0746218610523896, 32'sd-0.07628506688487968, 32'sd-0.031897751601679514, 32'sd0.1378062583788809, 32'sd0.0547910209651621, 32'sd-0.09538550652788284, 32'sd-0.05887084646605342, 32'sd-0.1456420549604964, 32'sd-0.03439818593438517, 32'sd0.1167479451002736, 32'sd0.1385520008768779, 32'sd-0.0474652003235659, 32'sd-0.10122776893208606, 32'sd-0.2762248869212814, 32'sd-0.022626672477705206, 32'sd-0.08383219809391569, 32'sd-0.08321584590525441, 32'sd-0.0304047754922741, 32'sd0.0802019042875601, 32'sd0.0396732526135802, 32'sd0.0720947090557025, 32'sd-0.014943213566876369, 32'sd-0.08722158602273354, 32'sd-0.017695010075157582, 32'sd-0.01470701678473311, 32'sd0.032956046561386086, 32'sd-0.008166485631524984, 32'sd0.03330894298837643, 32'sd-0.017901510393794423, 32'sd-0.06474110588713249, 32'sd-0.010070489008205463, 32'sd0.06222950573032339, 32'sd0.10454911292595194, 32'sd-0.0861599685799782, 32'sd-0.17042010315274916, 32'sd0.09758807608120755, 32'sd0.03640615254655544, 32'sd0.2167770513140066, 32'sd0.13118484281064766, 32'sd-0.06714053637699631, 32'sd-0.009258149224222807, 32'sd-0.19514808107257045, 32'sd-0.19467103878440634, 32'sd-0.05217111977814892, 32'sd-0.038865130816981966, 32'sd0.15465386563855277, 32'sd0.04871315557752495, 32'sd0.006696947473901776, 32'sd0.04468090010032653, 32'sd0.06310331113737239, 32'sd0.04324091017775794, 32'sd-0.10188702267154008, 32'sd-0.009361290992089162, 32'sd-0.06261513729017326, 32'sd-0.01770301975108993, 32'sd-0.09069621416136325, 32'sd-0.09118464448311, 32'sd0.016275395046746532, 32'sd-0.08931384932598145, 32'sd-0.021714112036509043, 32'sd0.08166858123748086, 32'sd0.11306661363320854, 32'sd-0.14950899990011837, 32'sd0.022332014243621103, 32'sd0.07279848411629768, 32'sd0.08904940184739196, 32'sd0.0075088461076780215, 32'sd-0.09659244371897446, 32'sd-0.15838039990136799, 32'sd-0.13538383242937563, 32'sd-0.13396216326646126, 32'sd0.06456155883943922, 32'sd0.0473565316230484, 32'sd0.16562308927961875, 32'sd0.16393462448114518, 32'sd0.06551354325917394, 32'sd-0.014875052717284551, 32'sd-0.039939084865941825, 32'sd0.058230926377228556, 32'sd0.0131050830797905, 32'sd-0.05776281592005427, 32'sd-0.008275184850761376, 32'sd0.04276878269143921, 32'sd-0.02876732722220552, 32'sd-0.0940537076783401, 32'sd-0.026900372306935403, 32'sd-0.13302816088485878, 32'sd-0.1222767316612284, 32'sd-0.0298942341948889, 32'sd-0.03577461759991588, 32'sd-0.06741385239471079, 32'sd-0.0394027806396159, 32'sd0.09643985693329385, 32'sd0.12383736329323293, 32'sd0.13058570550770993, 32'sd-0.07491064713751922, 32'sd-0.1589773964961973, 32'sd-0.08995492937740035, 32'sd0.06541136185093954, 32'sd0.09373463610766548, 32'sd0.04070573181215546, 32'sd0.033172343031103974, 32'sd0.05512008442924865, 32'sd0.10878360599758517, 32'sd-0.06506882803681895, 32'sd-0.10668510262765377, 32'sd-0.01115371534924713, 32'sd-0.11338613916456429, 32'sd-0.08540286073104077, 32'sd-0.03902297563729615, 32'sd0.04072800529781803, 32'sd0.0631410261988912, 32'sd0.03556648211560505, 32'sd-0.03779460853099734, 32'sd0.022379940264247666, 32'sd-0.061195049271389225, 32'sd-0.09844001651231579, 32'sd-0.026474633003374114, 32'sd-0.11020470551823766, 32'sd0.0652554965223908, 32'sd0.13318517926749013, 32'sd0.20379596510944722, 32'sd0.2117649416592513, 32'sd-0.0051257646135596515, 32'sd-0.07557784751079076, 32'sd-0.07097149345562603, 32'sd-0.17738640095116562, 32'sd0.029444378046130964, 32'sd0.007069756218174829, 32'sd0.05791029549012771, 32'sd-0.08494697695611533, 32'sd-0.00567816550165506, 32'sd-0.07659781854834088, 32'sd-0.10486441318287165, 32'sd-0.007356024524387509, 32'sd0.1809068228302831, 32'sd-0.10736121256183916, 32'sd0.08618018535064212, 32'sd0.08244413872987807, 32'sd-0.002753179016693258, 32'sd0.019380585993165465, 32'sd-0.08729892041198367, 32'sd-0.01700315331899095, 32'sd-0.050755410739953495, 32'sd0.03965713812956784, 32'sd-0.1730925700855911, 32'sd-0.14880441071488104, 32'sd-0.046047485798401296, 32'sd0.05842495657209736, 32'sd-0.0036764448293845533, 32'sd0.00381411713290904, 32'sd-0.041621695650952695, 32'sd-0.06967706945662921, 32'sd-0.016660466198472126, 32'sd-0.0029322959124100036, 32'sd0.027240592577847805, 32'sd-0.015658207416664148, 32'sd-0.13040834934818418, 32'sd-0.04526675127095689, 32'sd-0.09233059939167328, 32'sd-0.13942472280111617, 32'sd-0.11396879690257584, 32'sd-0.07206014554477543, 32'sd-0.01926960460578493, 32'sd0.035739698658100345, 32'sd0.02468842749269222, 32'sd0.02567313349197552, 32'sd-0.007271213257714425, 32'sd-0.016179673407889044, 32'sd-0.0033147511021208356, 32'sd-0.19370429853191887, 32'sd-0.10294490226825172, 32'sd-0.06089497343015626, 32'sd-0.055251748494943756, 32'sd-0.06749801718796512, 32'sd-0.004354255911398243, 32'sd-0.013772111696935877, 32'sd0.09911633173646582, 32'sd0.022338551337674477, 32'sd0.0371163355656294, 32'sd0.12236732529228377, 32'sd0.05206378100313377, 32'sd0.018380935165458245, 32'sd0.017922458330887462, 32'sd-0.12032586459479479, 32'sd-0.17686193029815392, 32'sd-0.0027681876578067983, 32'sd-0.04402538843000417, 32'sd-0.10998259217915458, 32'sd-0.01742875528120142, 32'sd0.050103532728715844, 32'sd0.038684674634083656, 32'sd0.04683012634638044, 32'sd0.008269015507922304, 32'sd0.01373675057837281, 32'sd-0.02907702016672356, 32'sd-0.09757816563421487, 32'sd-0.11137722323124188, 32'sd-0.1540727267633703, 32'sd0.03597931734238839, 32'sd-0.06897581314675161, 32'sd0.03492440022870488, 32'sd0.011130374960891734, 32'sd0.004639041842224572, 32'sd0.006520536430408161, 32'sd0.1355936033386895, 32'sd0.08364137184535471, 32'sd0.059915551157072575, 32'sd0.10424433566048696, 32'sd0.1374593812111519, 32'sd0.06746027225016443, 32'sd0.09106888875840762, 32'sd-0.07399181117666216, 32'sd-0.10242542617824694, 32'sd0.0018281484994073505, 32'sd0.008112709556467784, 32'sd0.09755827848624114, 32'sd0.055453467362242374, 32'sd0.07625588696126472, 32'sd-0.11057528991920504, 32'sd-0.09513158837806988, 32'sd0.03776967392303786, 32'sd0.026499848468161093, 32'sd0.004672390596117501, 32'sd-0.007848465030696278, 32'sd-0.00870307439215297, 32'sd-0.03596926127553439, 32'sd0.05206013101293519, 32'sd-0.058572852929389185, 32'sd-0.06209174854318576, 32'sd0.015169830013461276, 32'sd-0.0386328244870414, 32'sd-0.07310061328830611, 32'sd-0.025512981655189112, 32'sd0.07091947484561247, 32'sd0.014317220294606501, 32'sd0.19116748808340414, 32'sd0.11562389970256545, 32'sd-0.023143487777707986, 32'sd-0.09205518622083486, 32'sd-0.03298772630428589, 32'sd0.004795124455569012, 32'sd-0.008601502804974648, 32'sd-0.08663506170992136, 32'sd-0.023602189105343965, 32'sd0.039372234901019564, 32'sd-0.050948666653499064, 32'sd-0.031041936135920375, 32'sd-0.04231275156587039, 32'sd-0.08128165602659612, 32'sd0.08345342534135633, 32'sd-0.017758988802306214, 32'sd-0.10015771465328377, 32'sd0.0728725320475788, 32'sd-0.009893311882513262, 32'sd-0.046845775992292234, 32'sd-0.012840286634340836, 32'sd-0.03045860683997439, 32'sd-0.07603611771497172, 32'sd-0.08280623643884097, 32'sd0.08531901126790477, 32'sd-0.014825214407410834, 32'sd0.03881995203933231, 32'sd-0.060632714200874946, 32'sd0.05219515285049804, 32'sd0.06276549694856921, 32'sd0.044468343765242085, 32'sd0.031167083635367174, 32'sd-0.03343419008087472, 32'sd0.04821533095572699, 32'sd0.005869088953757197, 32'sd-0.07176243998437695, 32'sd0.01601839185847351, 32'sd0.03570145964326144, 32'sd-0.014636710884839532, 32'sd-0.060900834240716545, 32'sd-0.0990833886649286, 32'sd0.022581978416474472, 32'sd-2.7244587398921172e-05, 32'sd0.031700346450323484, 32'sd-0.13684529214429247, 32'sd0.008806259502982219, 32'sd0.050652623875664826, 32'sd0.04610190056892875, 32'sd0.04422281450814868, 32'sd0.046135284653606376, 32'sd-0.004586146763232652, 32'sd-0.042621897471347515, 32'sd-0.08570225086711704, 32'sd-0.11936248607629658, 32'sd0.030591825257584422, 32'sd-0.0010141608779796168, 32'sd0.056347577572630723, 32'sd0.17613723300424833, 32'sd0.103195776071758, 32'sd-0.0036068895267662967, 32'sd-0.007569214471897723, 32'sd0.031451350074891415, 32'sd-0.06922498256748276, 32'sd0.10362283800107507, 32'sd-0.03639252386893142, 32'sd-0.013456667237910233, 32'sd-0.18623220355931444, 32'sd-0.09792995347665384, 32'sd-0.08756400924312611, 32'sd-0.008183754670873958, 32'sd2.842581798485633e-119, 32'sd0.034684787251950656, 32'sd-0.06606009254925872, 32'sd-0.04123200039139033, 32'sd0.08770882697502616, 32'sd0.02092067073278719, 32'sd0.11651154081818976, 32'sd0.02084500555617491, 32'sd0.03861022056924756, 32'sd-0.0025369412462839186, 32'sd-0.11377924084856143, 32'sd-0.15502964330388114, 32'sd-0.14495728418516207, 32'sd0.08786418574585289, 32'sd0.09919513348579427, 32'sd0.13976689878881246, 32'sd0.09025434998327424, 32'sd-0.055549777520737205, 32'sd-0.054948802177404374, 32'sd-0.1518721194555557, 32'sd-0.050638507189532174, 32'sd-0.009154032406897633, 32'sd-0.08359716097768573, 32'sd-0.0504651158072524, 32'sd-0.032689637168816496, 32'sd0.004353595676666021, 32'sd0.021564751253938422, 32'sd-0.07404757385624991, 32'sd0.04786312754206415, 32'sd0.07338451661805759, 32'sd-0.016951127677222115, 32'sd0.035943921161184895, 32'sd0.03483937573123516, 32'sd0.04091161355648249, 32'sd-0.09756968971322441, 32'sd-0.06557289299517452, 32'sd-0.05005946452765383, 32'sd-0.13881852467769576, 32'sd-0.04246467597404545, 32'sd-0.16560366894590878, 32'sd-0.1457229244420884, 32'sd0.10370158434052679, 32'sd0.08748596360853131, 32'sd0.02600527461058175, 32'sd0.10665046139110408, 32'sd-0.11796996880551902, 32'sd-0.0596361946499166, 32'sd0.0903881030340926, 32'sd0.11168949712435554, 32'sd-0.003029150398291333, 32'sd-0.11501171484496778, 32'sd-0.04544198120408254, 32'sd-0.0736995780127541, 32'sd-0.08602455701652015, 32'sd-0.02552642114877972, 32'sd0.04533413337248449, 32'sd0.038578661680983374, 32'sd-0.07661455172169516, 32'sd0.04470677527346672, 32'sd0.011902355827223111, 32'sd-0.09504773317311457, 32'sd-0.07387674571327298, 32'sd-0.18348811652489852, 32'sd-0.02809112072145557, 32'sd-0.05152199665358036, 32'sd-0.024446723492007532, 32'sd-0.1877746317703757, 32'sd-0.19669099887938982, 32'sd-0.20259043397191928, 32'sd-0.022903620248077346, 32'sd0.0994348536711399, 32'sd0.06485943851343726, 32'sd0.07198679139784891, 32'sd-0.007708888951495728, 32'sd-0.0683066182759423, 32'sd-0.006033024967874752, 32'sd0.05358904780664846, 32'sd-0.12776702145613988, 32'sd-0.09068386801179426, 32'sd-0.1775014818643829, 32'sd-0.0046122639536814065, 32'sd0.08387358243755737, 32'sd-0.06853183066224915, 32'sd0.04521413253473161, 32'sd-3.5074676356342164e-126, 32'sd-0.0010509349008255473, 32'sd0.027166748934014717, 32'sd0.014995484270314179, 32'sd-0.056831226815244745, 32'sd-0.06051842863654156, 32'sd-0.11423421531457521, 32'sd-0.15398462337652363, 32'sd-0.03674341629210551, 32'sd-0.09032704757893019, 32'sd-0.10304204849702857, 32'sd-0.096809406613128, 32'sd-0.014388453463018177, 32'sd-0.12716047341595343, 32'sd0.037094624231710324, 32'sd0.08592264444607528, 32'sd0.050326669167900205, 32'sd-0.034295755010815505, 32'sd0.04457426434321468, 32'sd0.04523383939143921, 32'sd-0.06252379430698968, 32'sd-0.20969584065397032, 32'sd-0.02584398282199836, 32'sd-0.08368528054553973, 32'sd-0.06922976315709231, 32'sd0.05675488604680825, 32'sd-0.04518214547320253, 32'sd0.0440718526396911, 32'sd0.03910246599902435, 32'sd0.04875769473457801, 32'sd0.094466799650861, 32'sd-0.035162182137970774, 32'sd0.002018106919849642, 32'sd0.06259988323357152, 32'sd-0.09411364171346288, 32'sd0.02107317544612215, 32'sd0.011175107645251928, 32'sd-0.00015921453975591487, 32'sd0.009600884992721666, 32'sd-0.06098747876813437, 32'sd0.0068131942137135346, 32'sd-0.09084733989415401, 32'sd0.05645467350986396, 32'sd0.1456083216936382, 32'sd-0.004338810475773, 32'sd0.015633232312542787, 32'sd0.07154877556062376, 32'sd0.0711721319870719, 32'sd-0.05855862611340893, 32'sd-0.07733709947338607, 32'sd-0.045444461237767755, 32'sd-0.01658052990544815, 32'sd0.07824587312743479, 32'sd0.0072963616668076, 32'sd-0.008578566149746898, 32'sd-0.01567990486354223, 32'sd0.03200244691534856, 32'sd0.10899196823675522, 32'sd-0.012206483009322268, 32'sd-0.017724206620377055, 32'sd0.09940225087357135, 32'sd0.11272945244200314, 32'sd0.047525276658377885, 32'sd-0.024936737109285196, 32'sd0.010045377910930797, 32'sd-0.04520873494432053, 32'sd-0.017953162407603154, 32'sd0.0922605004426851, 32'sd0.018241389683609104, 32'sd-0.03321075279715933, 32'sd-0.09228263060999439, 32'sd0.04755976238465748, 32'sd0.06933747831496663, 32'sd-0.0386581581665663, 32'sd0.12036415458297872, 32'sd-0.06774860859177431, 32'sd-0.02988277857031533, 32'sd-0.03419205800812217, 32'sd-0.12015403893857333, 32'sd0.030463034699172192, 32'sd0.10671325550142763, 32'sd-0.0677701910987634, 32'sd0.0139027031767921, 32'sd0.02006302364132956, 32'sd5.704888909833532e-118, 32'sd0.03908243707160425, 32'sd0.05300573511842238, 32'sd-0.025008496600809203, 32'sd0.05885695988557521, 32'sd0.11334753076295523, 32'sd0.07112167941635973, 32'sd0.07275030194725388, 32'sd0.015039839120455072, 32'sd0.09479685157886383, 32'sd0.042110478274203965, 32'sd-0.009206026582827227, 32'sd-0.0015986701407486358, 32'sd0.04248243577936828, 32'sd-0.10055167345874301, 32'sd0.024596017972581034, 32'sd0.1060564048665203, 32'sd0.008669711154411312, 32'sd0.00786452178539001, 32'sd0.02200346136278297, 32'sd-0.049706975451154975, 32'sd0.09389627496212696, 32'sd0.0240958166946977, 32'sd0.004371891122916338, 32'sd-0.015336845382152811, 32'sd-0.03363872472044304, 32'sd-0.038948601793686644, 32'sd-7.770721669817988e-125, 32'sd1.2812849731199874e-115, 32'sd1.4927977759121926e-117, 32'sd0.021106528745860012, 32'sd-0.09048918133916156, 32'sd-0.06178808747083429, 32'sd0.024952127203333816, 32'sd-0.08296832297179373, 32'sd-0.01607214822113686, 32'sd-0.0004861504819649105, 32'sd0.1200903695452392, 32'sd-0.0361266344994614, 32'sd-0.044695028215325575, 32'sd0.02498201104701246, 32'sd-0.07065526681145388, 32'sd-0.1940184400667573, 32'sd-0.13445710641655848, 32'sd-0.02937829328568124, 32'sd-0.06991453054829816, 32'sd0.07371879847963968, 32'sd-0.01245295872042482, 32'sd0.07285885901482458, 32'sd-0.014059302911071487, 32'sd0.024158203228767015, 32'sd-0.016454568416084527, 32'sd-0.0035549958121091417, 32'sd0.02201904582601728, 32'sd0.0029643721867906804, 32'sd3.938712299254607e-121, 32'sd-1.3301726905901488e-126, 32'sd6.920467521602352e-121, 32'sd-0.021336821337154678, 32'sd-0.02368440374365842, 32'sd-0.03763424054589833, 32'sd-0.011844237739634703, 32'sd0.005853208158484318, 32'sd0.06860143471295237, 32'sd0.045336754915170314, 32'sd0.0594999408493785, 32'sd-0.06755339130374978, 32'sd-0.08919583211631929, 32'sd0.023644305055831986, 32'sd0.007191039931879476, 32'sd0.07926490264531741, 32'sd0.04098320075868157, 32'sd-0.013284845049387957, 32'sd-0.18526029832531046, 32'sd-0.02260924745917737, 32'sd-0.061951563340819686, 32'sd-0.01983841523407767, 32'sd-0.02124866439936182, 32'sd-0.01004414731239339, 32'sd-0.020887883629144156, 32'sd0.0388869408576278, 32'sd-0.0060240093838369695, 32'sd0.022957616240840698, 32'sd1.033484019341135e-117, 32'sd2.446739284874442e-124, 32'sd-1.4806280655386043e-117, 32'sd5.406043313363137e-118, 32'sd0.016021547829558103, 32'sd-0.0240067289473247, 32'sd-0.07453614811144343, 32'sd-0.07715435005850876, 32'sd-0.0008247499612919147, 32'sd0.08625232982484574, 32'sd-0.04428567099942735, 32'sd0.03437983560817559, 32'sd-0.024229542958360818, 32'sd-0.12561746779481767, 32'sd-0.2107153082403665, 32'sd-0.12517350651757073, 32'sd-0.18056094763996142, 32'sd0.0698072532421461, 32'sd0.08270278453869716, 32'sd-0.13299098106355173, 32'sd-0.06736971234788172, 32'sd0.010177484423453557, 32'sd0.0626454333198484, 32'sd-0.13213931669703777, 32'sd-0.005302426135575083, 32'sd0.03146039627641073, 32'sd-0.03838351209856335, 32'sd2.8918069514322767e-124, 32'sd6.449889627095274e-125, 32'sd5.367600632066392e-118, 32'sd7.43551005865449e-127, 32'sd-3.354806160184157e-120, 32'sd6.843529725095803e-126, 32'sd0.037998048571887884, 32'sd-0.00294188826552252, 32'sd0.04180571818200647, 32'sd0.06752836441650913, 32'sd-0.09574898897734249, 32'sd-0.00706188500344572, 32'sd-0.040627277499205264, 32'sd-0.046514526297191626, 32'sd-0.03965782634604719, 32'sd-0.04064763488694401, 32'sd-0.038564416154579964, 32'sd-0.02693031700920692, 32'sd-0.02868872033923326, 32'sd-0.006883446436503786, 32'sd0.05803356570690049, 32'sd-0.003975830463763209, 32'sd0.12021047902474498, 32'sd-0.032958191954718406, 32'sd-0.04463219672849858, 32'sd0.027251966655243202, 32'sd-1.6058876066526428e-115, 32'sd-1.1862470805763829e-117, 32'sd-3.695123958250809e-126, 32'sd6.399539835691115e-126}
    };

    localparam logic signed [31:0] layer0_biases [0:127] = '{
        32'sd-0.1274994600276725, 32'sd-0.003646774188560244, 32'sd-0.16192743681966934, 32'sd0.08888217424466142, 32'sd-0.1207546770002809, 32'sd0.05803170772379196, 32'sd-0.006783942540424067, 32'sd-0.1115440861277134, 32'sd-0.14291038276818901, 32'sd-0.06647181287754239, 32'sd0.0012949793965979228, 32'sd-0.07302080777802811, 32'sd-0.004665507798726913, 32'sd-0.10229298136792793, 32'sd0.006731991123545049, 32'sd-0.006053089393871269, 32'sd0.01577932996450472, 32'sd-0.04910846172625988, 32'sd-0.04439189848869223, 32'sd0.022326044234423623, 32'sd-0.15052743291898707, 32'sd-0.040498149186010475, 32'sd-0.03587981532198645, 32'sd-0.031080787917183526, 32'sd0.012796973253402089, 32'sd0.008533689585010497, 32'sd-0.022504421093454397, 32'sd-0.0035268285551300817, 32'sd-0.14411727788595954, 32'sd-0.043939291758134255, 32'sd-0.08899949748458673, 32'sd0.04198122663663008, 32'sd-0.12076629843185153, 32'sd-0.1281421977871082, 32'sd-0.025049643453214775, 32'sd-0.06725399910082135, 32'sd0.08803948573845596, 32'sd-0.11241570751544426, 32'sd-0.027304628676563664, 32'sd-0.030349169078289735, 32'sd-0.02013842711809301, 32'sd-0.0757804403680299, 32'sd0.006559094756808764, 32'sd0.043798322779020904, 32'sd-0.18649961839716703, 32'sd-0.08629198039563002, 32'sd-0.09253991059043938, 32'sd-0.10174260132323143, 32'sd-0.03651596266996245, 32'sd-0.04055648387934882, 32'sd-0.08087449946351523, 32'sd-0.16036305508639329, 32'sd-0.10323910144640676, 32'sd-0.1570358100144523, 32'sd-0.12460371179664088, 32'sd-0.08482082695240674, 32'sd0.03817038508456822, 32'sd0.08181228091424238, 32'sd-0.15965268223906923, 32'sd-0.05120488004883541, 32'sd-0.09248119727421947, 32'sd-0.09010086427743642, 32'sd0.04621896508852529, 32'sd-0.052234453155004315, 32'sd-0.12870401860841665, 32'sd-0.10410683284618044, 32'sd0.07009245764449865, 32'sd-0.05198920116536711, 32'sd-0.05178026920206926, 32'sd-0.02852455112827102, 32'sd0.046015374531435976, 32'sd0.07582805985455515, 32'sd-0.04411987386463083, 32'sd-0.026226269462935926, 32'sd-0.03364041491860055, 32'sd-0.006988825380293652, 32'sd-0.017111049036087945, 32'sd0.09693538202456403, 32'sd-0.15549933690799836, 32'sd-0.03628769878596967, 32'sd-0.10990775974806131, 32'sd0.1433282508530998, 32'sd-0.18116806632139015, 32'sd-0.0471925714076758, 32'sd-0.03375451336760963, 32'sd-0.04678926534175538, 32'sd-0.0623609846620864, 32'sd-0.010967105581607859, 32'sd-0.11782739803803459, 32'sd-0.04875053202686785, 32'sd-0.13410120340031648, 32'sd-0.023124392087522226, 32'sd-0.25703731651113815, 32'sd-0.004044595443971369, 32'sd-0.11006231845424495, 32'sd-0.15076073302585766, 32'sd-0.22354359795271028, 32'sd-0.10498900764441685, 32'sd-0.1106700533678615, 32'sd-0.044132053081405685, 32'sd-0.10054440205822845, 32'sd-0.029404570476876557, 32'sd-0.11315368980100217, 32'sd-0.003176837251123398, 32'sd-0.23596995438667925, 32'sd-0.06426079525017096, 32'sd0.05710338377197297, 32'sd-0.13678692301957981, 32'sd-0.1281503967159463, 32'sd0.0730769816968679, 32'sd0.07266261164247616, 32'sd-0.02552069179272736, 32'sd-0.04497728816846758, 32'sd0.0053204659476943795, 32'sd-0.02045724441322341, 32'sd-0.09864582718829057, 32'sd-0.04565665816600751, 32'sd-0.06689352644502777, 32'sd-0.00792033309484825, 32'sd0.0504085076154707, 32'sd0.07535057826156415, 32'sd-0.10396417813747179, 32'sd-0.26607963068485185, 32'sd-0.10466365183019413, 32'sd0.08680842334081124, 32'sd-0.005226528412602603, 32'sd-0.00215683829602922, 32'sd-0.01680075971318795
    };

    //Layer 1: 128 inputs, 64 neurons
    localparam logic signed [31:0] layer1_weights [0:63][0:128] = '{
        '{32'sd-0.15273142326367378, 32'sd0.26149938626919655, 32'sd-0.10868876209618741, 32'sd-0.18777363880401537, 32'sd-0.10817528750446707, 32'sd0.05081522011408665, 32'sd0.09212760507142818, 32'sd-0.0017158409535134578, 32'sd-0.2560276148764181, 32'sd0.0057362177700067485, 32'sd0.05795883764901562, 32'sd-0.15042862389756986, 32'sd0.031908363963040906, 32'sd0.19012709291093013, 32'sd-0.07504375865604482, 32'sd0.18651678834743282, 32'sd0.0002002840681841636, 32'sd0.03029394214964148, 32'sd0.10103541914668707, 32'sd0.06788662076128217, 32'sd-0.10747226922803099, 32'sd0.1812604525660162, 32'sd-0.074334914638571, 32'sd-0.16076486491191935, 32'sd0.02477571970593909, 32'sd0.21619904770886764, 32'sd0.17232765576559947, 32'sd0.06513568777347803, 32'sd0.025771842124057975, 32'sd0.14300638021434173, 32'sd0.2770822112830966, 32'sd0.17505012001576825, 32'sd-0.10683349133009126, 32'sd0.009527390551789578, 32'sd-0.06643402741695614, 32'sd0.1396752246137521, 32'sd-0.040529338951676416, 32'sd-0.05843669366338652, 32'sd0.040474706538432464, 32'sd-0.15748164085450678, 32'sd0.004628545093690512, 32'sd0.09475015914424416, 32'sd-0.19446612681013137, 32'sd-0.0327718595624467, 32'sd0.05166593523057306, 32'sd-0.12330964166144898, 32'sd-0.10868356913252107, 32'sd-0.158744427951353, 32'sd0.05436067327487298, 32'sd-0.004638675561480709, 32'sd-0.09168545818954749, 32'sd-0.10394421372375426, 32'sd-0.019378735025439242, 32'sd-0.16948156294198455, 32'sd0.07720333779310315, 32'sd-0.3588063850461922, 32'sd-0.07959224596414503, 32'sd0.1967333230314521, 32'sd0.11352435855945654, 32'sd0.08119677752728405, 32'sd-0.17738037723175423, 32'sd0.00208921485505078, 32'sd-0.0008610629495081039, 32'sd0.036996907342511196, 32'sd0.02264086519614492, 32'sd0.026022122745923203, 32'sd-0.08198702687234448, 32'sd0.12648705999676554, 32'sd0.020081247751300175, 32'sd0.0077559165436248256, 32'sd0.10540827269235972, 32'sd0.2641216112698168, 32'sd0.15997519219612064, 32'sd0.04738142735489043, 32'sd0.229666711866095, 32'sd0.03293807455646622, 32'sd-0.13726225725759922, 32'sd0.11015411343160497, 32'sd-0.222255248802646, 32'sd0.03817738475273335, 32'sd-0.09437070241587468, 32'sd0.16617197476688372, 32'sd0.08649900392958584, 32'sd0.09175132721352916, 32'sd0.1225452935496609, 32'sd0.08998608460007972, 32'sd-0.03952152656244126, 32'sd0.16500006303020623, 32'sd-0.014082330414603217, 32'sd0.12797799262816337, 32'sd0.14507542705831927, 32'sd0.14869463846490955, 32'sd-0.07179521060174975, 32'sd-0.18247325775958848, 32'sd0.17713804066526317, 32'sd-0.20417201710105098, 32'sd0.11334509321466271, 32'sd-0.22311814251690715, 32'sd0.26009840613017854, 32'sd0.031381570488538464, 32'sd-0.11058697583506256, 32'sd-0.08789679698327575, 32'sd0.07723476513320032, 32'sd0.04090723903169519, 32'sd-0.004985513681630706, 32'sd0.26399321424058486, 32'sd-0.17186389046782283, 32'sd0.047869975420649115, 32'sd-0.0339468114553219, 32'sd0.17115151563455788, 32'sd-0.009556596496747088, 32'sd-0.21034363203347695, 32'sd0.12552715954059707, 32'sd0.07617406236504261, 32'sd-0.12255326215324826, 32'sd-0.00811383144265341, 32'sd0.2716154758950459, 32'sd-0.031533142552272, 32'sd0.2510185967919448, 32'sd0.03459594399168692, 32'sd0.06626759231152735, 32'sd-0.048864617112110785, 32'sd0.00911489613781678, 32'sd-0.07712990885758332, 32'sd0.18266952487783075, 32'sd0.15327592884317753, 32'sd0.15147641684344262, 32'sd0.12227384807235125},
        '{32'sd0.10975691960873556, 32'sd-0.14177829354090163, 32'sd-0.1252030755256691, 32'sd-0.10801236425749118, 32'sd-0.16908002627708196, 32'sd-0.15795111986449287, 32'sd-0.08850430284508505, 32'sd-0.208539913251069, 32'sd-0.19946627689138854, 32'sd-0.0997723560043654, 32'sd0.15253760161159385, 32'sd-0.16536480354213684, 32'sd-0.046287930622266375, 32'sd0.0652221182955053, 32'sd0.2791018802337828, 32'sd-0.09156927107127964, 32'sd0.20875900816128456, 32'sd-0.0814199390554192, 32'sd0.2048702522953877, 32'sd0.2002614545717881, 32'sd-0.191882199100007, 32'sd0.1442027242849568, 32'sd0.0685012819102546, 32'sd-0.26508275037841816, 32'sd0.17655707056497116, 32'sd0.004367978064092833, 32'sd0.1877305964245718, 32'sd0.23598279457441781, 32'sd-0.1737014685266447, 32'sd-0.07243268496007087, 32'sd0.12605116061623628, 32'sd0.0766257516564565, 32'sd0.146486918696988, 32'sd0.10890823448740848, 32'sd0.09909889696869312, 32'sd-0.16994382291384838, 32'sd-0.24203127561596374, 32'sd-0.08759584739418798, 32'sd-0.053612103214124886, 32'sd-0.04048826540698791, 32'sd-0.20800162406283015, 32'sd-0.10387474214566884, 32'sd0.19743758036298517, 32'sd0.21926206287975475, 32'sd-0.02761924727931787, 32'sd-0.15135388397725033, 32'sd-0.19812081859864916, 32'sd0.09672956992096603, 32'sd0.03551084808050983, 32'sd0.07131749155301448, 32'sd0.12903500818588107, 32'sd0.29953685407920566, 32'sd-0.03148126961093755, 32'sd-0.03309028786295232, 32'sd0.04042820030624025, 32'sd0.022500978314299497, 32'sd-0.16506493045979131, 32'sd-0.13355309707173924, 32'sd0.019571638764096806, 32'sd0.2541241574309458, 32'sd0.1457234219103149, 32'sd-0.10710160442378011, 32'sd-0.14598310071953002, 32'sd-0.09324169774138172, 32'sd-0.018782932881060723, 32'sd-0.024248664694464562, 32'sd-0.1576329441447806, 32'sd0.04994721874943533, 32'sd-0.09195088565936857, 32'sd0.05267792668026924, 32'sd-0.23312224377767093, 32'sd0.0038443054295855335, 32'sd0.1089628640180074, 32'sd0.13725118058170996, 32'sd-0.04032409569872764, 32'sd0.21113799539425362, 32'sd0.05885524231065797, 32'sd0.04249386276580053, 32'sd0.1745427209085622, 32'sd-0.010106419250333358, 32'sd0.1751317145716208, 32'sd-0.019339440227819735, 32'sd0.012737482634413903, 32'sd-0.03354689524232259, 32'sd-0.10611802011462776, 32'sd0.08533745664910075, 32'sd-0.12131218140527097, 32'sd-0.08468518978255861, 32'sd0.04290828853929029, 32'sd0.04517674584465726, 32'sd0.18612603608521563, 32'sd0.24929082926241486, 32'sd0.11597675313859127, 32'sd0.11612951893421164, 32'sd-0.11526688292488113, 32'sd0.06062393203522736, 32'sd-0.05368708741987141, 32'sd0.05090557465259694, 32'sd0.16245949334125315, 32'sd0.0938190483002193, 32'sd-0.037776449767807724, 32'sd0.09297096672275697, 32'sd-0.13783613536033626, 32'sd0.07645240238413765, 32'sd-0.10474544662921674, 32'sd0.021007245195354952, 32'sd-0.17693401525716165, 32'sd-0.11670644945199464, 32'sd-0.010836084445407493, 32'sd-0.004377073212913745, 32'sd-0.19360007065999657, 32'sd-0.16365764590750564, 32'sd0.06668445524130354, 32'sd0.02562514713819387, 32'sd0.14426640385874887, 32'sd-0.15510047536901259, 32'sd0.10557440994219226, 32'sd-0.08613936414635162, 32'sd0.17638757542018157, 32'sd-0.0020123754263379335, 32'sd0.004789343446348418, 32'sd0.0847054971488628, 32'sd0.14156459798337942, 32'sd-0.09615553225188557, 32'sd0.04396702982026821, 32'sd0.08278975949639007, 32'sd-0.046058992950848955, 32'sd-0.25904992919016745},
        '{32'sd0.10382804429021379, 32'sd0.08433036807022146, 32'sd-0.03766037621822127, 32'sd-0.13615644225104306, 32'sd-0.2846320280488836, 32'sd0.16690956609756372, 32'sd0.0962823776803214, 32'sd-0.013639114615588121, 32'sd0.18802270270692484, 32'sd0.04734136170291328, 32'sd0.0219194207979705, 32'sd-0.11457833818907846, 32'sd0.21904681489380973, 32'sd0.06371135566739726, 32'sd-0.0626979860521054, 32'sd-0.09520431693050001, 32'sd0.09455103199946047, 32'sd-0.024715113329419492, 32'sd0.028638270987968988, 32'sd-0.006966521846971074, 32'sd-0.03799005142339417, 32'sd-0.23193802384724713, 32'sd0.18948149929093427, 32'sd-0.19648869754200038, 32'sd0.21647166876835092, 32'sd-0.2190129586792082, 32'sd-0.013266190620600315, 32'sd-0.02437671345014064, 32'sd-0.1866432175848466, 32'sd0.06265115861006995, 32'sd-0.15377801905336416, 32'sd-0.17544581348763388, 32'sd0.052702379569915934, 32'sd-0.06008720724630219, 32'sd0.054234206597912046, 32'sd0.12982885797422852, 32'sd0.010169555081832236, 32'sd0.07398645552295896, 32'sd-0.14496956112410186, 32'sd0.1523195354207589, 32'sd0.14194729897115, 32'sd-0.09759798413660369, 32'sd-0.02954834089496485, 32'sd0.13253127540761547, 32'sd-0.047554506911188, 32'sd-0.04067497084866155, 32'sd-0.07198372413468118, 32'sd0.0876764237311551, 32'sd0.28436070018338666, 32'sd0.24189363560020952, 32'sd0.14409600962510533, 32'sd0.3715370000065665, 32'sd0.08835754274347855, 32'sd-0.13982219138344615, 32'sd-0.2657173489173034, 32'sd-0.23361107976815143, 32'sd0.034397019167875784, 32'sd0.05944505043746445, 32'sd0.054884473765441345, 32'sd-0.05464567602935361, 32'sd-0.19972925616826046, 32'sd0.12250329261764571, 32'sd-0.07413781111131368, 32'sd0.057634158555011215, 32'sd0.07025607304371642, 32'sd0.10060947250292449, 32'sd0.010958733588409108, 32'sd-0.05077027505381978, 32'sd0.12697736417040936, 32'sd-0.07148164051367212, 32'sd0.18462319803300267, 32'sd0.02417628446454927, 32'sd-0.23935492559987603, 32'sd0.1703958406058692, 32'sd0.11683115190495699, 32'sd-0.10068634169109687, 32'sd0.1478786805338412, 32'sd-0.05065516786650295, 32'sd-0.3010059220304603, 32'sd-0.09462060356431075, 32'sd0.09512550497693995, 32'sd0.2325968118631822, 32'sd0.2855169049882759, 32'sd0.1620188576922659, 32'sd-0.13477985003342652, 32'sd0.17807845613477147, 32'sd-0.00538649963398246, 32'sd0.018450547168919047, 32'sd0.017197813386365057, 32'sd-0.029078770380443694, 32'sd0.10678684579567499, 32'sd-0.11866032320518159, 32'sd-0.14573203069918972, 32'sd-0.2542466860077006, 32'sd0.11146577931949334, 32'sd-0.05882719744275309, 32'sd0.07813280720661128, 32'sd0.17405758224989687, 32'sd0.2511951508864771, 32'sd0.08577620616220052, 32'sd0.047616777251833664, 32'sd-0.0460376881433088, 32'sd-0.05013946442822148, 32'sd-0.24931590810485219, 32'sd0.04301176322625287, 32'sd0.07347315658799082, 32'sd-0.0015796554936328645, 32'sd-0.05169707102479825, 32'sd-0.10961308074511607, 32'sd-0.10554635297342081, 32'sd0.12586608307068411, 32'sd-0.026090454117849275, 32'sd-0.12329111043598921, 32'sd0.1977651666246206, 32'sd0.007243605864202731, 32'sd-0.03612150851255095, 32'sd-0.08132695885872339, 32'sd0.051761834404049904, 32'sd0.19191363900824684, 32'sd0.07980263343228379, 32'sd0.019527309573472307, 32'sd-0.09818002085484101, 32'sd-0.2011619611939584, 32'sd0.09720894399645694, 32'sd-0.03412555990618314, 32'sd0.183897920374837, 32'sd-0.18158362480000412, 32'sd-0.16062744530939185},
        '{32'sd0.04930627727635218, 32'sd-0.0162810523307647, 32'sd0.22118830405739875, 32'sd-0.0183210886692588, 32'sd-0.1264488604211499, 32'sd-0.060112201892443054, 32'sd0.12408039197466458, 32'sd-0.050372195602745584, 32'sd-0.15337571082185691, 32'sd0.1490885751833704, 32'sd0.12233573612024967, 32'sd0.23809990668845177, 32'sd0.19272321522081112, 32'sd-0.21572835578985966, 32'sd-0.034826784156669864, 32'sd-0.009879153378034109, 32'sd-0.3860119785784381, 32'sd0.0171524368166602, 32'sd0.0712323114088579, 32'sd-0.08738247291881032, 32'sd-0.2560718585001552, 32'sd-0.08956042892453032, 32'sd-0.017698806727925998, 32'sd0.005082076224633119, 32'sd0.133011609047143, 32'sd0.2758760206695822, 32'sd-0.010204171911248236, 32'sd0.11399826282034521, 32'sd0.11130450957320895, 32'sd-0.08027785235512465, 32'sd-0.06445759310240322, 32'sd0.15055179526658907, 32'sd0.12471285928103565, 32'sd-0.10756926350681187, 32'sd-0.08030839431385146, 32'sd0.038616079400611424, 32'sd0.014046717773948168, 32'sd0.1863195700861848, 32'sd-0.04816556412114351, 32'sd0.08365008206948377, 32'sd0.23000047149704028, 32'sd0.18828424918163952, 32'sd-0.25181355655067644, 32'sd-0.032311168327299154, 32'sd-0.18756025244892477, 32'sd0.03529084215690848, 32'sd-0.04847242217095089, 32'sd0.1485202060145715, 32'sd0.032415334010370556, 32'sd0.10116853826863254, 32'sd0.07880522186312804, 32'sd0.13873771119692693, 32'sd0.2156102810633606, 32'sd-0.08779834788086896, 32'sd-0.16424676565425114, 32'sd0.1108955922692109, 32'sd-0.024758917643914212, 32'sd0.09031388663689703, 32'sd-0.09507566209493834, 32'sd0.04009589380122175, 32'sd-0.011111120214362056, 32'sd-0.20336982909691712, 32'sd-0.2576737147121182, 32'sd-0.173296186111565, 32'sd0.135360927024912, 32'sd0.29591342217149114, 32'sd0.003715472837116173, 32'sd0.019780143455082708, 32'sd0.08262982795842269, 32'sd0.013750867743259976, 32'sd-0.16027565966444177, 32'sd0.00545063889774374, 32'sd-0.17160552871335258, 32'sd-0.06865791028838691, 32'sd0.04314714784539009, 32'sd0.22364005364650952, 32'sd-0.017675208695571827, 32'sd-0.18328202504497842, 32'sd-0.08478335907461661, 32'sd-0.09784950329856443, 32'sd-0.00024299212438487494, 32'sd0.12501193075870862, 32'sd-0.011148296562454375, 32'sd-0.14384090793681778, 32'sd0.13213962303921029, 32'sd0.12394832885850908, 32'sd-0.0035300977634893736, 32'sd-0.03484287022882493, 32'sd-0.0601117232139244, 32'sd0.15479285182437583, 32'sd0.015549729404730792, 32'sd-0.15633530513929234, 32'sd0.17141653241745966, 32'sd0.13296454395406115, 32'sd-0.15932031717566245, 32'sd0.3353533203244553, 32'sd0.28119196732563606, 32'sd-0.014054775636857813, 32'sd-0.06994331558290065, 32'sd0.09894644250413748, 32'sd-0.10332216982500281, 32'sd-0.08439697085556458, 32'sd0.07725742239597207, 32'sd-0.13745410589616533, 32'sd-0.07191351702233952, 32'sd-0.007576931899961624, 32'sd-0.14714160183950037, 32'sd-0.08061837954363964, 32'sd0.01035066251618813, 32'sd-0.06836843423961561, 32'sd-0.16975689815147113, 32'sd0.05804266003777638, 32'sd-0.23512993710143804, 32'sd0.07534976958194597, 32'sd0.16903044098779954, 32'sd-0.15814342684484173, 32'sd-0.15374440203545384, 32'sd-0.09049847713777194, 32'sd0.19742596930439174, 32'sd-0.015139557083108832, 32'sd0.21707585934212206, 32'sd0.08656340719381028, 32'sd-0.05704472598853245, 32'sd0.048785889748446956, 32'sd-0.24009892208921618, 32'sd0.0016983138077593472, 32'sd0.1093828943548637, 32'sd-0.08157858641987659},
        '{32'sd0.1124373716575407, 32'sd-0.08965583883691124, 32'sd0.20161822921288897, 32'sd0.17788529701582018, 32'sd0.10189092073593768, 32'sd-0.11487776707693911, 32'sd0.08580200889777312, 32'sd-0.09637267693039639, 32'sd-0.015782798246089434, 32'sd0.10341476236701755, 32'sd0.12424747264268358, 32'sd-0.12204011511279475, 32'sd0.19348835830033015, 32'sd0.12363366908525972, 32'sd-0.1633452985304775, 32'sd-0.11842571707622034, 32'sd-0.13442128755460017, 32'sd0.14626650981805966, 32'sd0.13889421985171937, 32'sd0.234128283517152, 32'sd0.058575780050669074, 32'sd0.033624302030074125, 32'sd0.1491040964609872, 32'sd0.19530287971254343, 32'sd0.02394431305447588, 32'sd-0.13359982202175313, 32'sd0.1393716747288832, 32'sd0.23857419794245155, 32'sd-0.1547217225092291, 32'sd-0.166841439057806, 32'sd-0.14511419965579303, 32'sd0.23461874367189767, 32'sd-0.13416336014535135, 32'sd-0.1229599222945017, 32'sd-0.14490740879011413, 32'sd-0.04024491854002757, 32'sd0.030713407205280725, 32'sd-0.006807473949639694, 32'sd0.08361752399510315, 32'sd-0.13943821663950304, 32'sd-0.0542947001717494, 32'sd-0.2054930124251525, 32'sd-0.040668338770631036, 32'sd0.05356455433726287, 32'sd-0.1832963713261383, 32'sd-0.284468158122977, 32'sd-0.10785097696467341, 32'sd-0.08641894957695684, 32'sd0.07440021575362588, 32'sd0.2315414967727155, 32'sd-0.2972194581668149, 32'sd0.12339808199495353, 32'sd-0.027994091776148037, 32'sd-0.0375767198197632, 32'sd0.1600101684694033, 32'sd0.039030291070727884, 32'sd-0.06894395539040137, 32'sd-0.11655738730868564, 32'sd0.17291192131352476, 32'sd-0.11697481243440874, 32'sd-0.2525082223588659, 32'sd-0.11419796461116402, 32'sd-0.05392424881129817, 32'sd0.12941622789878585, 32'sd0.029926784909485755, 32'sd-0.04276336228788155, 32'sd-0.3289119694027408, 32'sd0.11101793580274016, 32'sd0.09836229980682476, 32'sd-0.17167228547350052, 32'sd0.11495965555440939, 32'sd0.16247950700538108, 32'sd-0.16840864381006312, 32'sd-0.13973478699662537, 32'sd-0.09208080005217872, 32'sd-0.10192767020662603, 32'sd-0.07108735660066162, 32'sd0.25860442950447726, 32'sd-0.13848716955757143, 32'sd-0.14972964332846814, 32'sd0.07844255720228947, 32'sd0.09298615640153705, 32'sd-0.21014220779040343, 32'sd-0.1767102516573198, 32'sd-0.2949762558283207, 32'sd0.19285295802783506, 32'sd0.14481720959257185, 32'sd-0.11316093595240337, 32'sd-0.13394945618125093, 32'sd0.21085389293059126, 32'sd0.22466036492394795, 32'sd-0.1777504040226612, 32'sd-0.004401361165652655, 32'sd0.14012794307750334, 32'sd-0.0802423816603494, 32'sd-0.12468146863756402, 32'sd-0.09604790362410018, 32'sd0.11808642436311173, 32'sd0.1672936429034814, 32'sd0.07136813396417398, 32'sd-0.11664076061849726, 32'sd0.01585079136821368, 32'sd0.2755150541730441, 32'sd-0.17424481571697914, 32'sd-0.08150574645594992, 32'sd-0.0847445438610497, 32'sd-0.07658515385033926, 32'sd0.09790004657872858, 32'sd0.18341345883600557, 32'sd0.0349257094523004, 32'sd-0.21154073028952491, 32'sd0.01636611416389696, 32'sd0.23145544188830378, 32'sd-0.12391508982189609, 32'sd-0.09506022121720353, 32'sd0.11426189914680854, 32'sd-0.1305863248325061, 32'sd-0.04597180710946029, 32'sd-0.003631732418436946, 32'sd-0.06073037898080771, 32'sd0.0028418768133472065, 32'sd-0.11430618523101811, 32'sd0.00016638127390843047, 32'sd0.051157838752907026, 32'sd0.19490671463352077, 32'sd-0.022587950548351547, 32'sd0.05135518499623232, 32'sd0.029809473558635186},
        '{32'sd0.1707845876542315, 32'sd0.009457298938095153, 32'sd0.06984417134933409, 32'sd0.21782514991947302, 32'sd-0.18721274519205758, 32'sd-0.23553803039032, 32'sd-0.023778001215121365, 32'sd-0.04084150223377124, 32'sd-0.19029667877671302, 32'sd0.12576281302490816, 32'sd-0.21723386422879104, 32'sd-0.14979166615238243, 32'sd-0.15997969770170206, 32'sd0.060042910432501165, 32'sd-0.0644012028002236, 32'sd-0.07758654690272491, 32'sd-0.1880658587086508, 32'sd0.04386024614165655, 32'sd-0.15112675265041747, 32'sd0.0026419712315686474, 32'sd0.018232255880611628, 32'sd-0.10981688699737285, 32'sd0.08991728084094333, 32'sd0.13415857380185622, 32'sd-0.19067031559264375, 32'sd-0.1951424507354095, 32'sd0.010916729631101586, 32'sd-0.202988874420359, 32'sd-0.045116021830951876, 32'sd0.14968860709494713, 32'sd0.038168736017156056, 32'sd-0.03605960998083315, 32'sd-0.05458993339103582, 32'sd-0.18712289016483818, 32'sd0.05129446311128519, 32'sd0.021271617363636124, 32'sd-0.09049539028181004, 32'sd-0.1633193086718253, 32'sd0.0733175540580431, 32'sd0.179458613665316, 32'sd-0.13249671521896278, 32'sd0.17231085310864935, 32'sd0.055386420217945605, 32'sd0.10434182627032806, 32'sd-0.04101425525247009, 32'sd-0.12574513204915636, 32'sd-0.11546506691383127, 32'sd0.1578127501879702, 32'sd0.16669681372072132, 32'sd0.20408976021360858, 32'sd0.16334010071611177, 32'sd0.1063639527645538, 32'sd0.021348881261629576, 32'sd-0.03676835535127439, 32'sd0.0057708873930424264, 32'sd0.09791427284378613, 32'sd0.07150304905785829, 32'sd-0.02310744040587287, 32'sd-0.25701863983468504, 32'sd-0.1561150712867298, 32'sd-0.08714971343387096, 32'sd-0.14042958991209212, 32'sd0.08013729023541717, 32'sd0.11318037055916835, 32'sd-0.028089471175362105, 32'sd0.3154364102377048, 32'sd-0.26871264877824286, 32'sd-0.07176109217195398, 32'sd-0.18144803431483583, 32'sd0.25046316460422685, 32'sd-0.12682915938915376, 32'sd-0.29538212481874926, 32'sd-0.06626114815071137, 32'sd0.006146959383821005, 32'sd0.04201701918990299, 32'sd0.26321432431850406, 32'sd0.18493361887032883, 32'sd0.09764278679324559, 32'sd0.19295903942282655, 32'sd-0.20576862432018822, 32'sd-0.03851514147998322, 32'sd0.18786839567609623, 32'sd-0.03453651280587535, 32'sd-0.06961588637431046, 32'sd0.14525447479529444, 32'sd0.06304592056063878, 32'sd0.037484553289298894, 32'sd-0.21049563120928605, 32'sd0.021045917790587978, 32'sd0.2991218324233297, 32'sd-0.011784033630529945, 32'sd0.1879244046036959, 32'sd0.006255165328030147, 32'sd-0.04806850463365353, 32'sd0.15914343694468114, 32'sd0.13194919074103365, 32'sd-0.03726198223537601, 32'sd0.03201950907587747, 32'sd-0.3829754245674079, 32'sd-0.21868240196586491, 32'sd-0.04148636532138329, 32'sd0.22438772697810644, 32'sd0.05062891537312202, 32'sd0.1921236907939827, 32'sd0.01610054173356144, 32'sd-0.1661909201217459, 32'sd0.20483974540264627, 32'sd0.07236774513079215, 32'sd-0.2387427568779503, 32'sd-0.23495763360479932, 32'sd-0.15945978640950023, 32'sd0.10290699464356644, 32'sd0.041265706950195734, 32'sd0.12326132416171913, 32'sd-0.010813331319478345, 32'sd-0.09210056863996238, 32'sd0.02752431937960304, 32'sd0.18852747707633022, 32'sd0.18744397115907702, 32'sd-0.03446563302677721, 32'sd0.06033297290795496, 32'sd0.068542090560791, 32'sd0.19724540342076738, 32'sd-0.0007176767488267533, 32'sd-0.24351236458206615, 32'sd-0.07698205226267162, 32'sd0.11303148963810354, 32'sd-0.18035721924517756},
        '{32'sd0.20704656357893284, 32'sd0.23383887037924864, 32'sd0.055142047416895976, 32'sd-0.15466906522027604, 32'sd-0.08814592645903448, 32'sd0.2307707359838878, 32'sd0.1874486429284825, 32'sd0.06125770692722799, 32'sd0.14158543298272896, 32'sd-0.04762227503415046, 32'sd0.08463225908167028, 32'sd0.0547280159797368, 32'sd0.1911912336994564, 32'sd0.11537988370934191, 32'sd-0.12532567443752735, 32'sd0.20712182983244565, 32'sd-0.00022352437430890316, 32'sd-0.24283143386008613, 32'sd-0.07138344669713666, 32'sd-0.13483047305003001, 32'sd-0.1791868301946381, 32'sd0.23982238162779496, 32'sd-0.09717004065299208, 32'sd-0.22151490013390668, 32'sd-0.10683155772976022, 32'sd-0.05411066227650934, 32'sd-0.05758959317821833, 32'sd-0.1347393554979241, 32'sd-0.017073408123221195, 32'sd0.09957020943471591, 32'sd0.1477001577367542, 32'sd0.18665120589903172, 32'sd-0.05713944791276128, 32'sd0.024510989116381048, 32'sd0.06223269528115148, 32'sd0.1555379048518935, 32'sd-0.04614228271201671, 32'sd0.14946532328995715, 32'sd0.1532001645447463, 32'sd0.036212457782577034, 32'sd-0.018810225145393152, 32'sd0.029854325104997068, 32'sd0.17745107554979453, 32'sd0.11279828318277538, 32'sd0.11655034269189977, 32'sd-0.009629261779657826, 32'sd-0.14551141757948927, 32'sd0.13185183800702913, 32'sd0.05285179687462755, 32'sd0.1505685877253394, 32'sd-0.12297609087943769, 32'sd0.0812294975796686, 32'sd-0.07487324070260128, 32'sd0.18605845580097677, 32'sd-0.048237948707223255, 32'sd0.14598370866143542, 32'sd0.14038660894572205, 32'sd0.13510387651921288, 32'sd0.12269884136474497, 32'sd0.011841577093375369, 32'sd0.024319548725700635, 32'sd0.1822669206379864, 32'sd-0.12023226367691735, 32'sd0.15520543935924852, 32'sd-0.12487829071365592, 32'sd0.22094385830878946, 32'sd0.2996755733356412, 32'sd-0.1294358275015372, 32'sd0.06539364279608686, 32'sd-0.051214994456109275, 32'sd-0.07874111972877364, 32'sd-0.2705054089371138, 32'sd-0.02994381465641963, 32'sd-0.09364738060937526, 32'sd-0.07745128691079471, 32'sd0.1685284118860415, 32'sd-0.01626029031002801, 32'sd-0.1254888144608041, 32'sd0.08497033191661049, 32'sd0.024871188637496353, 32'sd-0.2018591940892871, 32'sd0.16385495707483955, 32'sd-0.09733502409983003, 32'sd0.07493766062171983, 32'sd-0.17469997247588906, 32'sd0.08814409310491583, 32'sd-0.3432602018221063, 32'sd-0.164488695150312, 32'sd-0.13238989197694076, 32'sd0.025655130115569618, 32'sd-0.21076166569469848, 32'sd-0.15512105376061897, 32'sd0.18034511607507575, 32'sd0.15551425790111195, 32'sd-0.04641221170204031, 32'sd0.21036572025040579, 32'sd-0.020954331084996253, 32'sd-0.007388373100180231, 32'sd-0.07061591935342677, 32'sd0.23237016976163402, 32'sd-0.06712554770932139, 32'sd-0.3196872127155091, 32'sd0.0029505287997528707, 32'sd0.023447062610615663, 32'sd0.0596624622335622, 32'sd0.19567673912611336, 32'sd-0.1299597080530256, 32'sd-0.08512302529563508, 32'sd-0.13371383879000473, 32'sd0.16109308259346422, 32'sd-0.002033021349338201, 32'sd-0.09552215924534518, 32'sd-0.16505446599280274, 32'sd-0.01354787635846547, 32'sd0.09067519258512721, 32'sd-0.18797610674506554, 32'sd-0.15659705339017332, 32'sd-0.19225273663201287, 32'sd-0.003144135499816484, 32'sd-0.03801249614501104, 32'sd0.19322151450311065, 32'sd0.11090032301031807, 32'sd0.016894488221231466, 32'sd-0.05581940700576331, 32'sd-0.006181773411102658, 32'sd-0.09469096819943755, 32'sd0.09176482600511732, 32'sd-0.13951864985529486},
        '{32'sd0.27441196768701287, 32'sd0.18901933988820976, 32'sd-0.04153087853185044, 32'sd-0.14983153297290994, 32'sd-0.18786467212477867, 32'sd0.04742320616833266, 32'sd0.27551054350228993, 32'sd-0.1080740742829519, 32'sd0.15063875663851772, 32'sd-0.07291618352736144, 32'sd0.19024122460773524, 32'sd0.02083707195884844, 32'sd-0.062089878345009286, 32'sd0.0910852208292761, 32'sd0.02636726811159371, 32'sd0.22883057946868973, 32'sd-0.08542248807138621, 32'sd-0.002551110944645974, 32'sd0.19910755314232131, 32'sd0.27036478999465535, 32'sd0.22504912906879151, 32'sd-0.12251341970507516, 32'sd0.19808203654443332, 32'sd0.06519489151975401, 32'sd-0.0016658718679486582, 32'sd-0.10561535171708343, 32'sd0.07409574572100662, 32'sd-0.06751001519397218, 32'sd-0.0904864000586876, 32'sd-0.1716659105252961, 32'sd-0.1107352802484748, 32'sd0.06954377139543949, 32'sd-0.06768177661120839, 32'sd-0.022882149163543045, 32'sd0.13309643521742945, 32'sd-0.08587248251384405, 32'sd-0.011914455260094596, 32'sd0.13172920863212081, 32'sd0.09151938013871957, 32'sd0.31087658524647505, 32'sd-0.14356419851456542, 32'sd-0.02633032169391683, 32'sd0.19316562893123515, 32'sd0.2202456547205115, 32'sd-0.18591234930817133, 32'sd0.15973950230060116, 32'sd0.08837873238825578, 32'sd0.15202060220184505, 32'sd-0.14871398665954558, 32'sd0.28651402038414175, 32'sd-0.2699372665309732, 32'sd-0.0640256588977805, 32'sd0.02815156144170802, 32'sd0.1833257500510615, 32'sd0.10213722712561972, 32'sd0.14257426454294106, 32'sd-0.1328352376676887, 32'sd-0.1136200094863475, 32'sd-0.034575182916908094, 32'sd0.08485432535827835, 32'sd-0.020004524482331112, 32'sd0.03739265513804528, 32'sd-0.08007285410094132, 32'sd0.04899138997381764, 32'sd0.1745605141884818, 32'sd0.12742039976458774, 32'sd-0.005055582709016114, 32'sd0.06379193882347764, 32'sd-0.14264928546032254, 32'sd0.011775469353423449, 32'sd-0.06929349561562982, 32'sd-0.07407639230141183, 32'sd0.12410404392125095, 32'sd-0.25149201053779346, 32'sd0.06443522305975699, 32'sd-0.017162565932962563, 32'sd0.20841270893698047, 32'sd-0.051501882663126546, 32'sd-0.11807304316072054, 32'sd0.04378779684326132, 32'sd0.012839168612847125, 32'sd0.2151625597910381, 32'sd-0.15287843686973504, 32'sd-0.04181925397473394, 32'sd-0.25025231777613255, 32'sd-0.1221212258177606, 32'sd0.033540577117628305, 32'sd-0.1688785338772455, 32'sd0.0030276691453271914, 32'sd-0.1315863372755496, 32'sd0.22769214463717594, 32'sd-0.16805501716882312, 32'sd0.18525837691638855, 32'sd-0.10711338285184971, 32'sd0.2886281079475856, 32'sd-0.2105115726334078, 32'sd-0.09506618625878567, 32'sd-0.06186312077834888, 32'sd0.11506742863091957, 32'sd0.10905504458262935, 32'sd0.23804072905341048, 32'sd0.06867999501232316, 32'sd-0.06718832508441737, 32'sd-0.05413030132044248, 32'sd0.13359004691986734, 32'sd-0.021553774213187674, 32'sd-0.03094120056116913, 32'sd0.041839320564826255, 32'sd-0.2943209092923158, 32'sd0.26728211822554615, 32'sd-0.07539419160591324, 32'sd-0.10062006121202281, 32'sd-0.16041028829794102, 32'sd-0.09557205751587368, 32'sd0.10459978007210176, 32'sd0.20680320646681388, 32'sd-0.07630122711481652, 32'sd0.11086144305851148, 32'sd-0.07172047176888548, 32'sd0.10235704616884665, 32'sd-0.2176024479280612, 32'sd-0.1033350718597839, 32'sd-0.3456120039226723, 32'sd0.16103239959655938, 32'sd0.17710275479176185, 32'sd-0.1255460185716462, 32'sd-0.1407575733150028, 32'sd0.005634205872129856},
        '{32'sd0.04479703978100399, 32'sd-0.18165731346131156, 32'sd-0.10839857883297001, 32'sd0.030437368372364406, 32'sd-0.192167744931782, 32'sd-0.18429941387362525, 32'sd-0.026346970334206788, 32'sd-0.14260804128288596, 32'sd0.039294363304972026, 32'sd0.14973010482585147, 32'sd0.04115189608504015, 32'sd-0.16214840113959225, 32'sd0.14757585392135877, 32'sd-0.015304322727343365, 32'sd-0.17778164140128, 32'sd-0.1498959181745771, 32'sd-0.00277022361281027, 32'sd-0.042670233235227735, 32'sd0.07715371969673582, 32'sd-0.08040336285114208, 32'sd-0.1795573233624698, 32'sd-0.08464416242120187, 32'sd-0.15693416286985548, 32'sd0.0188328104778218, 32'sd-0.0669253217053369, 32'sd0.12620837029282064, 32'sd-0.15697485499718591, 32'sd-0.11051526142140228, 32'sd-0.03876221380963746, 32'sd-0.20545424079661564, 32'sd-0.26232819460796447, 32'sd-0.11622854285291499, 32'sd-0.17692514195499134, 32'sd0.08998057854884886, 32'sd0.08870703335309998, 32'sd0.14336368339491726, 32'sd0.01860823209965293, 32'sd0.07495801009608963, 32'sd0.08365794711466334, 32'sd0.09011642518462479, 32'sd0.06587698425399267, 32'sd0.08330119233871915, 32'sd-0.28167310429669157, 32'sd-0.10651082173472613, 32'sd-0.15646228777427781, 32'sd0.04108369462504129, 32'sd0.037776572190894954, 32'sd-0.09737376781329386, 32'sd-0.06972842606378607, 32'sd-0.01258733184165488, 32'sd-0.07079144502677688, 32'sd-0.20275797013532254, 32'sd0.16218944803453636, 32'sd0.0647662636557683, 32'sd-0.1422042243537877, 32'sd0.1335901320564553, 32'sd-0.12841390217356266, 32'sd0.12986631937140847, 32'sd-0.10802894346302917, 32'sd0.17771299762916515, 32'sd0.018813023460133665, 32'sd0.14236426004569389, 32'sd0.18575881805466252, 32'sd0.12359348307925408, 32'sd-0.22671951348540562, 32'sd-0.13127038190831727, 32'sd0.16592318767423533, 32'sd0.25294949029907676, 32'sd-0.15025367511431317, 32'sd-0.19707478153091004, 32'sd0.15380188315891619, 32'sd-0.13870818784360858, 32'sd-0.18511810745365298, 32'sd-0.261674381893497, 32'sd-0.15159219690607972, 32'sd0.12012950436945188, 32'sd0.06371474491255885, 32'sd0.1217808678120736, 32'sd-0.15273992492551494, 32'sd0.059042822707969816, 32'sd-0.08720780629915352, 32'sd0.042104743199338594, 32'sd0.03785268374223804, 32'sd0.1333082548899647, 32'sd0.03953116279987161, 32'sd0.039944938038520277, 32'sd0.05343883957675769, 32'sd0.1757604719457457, 32'sd0.06682524132504256, 32'sd-0.3247358903737031, 32'sd-0.18090408997712226, 32'sd0.08665394418817643, 32'sd-0.04972647845012825, 32'sd-0.18401603654003298, 32'sd-0.1423911173936297, 32'sd0.004466012478848466, 32'sd0.15794181388872092, 32'sd-0.1730626885460903, 32'sd-0.03144727135197693, 32'sd-0.0036966900582920915, 32'sd-0.18866167729867486, 32'sd0.2651556000490465, 32'sd0.06878330456959436, 32'sd0.23377242589621725, 32'sd-0.030685973669659677, 32'sd0.21738346355325158, 32'sd0.022611901317313592, 32'sd0.12582766837700082, 32'sd-0.07041211278839832, 32'sd0.20452342729833264, 32'sd0.04950146134178328, 32'sd0.08057255883778332, 32'sd-0.03910948188286045, 32'sd0.2592178325353151, 32'sd-0.053150286200789966, 32'sd-0.14647672527327815, 32'sd0.23594066667859848, 32'sd-0.1625099836936615, 32'sd0.2573668467847582, 32'sd-0.007854327300389418, 32'sd0.15639459318700147, 32'sd-0.12753325058377682, 32'sd-0.14471196313816007, 32'sd0.2001860801627695, 32'sd-0.04557217473965701, 32'sd0.085981377670328, 32'sd0.10847701253673299, 32'sd0.06775949337834583},
        '{32'sd-0.03634399866884172, 32'sd-0.01659451467993783, 32'sd-0.10377117464934714, 32'sd0.23384134107951407, 32'sd0.075041629459985, 32'sd-0.05001879054985769, 32'sd0.059544753445625744, 32'sd-0.17790606782938934, 32'sd0.04712629221772376, 32'sd-0.10992674863504934, 32'sd-0.16886115546174008, 32'sd-0.09496458332526343, 32'sd0.16020424438442404, 32'sd0.23078609422221186, 32'sd0.2637470707363152, 32'sd0.13327431232939146, 32'sd0.10711915861379634, 32'sd0.1255566460114549, 32'sd0.16616965748734433, 32'sd0.17244905527432727, 32'sd-0.11562189407449418, 32'sd0.14301507763234375, 32'sd-0.14068069434010352, 32'sd0.09589322066891369, 32'sd-0.2950642260571499, 32'sd-0.16076745447977867, 32'sd0.22647905606213697, 32'sd-0.14989362636083242, 32'sd-0.0796141689996489, 32'sd-0.11792573269337119, 32'sd0.0390215699865096, 32'sd0.0058339439624001364, 32'sd-0.024988129389665614, 32'sd0.19236681155619373, 32'sd0.23365819915585004, 32'sd0.13558809066503447, 32'sd0.16312547912303524, 32'sd-0.1263578234498345, 32'sd0.09543268309031634, 32'sd-0.1151375479707443, 32'sd0.06328635647746438, 32'sd0.21321386936006081, 32'sd0.11415925019512936, 32'sd-0.2822974922523229, 32'sd0.014527882969165278, 32'sd-0.17910858446067876, 32'sd-0.1128774563496717, 32'sd-0.11224394627444843, 32'sd-0.2079095495002772, 32'sd-0.06894726189301453, 32'sd-0.0421795306173492, 32'sd-0.0027370656701615034, 32'sd-0.15861788403458835, 32'sd0.06340907973130679, 32'sd-0.08778797303135451, 32'sd-0.06528588346836289, 32'sd-0.07602537511656936, 32'sd-0.08192870159704252, 32'sd0.058390246515190244, 32'sd0.1828710836008575, 32'sd0.13080397272082225, 32'sd0.04069393078352358, 32'sd0.15295627769104445, 32'sd-0.041098077376173034, 32'sd0.014900690742272215, 32'sd-0.17392386119964223, 32'sd0.05085913088368157, 32'sd0.2643835374168539, 32'sd-0.03523328520430831, 32'sd0.018856519949508842, 32'sd-0.12969350658659037, 32'sd0.05079394074185103, 32'sd-0.11606463952115162, 32'sd0.10000758961417004, 32'sd-0.04358675778494082, 32'sd-0.0687060737055748, 32'sd-0.18828501112461213, 32'sd-0.0804369480423773, 32'sd-0.05779994642751452, 32'sd0.14714715860128416, 32'sd0.11167955460128053, 32'sd-0.13381530625300117, 32'sd-0.07131430513913953, 32'sd0.17788747986062653, 32'sd-0.06548539941745113, 32'sd0.2252596689585564, 32'sd-0.10351241062582932, 32'sd-0.22511456984577422, 32'sd0.03982168316368124, 32'sd0.13038679548273513, 32'sd0.028990364814292915, 32'sd0.10717169952495352, 32'sd0.07984562845133397, 32'sd0.2210874822469563, 32'sd-0.09165620677140358, 32'sd-0.19970620938528472, 32'sd-0.2152037212439353, 32'sd0.030247521076813607, 32'sd-0.09563146198634956, 32'sd-0.22620342838149893, 32'sd-0.28773456753006854, 32'sd0.19085831467482356, 32'sd-0.14506553345538536, 32'sd0.12726538341251745, 32'sd-0.07903147645359583, 32'sd-0.032247217467948806, 32'sd-0.12060117035573154, 32'sd0.19405769794495864, 32'sd0.11081472662442741, 32'sd0.16762146074311346, 32'sd0.06880614766759835, 32'sd0.11044424459207053, 32'sd-0.055171284435125416, 32'sd-0.055729190819794314, 32'sd0.129224959423768, 32'sd-0.04084271752977519, 32'sd0.1043566393071485, 32'sd0.009679854677197331, 32'sd0.18370759234890266, 32'sd0.04168815283592808, 32'sd0.060738380056297496, 32'sd-0.09184593548843753, 32'sd0.15070127994597932, 32'sd-0.004022921685463369, 32'sd-0.04315813961648193, 32'sd-0.2553864558157467, 32'sd0.18239490641535425, 32'sd0.0016047283523625585},
        '{32'sd0.08865663691821672, 32'sd-0.21409649491039598, 32'sd-0.09786214686916062, 32'sd0.043836897196878985, 32'sd0.15151664141540777, 32'sd0.038604084083607854, 32'sd-0.16367270267720643, 32'sd-0.2224944133724347, 32'sd0.25988808979099615, 32'sd-0.12743009645678133, 32'sd0.22745262354794285, 32'sd0.2190873669942652, 32'sd0.05053898477435882, 32'sd0.2004567458312615, 32'sd0.0866090411778341, 32'sd-0.1956298138338499, 32'sd-0.18002667545153206, 32'sd0.09574009472969318, 32'sd-0.1048515315443082, 32'sd-0.16619550613814005, 32'sd-0.1184986773879043, 32'sd0.08647782656671692, 32'sd-0.1765614033219924, 32'sd0.12136986880503378, 32'sd-0.13060181838171134, 32'sd0.061222814807808223, 32'sd-0.27311714865572856, 32'sd-0.13094144541022235, 32'sd-0.07427709966860568, 32'sd-0.07915441924840075, 32'sd-0.2634355080051492, 32'sd0.08776743161760196, 32'sd0.08348770555726809, 32'sd-0.16818977127464504, 32'sd-0.05936238917523251, 32'sd-0.07219945449912661, 32'sd-0.21398229551854003, 32'sd0.16642671412678128, 32'sd-0.14406842945729936, 32'sd0.1238159257909169, 32'sd-0.08895631129495607, 32'sd0.00799725685730345, 32'sd-0.046830672160588886, 32'sd-0.03845468208060102, 32'sd-0.07663601130514049, 32'sd-0.17598693879526806, 32'sd-0.04109733371397508, 32'sd-0.20391522071291276, 32'sd-0.0435157031029633, 32'sd-0.2013132855780338, 32'sd0.19247431463456935, 32'sd0.035337153500294365, 32'sd-0.254768373045211, 32'sd0.12889641497932286, 32'sd-0.04575660216148887, 32'sd0.19689183954549608, 32'sd0.12211904623663968, 32'sd0.08886453557138407, 32'sd0.1958362903573727, 32'sd0.16236496997591768, 32'sd0.02175342843655618, 32'sd-0.13651758830711774, 32'sd-0.08653986946757711, 32'sd0.09564675952523992, 32'sd0.1120716042931062, 32'sd0.06926584148934692, 32'sd0.1926680794357959, 32'sd0.13422316055676684, 32'sd-0.2333294337550751, 32'sd-0.14876493162021884, 32'sd0.1782629189016151, 32'sd-0.04900937289582079, 32'sd0.21519064717995895, 32'sd0.04113476386380414, 32'sd0.1720731600045838, 32'sd-0.06590520625181887, 32'sd-0.20521489393203776, 32'sd0.15056587083314762, 32'sd0.1572780401449927, 32'sd0.20640234639980656, 32'sd-0.16193754172193445, 32'sd-0.08116845182825536, 32'sd-0.03884205526852025, 32'sd0.09047885854859503, 32'sd0.06213924147548526, 32'sd-0.1635305045676188, 32'sd0.0036179019822959145, 32'sd0.035049138444811424, 32'sd0.09952181486502071, 32'sd0.17737028123065404, 32'sd0.05028780976261, 32'sd-0.07639434980650839, 32'sd0.06895846342034552, 32'sd0.2578057093333824, 32'sd-0.14672139297488118, 32'sd0.22888716584393934, 32'sd-0.05733787623567155, 32'sd0.06728024062491568, 32'sd0.20640913470558656, 32'sd-0.16959080613686614, 32'sd0.1556251293261971, 32'sd-0.05956153616838975, 32'sd-0.19072914346718983, 32'sd-0.18509770369446546, 32'sd-0.21280722432198523, 32'sd0.11901805605221416, 32'sd0.005396805703964412, 32'sd-0.25757540780480304, 32'sd-0.09210971528071366, 32'sd0.09470977790458092, 32'sd-0.29204628039114017, 32'sd-0.1603754436667794, 32'sd-0.10821259023228032, 32'sd0.05910815695233198, 32'sd0.2301711074299455, 32'sd0.2465950759713846, 32'sd0.17058171879135747, 32'sd0.24698051065518747, 32'sd-0.12055068886611447, 32'sd-0.0038427637378415733, 32'sd0.23119010038162607, 32'sd0.0654900508469528, 32'sd-0.03269169541238802, 32'sd-0.015870791109908706, 32'sd-0.16270825724074947, 32'sd0.1079831494801094, 32'sd-0.2579055229589065, 32'sd0.15527863623134788},
        '{32'sd0.17742526874134187, 32'sd0.21144767508459586, 32'sd-0.12933445107060923, 32'sd0.08190099159688709, 32'sd0.07353045591628364, 32'sd0.15339732604605805, 32'sd-0.09508323400527756, 32'sd-0.18659367460295243, 32'sd0.0894134259066565, 32'sd-0.11843923644069809, 32'sd-0.02030083124405215, 32'sd-0.030190138036411452, 32'sd-0.1795706057698076, 32'sd-0.01268364073682013, 32'sd0.14314070425158187, 32'sd0.13764957126058316, 32'sd-0.10648614447233225, 32'sd0.10005396773612084, 32'sd0.06495043724286215, 32'sd0.033496516018611006, 32'sd-0.06976597466626248, 32'sd0.09270621414059739, 32'sd0.19956261525854543, 32'sd0.0765117005625103, 32'sd0.0021586720381291035, 32'sd0.1506103336862878, 32'sd0.09690891010051554, 32'sd-0.15561377458851428, 32'sd-0.01735333799684215, 32'sd-0.10948414449946077, 32'sd0.15335169491564055, 32'sd-0.025615576197388797, 32'sd-0.215921471511173, 32'sd0.008542427667225634, 32'sd-0.07516218966080145, 32'sd0.19024119106436543, 32'sd-0.15609881883376056, 32'sd-0.0493571843387178, 32'sd0.09207225273105031, 32'sd0.3200468952677558, 32'sd-0.10357649029302526, 32'sd-0.004121795628869522, 32'sd-0.06757283299589438, 32'sd-0.0669768380614784, 32'sd0.2990338082602594, 32'sd-0.003092052108960158, 32'sd0.05267373131199814, 32'sd0.16227200890285667, 32'sd-0.16623585408507122, 32'sd0.012356758390852873, 32'sd-0.2514078335638942, 32'sd0.013066244044145511, 32'sd0.18295323469721855, 32'sd0.1260339792128059, 32'sd-0.05454715229810053, 32'sd-0.1964680821472705, 32'sd-0.14204801027121763, 32'sd0.012939795214823352, 32'sd0.028658991992145253, 32'sd0.06841050016074549, 32'sd-0.1919368458650409, 32'sd-0.0004886646391829675, 32'sd0.0973822648747305, 32'sd-1.4826266863332061e-05, 32'sd0.04492822486470792, 32'sd-0.1546418314224339, 32'sd0.16185484739352504, 32'sd-0.25554483416296736, 32'sd0.13146236182872656, 32'sd-0.09702834888196965, 32'sd0.18119878028064088, 32'sd-0.010104965397526453, 32'sd-0.05652882393228828, 32'sd-0.06744432330345465, 32'sd0.016836904632322198, 32'sd0.0060116849188752205, 32'sd0.07599869170982039, 32'sd-0.09588775230948084, 32'sd-0.07836214317709816, 32'sd0.11791748405559013, 32'sd-0.14813038004036866, 32'sd-0.11108191346388403, 32'sd0.31711178801436735, 32'sd-0.04398318700399931, 32'sd-0.20008595417156053, 32'sd0.08915357718610718, 32'sd0.1582709477912594, 32'sd-0.09679776676525738, 32'sd0.0851230411090462, 32'sd0.15481810138634272, 32'sd-0.21601049138496167, 32'sd-0.23030325907201254, 32'sd0.06534186941943375, 32'sd0.1968862385870539, 32'sd-0.13522056925325748, 32'sd-0.11255983194122265, 32'sd0.03283702659570774, 32'sd0.007342500228033401, 32'sd-0.09915931694599814, 32'sd0.08856071936152725, 32'sd0.18780684404867895, 32'sd0.06551133203745568, 32'sd0.1433231068509163, 32'sd-0.20984440563885778, 32'sd0.15666693566645445, 32'sd0.09531484285817568, 32'sd-0.2165556515458485, 32'sd0.011628584810332023, 32'sd-0.2397613424382458, 32'sd0.2347543306053016, 32'sd-0.05828368527603044, 32'sd-0.017193739375735206, 32'sd-0.08644754336524958, 32'sd0.2472596229088162, 32'sd0.15904699310871742, 32'sd-0.17809593118078476, 32'sd-0.02077348750823937, 32'sd-0.10980185310149095, 32'sd0.14089257141416292, 32'sd0.18561464607877168, 32'sd-0.1973443785041712, 32'sd0.10291582345646381, 32'sd-0.15698488706714384, 32'sd-0.1892438336852554, 32'sd0.19565495035090424, 32'sd-0.17120333702050836, 32'sd0.05888676305864618, 32'sd0.009499491367882983},
        '{32'sd0.17087831616269286, 32'sd0.13421987483478942, 32'sd-0.15641987920033723, 32'sd-0.01774235582995582, 32'sd-0.22628889653049666, 32'sd0.2166920367479275, 32'sd0.05582355431398279, 32'sd0.2067412856525253, 32'sd0.10645241565291254, 32'sd-0.1453821455362384, 32'sd0.020652447399692086, 32'sd0.05720231997663302, 32'sd0.16603928955610137, 32'sd-0.02473428188755126, 32'sd-0.01989624907519309, 32'sd0.13861333497196182, 32'sd0.035306707090899545, 32'sd-0.1538500439350062, 32'sd-0.14086756665977154, 32'sd-0.2274306202468654, 32'sd-0.02702088837773562, 32'sd-0.044781038696651135, 32'sd-0.11734865023928241, 32'sd0.08267439327030686, 32'sd-0.26454479100784445, 32'sd-0.05052736341638224, 32'sd0.04193044642972785, 32'sd-0.1674444567631864, 32'sd-0.013192878927761529, 32'sd0.21713380128005003, 32'sd-0.20434555670448928, 32'sd0.07084684777519336, 32'sd0.07285865593509991, 32'sd0.05953200876911039, 32'sd-0.045427580475171266, 32'sd0.07103574075991466, 32'sd0.21859872662338214, 32'sd0.16815644124906678, 32'sd0.025389357932768763, 32'sd-0.172491590632691, 32'sd-0.12110071165449787, 32'sd0.07242727937225749, 32'sd0.16713861121399415, 32'sd-0.13868601918598225, 32'sd0.11294831506191114, 32'sd0.12341764284227254, 32'sd0.22942562377343473, 32'sd-0.18728582002095864, 32'sd0.04317543943180642, 32'sd0.18005119292667318, 32'sd0.19598821490205254, 32'sd-0.2728214537773017, 32'sd-0.12599119102587172, 32'sd-0.21050163835734548, 32'sd-0.08991314832037943, 32'sd-0.018846122434576038, 32'sd0.14158243181299884, 32'sd-0.03264528556125997, 32'sd-0.2751087959470973, 32'sd0.07845014576517777, 32'sd0.009573188989180071, 32'sd0.20084216859065782, 32'sd-0.010557580490140363, 32'sd0.268894293922562, 32'sd0.043576267594235045, 32'sd-0.05180626391602011, 32'sd-0.13286137649275773, 32'sd0.1373221378656134, 32'sd0.07204673404985414, 32'sd-0.17372231413541633, 32'sd-0.008819756883188472, 32'sd0.15024939661221878, 32'sd0.08866842438172967, 32'sd0.08414282967101044, 32'sd0.21062597797602373, 32'sd-0.17353290541011232, 32'sd0.03860964910094717, 32'sd0.12152442886200733, 32'sd0.13392833343467214, 32'sd-0.038722898471245874, 32'sd0.08395704954110117, 32'sd-0.05402949435242756, 32'sd-0.09932640924695281, 32'sd-0.19320798992599567, 32'sd-0.05282418405332343, 32'sd0.07812790223590924, 32'sd-0.14762964512668744, 32'sd-0.2060246635154726, 32'sd0.24971740759904495, 32'sd-0.024518934105597003, 32'sd-0.1050319704924548, 32'sd0.3004176101689115, 32'sd-0.2640470614740921, 32'sd0.311069253727997, 32'sd-0.15678347779657445, 32'sd0.1273006757738421, 32'sd-0.17935074016452432, 32'sd-0.19643346133912762, 32'sd-0.07229798882624695, 32'sd-0.1864541467867217, 32'sd-0.20039653431135618, 32'sd-0.14440439464749769, 32'sd0.043844938810589436, 32'sd-0.021219999118073797, 32'sd-0.1166840901077614, 32'sd0.03358947637855281, 32'sd-0.050781877541589526, 32'sd0.0775670492766821, 32'sd-0.15654028364953773, 32'sd0.2728992614729893, 32'sd0.06842846918660989, 32'sd0.092066938012969, 32'sd0.20717401996117155, 32'sd0.03804671270642592, 32'sd0.055438279138616, 32'sd0.14099368052647587, 32'sd-0.1445424726716564, 32'sd-0.1350503516611676, 32'sd0.09190002478847782, 32'sd0.18098947520205735, 32'sd0.04185432518526838, 32'sd0.08208351163434116, 32'sd-0.031794560801495425, 32'sd0.07944379558187196, 32'sd0.04443212277395301, 32'sd-0.17324909738959782, 32'sd0.09280278146322923, 32'sd0.20037750608427563},
        '{32'sd0.23016294709578147, 32'sd0.1725522966513939, 32'sd0.12734452337140056, 32'sd0.2499518236168741, 32'sd-0.10484369212886728, 32'sd-0.22954985910242315, 32'sd-0.1146322671187505, 32'sd-0.058364198029016684, 32'sd0.024933458134783093, 32'sd0.028896547258357896, 32'sd0.07573121231747704, 32'sd0.10405465318375508, 32'sd0.029960777913754358, 32'sd-0.10597080742498369, 32'sd0.03865941307306001, 32'sd-0.07125467239883929, 32'sd-0.1486982357635464, 32'sd-0.2184245635320736, 32'sd-0.043422107199191984, 32'sd-0.22241798443689811, 32'sd0.10918560701785353, 32'sd-0.012887594227281753, 32'sd-0.1936330584086619, 32'sd0.20265042698648697, 32'sd-0.06567976849891789, 32'sd0.1623126342140267, 32'sd-0.1283997045389111, 32'sd-0.3335294130536792, 32'sd-0.07437487195491264, 32'sd0.025948518128433462, 32'sd-0.22308241727849717, 32'sd0.1483242520278168, 32'sd0.16631424854693827, 32'sd-0.18390743868263892, 32'sd0.1132636060631204, 32'sd-0.20467886862294155, 32'sd-0.08139908876310971, 32'sd-0.04840367891709102, 32'sd0.06352214992430386, 32'sd-0.03068284526909977, 32'sd0.02018053044409045, 32'sd0.1624450665433696, 32'sd-0.16665484809950318, 32'sd-0.020333411346155777, 32'sd0.09371158597681274, 32'sd0.15848447429758597, 32'sd0.1778295844320063, 32'sd-0.03798635749848519, 32'sd0.017981476637671495, 32'sd-0.21571985149350403, 32'sd0.09845132573187695, 32'sd-0.26021259926804213, 32'sd0.1576617769870208, 32'sd-0.001046252190024784, 32'sd-0.16834884681875678, 32'sd-0.16750958204961405, 32'sd0.08505541675766064, 32'sd-0.07005723442461212, 32'sd0.10585429997528714, 32'sd-0.15428011297267233, 32'sd0.08254756578369607, 32'sd-0.026288146786488026, 32'sd0.03484572812252977, 32'sd0.05172673605768431, 32'sd0.060346111376816704, 32'sd0.09077992903571148, 32'sd0.03228323060931054, 32'sd0.11469062400462887, 32'sd0.010499138292978402, 32'sd0.18311086500213725, 32'sd0.0315435255810436, 32'sd-0.07878780110942614, 32'sd-0.031557038208377415, 32'sd-0.032677599636354485, 32'sd0.023614386176526305, 32'sd0.1996161306309547, 32'sd-0.029069302624684143, 32'sd0.31261391809764794, 32'sd0.12565654243106195, 32'sd-0.19603702162636463, 32'sd0.16958034017163476, 32'sd0.25231069376684956, 32'sd-0.15109956005398031, 32'sd-0.1682002839249846, 32'sd0.02841031835273748, 32'sd-0.14172057845443967, 32'sd0.12546123805873838, 32'sd0.05328546392585652, 32'sd0.173754260417429, 32'sd0.024456828405839157, 32'sd-0.10912796918993677, 32'sd0.24535977582149074, 32'sd-0.05890379161543273, 32'sd-0.10579681378556348, 32'sd0.11899459308932259, 32'sd-0.0801897022177889, 32'sd-0.14089062682512754, 32'sd0.022105487567868783, 32'sd-0.12985243796660348, 32'sd-0.06018482800775345, 32'sd0.12840779637988986, 32'sd0.02112141194109116, 32'sd0.29966248819289126, 32'sd0.19006794743591635, 32'sd0.11256219258192415, 32'sd0.16054333689881772, 32'sd0.029796172278211217, 32'sd-0.13270827417659853, 32'sd-0.20771358286573635, 32'sd0.1958781193894345, 32'sd0.20675187047826005, 32'sd-0.15625610791627267, 32'sd-0.0507968228040756, 32'sd0.12238264893880262, 32'sd0.10209243747246163, 32'sd0.15311857349388697, 32'sd-0.188532540606382, 32'sd-0.01124000493498724, 32'sd0.15575410784252935, 32'sd0.09551986898454123, 32'sd0.1261844051511057, 32'sd0.06563269063050405, 32'sd-0.2181055101623067, 32'sd0.05675125852884597, 32'sd0.006770359705951636, 32'sd0.021937806902314897, 32'sd-0.09971079056812027, 32'sd-0.06543649299232544},
        '{32'sd-0.2449870022723994, 32'sd0.08563403311349398, 32'sd0.14194420763598178, 32'sd0.20899393173379097, 32'sd-0.22128439428246807, 32'sd0.13521610393116662, 32'sd0.16438797967270036, 32'sd0.10981744569006188, 32'sd-0.2468665197447044, 32'sd0.07562181892851547, 32'sd-0.08039187066517085, 32'sd-0.014550283867100408, 32'sd0.18194601875021127, 32'sd0.05073013596836702, 32'sd-0.042330666193550935, 32'sd0.2372931950542768, 32'sd-0.017685591257882268, 32'sd-0.1513511972549094, 32'sd0.0707703323794637, 32'sd-0.2989578274925079, 32'sd-0.13132679545234666, 32'sd0.2081311460288318, 32'sd-0.09895042071624818, 32'sd0.026497760617440972, 32'sd-0.01722699017439275, 32'sd-0.15082383735989566, 32'sd0.10759126769176185, 32'sd-0.07862880242115361, 32'sd-0.010177970277447417, 32'sd0.056058600363107954, 32'sd-0.14172382534929176, 32'sd0.1973334678594927, 32'sd0.023502088422235702, 32'sd-0.1458851892925414, 32'sd0.08973745165479785, 32'sd0.23407195712331613, 32'sd-0.05127264608806441, 32'sd0.18449097883082707, 32'sd0.06441890487882342, 32'sd-0.1409358898189393, 32'sd0.008571898316971225, 32'sd0.011871685804914274, 32'sd0.17417633191210777, 32'sd0.09775005850878082, 32'sd-0.24776446762785592, 32'sd0.06575555534784662, 32'sd0.06944066799483178, 32'sd-0.04436463849355884, 32'sd0.04279318341484799, 32'sd0.044884199576684845, 32'sd-0.0453013631438247, 32'sd-0.02178336812042685, 32'sd0.1069125162100456, 32'sd-0.06086329311133553, 32'sd-0.2666353834450941, 32'sd0.0179991912800561, 32'sd0.19835177833371648, 32'sd0.21824789117907448, 32'sd-0.16975672260655886, 32'sd-0.060294328133392444, 32'sd0.06692828547985918, 32'sd0.014181730073500194, 32'sd-0.15938556509201957, 32'sd-0.012593937049892647, 32'sd-0.05864113001445474, 32'sd0.18303990120304708, 32'sd-0.0487455162950437, 32'sd-0.06544489524312823, 32'sd-0.11196187701149365, 32'sd0.09384857958844067, 32'sd0.17045441118749793, 32'sd0.03163472942390505, 32'sd-0.08500256318663718, 32'sd-0.15330885996911545, 32'sd-0.015307840912515865, 32'sd0.08682259153569946, 32'sd0.1102516018775524, 32'sd0.1827396334879431, 32'sd-0.1957992042830822, 32'sd-0.09586079007903744, 32'sd-0.17996704334870114, 32'sd0.005679321453226243, 32'sd0.1633746197626654, 32'sd-0.0259664970252552, 32'sd0.07574558347473412, 32'sd0.18635142192862658, 32'sd-0.04837761979294687, 32'sd0.12293701423772119, 32'sd0.11589387075539265, 32'sd-0.15609965150954266, 32'sd0.06116963937554861, 32'sd-0.09951050586249996, 32'sd0.05502365620065216, 32'sd0.051528542268347494, 32'sd-0.15929290471762086, 32'sd0.0950612093751319, 32'sd0.06652555786455863, 32'sd0.04803293917968261, 32'sd-0.008406958893623752, 32'sd-0.1290022700127286, 32'sd0.13727890103478274, 32'sd0.11904141169219698, 32'sd0.15728885628820644, 32'sd0.14968929100012324, 32'sd-0.17622228038437998, 32'sd0.02109839556915034, 32'sd0.16094103239283802, 32'sd0.015412860579054482, 32'sd-0.16087964436892152, 32'sd-0.0804090883090474, 32'sd0.1745902438684875, 32'sd0.07068383321198674, 32'sd-0.2695957496994674, 32'sd0.34470518522190097, 32'sd0.11248132620468518, 32'sd-0.1284544970313136, 32'sd-0.10741256443370152, 32'sd-0.04138947545460984, 32'sd0.10096116157821719, 32'sd-0.1472656835439975, 32'sd0.15853568388777775, 32'sd0.004104763649111407, 32'sd-0.07290361803404903, 32'sd0.06840180532034032, 32'sd0.09140059345027855, 32'sd0.06685814381301294, 32'sd-0.12392274840037341, 32'sd-0.012470234804287715},
        '{32'sd0.014109771689433245, 32'sd0.16402890121687555, 32'sd0.10180156079719242, 32'sd-0.21747126749327816, 32'sd-0.042262479780604434, 32'sd0.12167514739967825, 32'sd-0.32112301211849603, 32'sd-0.02561101519095785, 32'sd0.22385296399387358, 32'sd-0.21627091446368224, 32'sd0.2311725135520952, 32'sd0.02699334359450985, 32'sd-0.15672005297972977, 32'sd0.10614147737847317, 32'sd0.13307201151679568, 32'sd-0.03288976944567041, 32'sd0.15901069286562972, 32'sd0.06391552657110836, 32'sd0.021080754285590503, 32'sd-0.11239658604507798, 32'sd0.033506923473298235, 32'sd0.030855622564037385, 32'sd0.25777780489616997, 32'sd0.13492648148253153, 32'sd-0.15075046551394577, 32'sd-0.023269741402238465, 32'sd-0.15418170561807668, 32'sd-0.06935119251938371, 32'sd-0.01766203955413607, 32'sd0.1885628417237425, 32'sd0.08032897065457514, 32'sd0.1033243327783656, 32'sd-0.1634577017546302, 32'sd0.11457203265792558, 32'sd-0.1814514775127235, 32'sd0.0687012572720078, 32'sd-0.21175450294691023, 32'sd-0.1422679249046747, 32'sd-0.10534703163957773, 32'sd0.14228446183328625, 32'sd-0.0809707418370771, 32'sd0.01469818002196955, 32'sd0.08284093976006882, 32'sd0.16334670571280638, 32'sd-0.20362847680214993, 32'sd0.061160056370395545, 32'sd-0.1912977794104771, 32'sd-0.027097732524889447, 32'sd-0.1689217547600314, 32'sd0.1564117787899061, 32'sd-0.054301926119068325, 32'sd0.10506129175544514, 32'sd-0.060653515654971124, 32'sd-0.05844562330849364, 32'sd0.07716014476060412, 32'sd0.1468553685428662, 32'sd-0.1767776897582758, 32'sd0.051684161188363005, 32'sd-0.17605393789577442, 32'sd0.12153383127259659, 32'sd-0.014034891312160801, 32'sd0.020652063622932294, 32'sd-0.04832746173499599, 32'sd0.17299578502856658, 32'sd0.0414759206581334, 32'sd-0.028252778650652483, 32'sd-0.08292140183600909, 32'sd-0.1169636089416623, 32'sd-0.1973300841130684, 32'sd-0.14184318541202368, 32'sd-0.1747163213333434, 32'sd-0.08272896810202518, 32'sd0.14075973096653574, 32'sd-0.14691496867718362, 32'sd0.2500002532620269, 32'sd-0.14665047837656395, 32'sd-0.058919486471954705, 32'sd0.035278201766675364, 32'sd0.08386663705443491, 32'sd0.0609827218049992, 32'sd0.15560882683876998, 32'sd-0.15056900366144224, 32'sd-0.0261385823247607, 32'sd0.044615320747348974, 32'sd0.0025276486609926863, 32'sd-0.02046171326335954, 32'sd-0.17559858297993927, 32'sd-0.024019422141517505, 32'sd-0.032740087504891935, 32'sd0.1804781071194742, 32'sd0.06786005809965708, 32'sd0.032722284688265456, 32'sd0.11127166813184317, 32'sd0.12913792570271376, 32'sd0.12886813172151285, 32'sd0.16233031350100494, 32'sd0.03498679292539721, 32'sd0.16201001778050986, 32'sd0.05654293837747564, 32'sd-0.055588626594799066, 32'sd-0.1389783427085918, 32'sd-0.15708686807245426, 32'sd-0.22360976575775696, 32'sd0.01575925092562057, 32'sd-0.13645543083754041, 32'sd-0.22209550176472062, 32'sd0.09571551167729395, 32'sd0.14553716727385663, 32'sd0.060835225684182925, 32'sd-0.06914496413305797, 32'sd-0.15135126566515375, 32'sd-0.10664760786055424, 32'sd0.2530741922667916, 32'sd-0.22061270835426336, 32'sd0.09555384601505604, 32'sd-0.056114580263698755, 32'sd0.11368375835960531, 32'sd0.05548090130751529, 32'sd-0.06182644479494501, 32'sd-0.22913913034225064, 32'sd0.14422646497012026, 32'sd0.05277153282738927, 32'sd0.18547877336089783, 32'sd-0.19919661896303179, 32'sd0.13904058407474654, 32'sd0.12984153421315514, 32'sd-0.1384805248069023, 32'sd0.24369069748057584},
        '{32'sd-0.2793604784829152, 32'sd0.18477771091592168, 32'sd-0.1164261983929463, 32'sd-0.23243144624533693, 32'sd-0.03184349822842852, 32'sd-0.030999212766479413, 32'sd0.11021715855456678, 32'sd0.1557583540811971, 32'sd-0.18087673166769166, 32'sd0.06951513090317571, 32'sd-0.07476642070536788, 32'sd-0.14952988196747619, 32'sd0.01004511897647611, 32'sd0.2177482516589916, 32'sd0.06840488700837766, 32'sd0.20430431757559664, 32'sd-0.0901629555791742, 32'sd0.054400767385028304, 32'sd0.07683137871277602, 32'sd-0.09303172287200834, 32'sd0.029673379659610147, 32'sd0.02924420692243451, 32'sd0.07766648089092715, 32'sd0.11795015076553662, 32'sd0.2166443722927861, 32'sd0.14788512914505622, 32'sd0.023095768140254425, 32'sd0.2253968919734878, 32'sd0.11295085611511535, 32'sd0.10430521971624353, 32'sd-0.021160724449313714, 32'sd-0.2014649799010926, 32'sd-0.17605081117390117, 32'sd-0.04374207008950783, 32'sd-0.05253968673639697, 32'sd-0.1624654685962775, 32'sd-0.2280905537672809, 32'sd-0.0706103905117005, 32'sd-0.23417923647606426, 32'sd-0.17478270965117818, 32'sd-0.06442424544031498, 32'sd0.0007053583906935941, 32'sd0.007752439283951759, 32'sd0.037544529298641494, 32'sd-0.13410467941329943, 32'sd-0.0031465360667117317, 32'sd0.15988976999658933, 32'sd-0.0233737450376205, 32'sd-0.08377409549687564, 32'sd0.1099086648977188, 32'sd0.13191928556585228, 32'sd0.14616609514961595, 32'sd0.012309724020709865, 32'sd0.05665720923972392, 32'sd0.10050643095579911, 32'sd0.1728373500274745, 32'sd-0.10286348771039622, 32'sd0.08906992991084788, 32'sd0.34016419504655016, 32'sd-0.005092416854662629, 32'sd-0.015928274430383027, 32'sd0.15594936899261863, 32'sd-0.07818822964299765, 32'sd0.1348638535592858, 32'sd0.12690056759071694, 32'sd0.06958662746628268, 32'sd-0.10307760023346998, 32'sd0.126684763901773, 32'sd-0.14878065237941926, 32'sd0.13400888033126637, 32'sd-0.08097364356413865, 32'sd0.25712819218515826, 32'sd0.17077043395232558, 32'sd-0.18225215990247398, 32'sd-0.05475454893754968, 32'sd-0.06893468472830985, 32'sd-0.08497237727769724, 32'sd-0.07373200057890636, 32'sd-0.06776922462886124, 32'sd0.18101686604800846, 32'sd-0.13955902774381237, 32'sd0.13517003065864547, 32'sd-0.07060760866720553, 32'sd-0.06312043889772284, 32'sd-0.09232243767462658, 32'sd-0.03542110478004137, 32'sd-0.018519779671784087, 32'sd0.26104277562639167, 32'sd-0.1769583739430435, 32'sd-0.13255990723065297, 32'sd0.06997397523234894, 32'sd0.12092574195278412, 32'sd-0.13801961116861794, 32'sd0.04888041897938664, 32'sd0.0037718475241656, 32'sd-0.04384823216134727, 32'sd-0.14951611684873428, 32'sd-0.17530816969163782, 32'sd0.12028141209304775, 32'sd0.15539707328811816, 32'sd-0.06751074244963326, 32'sd-0.14182588519541023, 32'sd-0.17570160609077343, 32'sd-0.11348575350209644, 32'sd-0.0013000223386858813, 32'sd0.27029183827583814, 32'sd-0.20861509578126017, 32'sd0.00790830729071328, 32'sd0.1557558663208587, 32'sd-0.2973669366483478, 32'sd-0.17052946905775826, 32'sd-0.2271435169307061, 32'sd-0.18062268341383708, 32'sd0.0032586076898713646, 32'sd0.18328189389712538, 32'sd0.18556876837117373, 32'sd0.06574206734028265, 32'sd0.20023277881350754, 32'sd-0.13801546775509196, 32'sd-0.15692180258341007, 32'sd0.0620899166227393, 32'sd-0.26795597891764567, 32'sd0.1432119930815346, 32'sd-0.10003600090277813, 32'sd-0.1034813585012209, 32'sd0.08683189711362743, 32'sd-0.06575815174413832, 32'sd-0.1140975037387616},
        '{32'sd0.05102389616215056, 32'sd0.18396713545560675, 32'sd0.11999750624925755, 32'sd-0.08418231912056975, 32'sd0.07603882266780837, 32'sd-0.11987094352963139, 32'sd0.24797352786710364, 32'sd-0.049557650457219354, 32'sd-0.16816793252000686, 32'sd-0.1743380742926509, 32'sd-0.07820382825040911, 32'sd-0.006612302855629537, 32'sd0.1760039378085692, 32'sd-0.15881915717333536, 32'sd0.036203493416909496, 32'sd-0.028608194946967713, 32'sd0.1825392981789336, 32'sd-0.12221354457968424, 32'sd0.07101793363326547, 32'sd-0.007000372542348702, 32'sd-0.0732317846709776, 32'sd-0.21869809373378796, 32'sd-0.04624711889931898, 32'sd-0.08414431321076478, 32'sd-0.1035904780612196, 32'sd-0.18596498856854787, 32'sd0.03209134051066571, 32'sd0.18966548131263622, 32'sd0.12058185668896529, 32'sd-0.15675488609092988, 32'sd-0.10458116771171282, 32'sd0.03870079721379544, 32'sd0.2833055736676461, 32'sd0.18757729645006083, 32'sd0.1625277548711801, 32'sd-0.15757231613317257, 32'sd0.12272372563288954, 32'sd-0.17088877534401575, 32'sd-0.1633341683808703, 32'sd0.054457436762997455, 32'sd-0.06743790384950023, 32'sd-0.1248995865717224, 32'sd-0.12938710184784785, 32'sd0.11305315872340164, 32'sd0.05597281814614679, 32'sd0.1420355796134515, 32'sd0.05602162460298283, 32'sd0.14112853339111298, 32'sd0.18039986957913456, 32'sd-0.024947649935800644, 32'sd-0.1217061541331796, 32'sd0.11424654879291536, 32'sd0.00011508367460630769, 32'sd-0.13112758701047542, 32'sd-0.07240133579365177, 32'sd0.020350682635106632, 32'sd0.05049194442374655, 32'sd0.14033258550886918, 32'sd-0.00540420753420056, 32'sd-0.18616237148141393, 32'sd-0.23941027392077002, 32'sd-0.15538508676015556, 32'sd0.22030860416096676, 32'sd0.046060212076557555, 32'sd-0.08556261550186946, 32'sd-0.3268453706854174, 32'sd-0.16184378981084044, 32'sd-0.13258368177333235, 32'sd0.24099677410442583, 32'sd0.10768080887525598, 32'sd0.22442629049256366, 32'sd0.19489335226817814, 32'sd0.017704526329258265, 32'sd-0.1647118779624579, 32'sd-0.003667689351312404, 32'sd0.0534902978662976, 32'sd-0.04037364279975738, 32'sd0.052054928241189145, 32'sd-0.12104931917082296, 32'sd0.08876038146073804, 32'sd0.12880787844494287, 32'sd0.128148274370199, 32'sd-0.15422149426750403, 32'sd0.13862719129729298, 32'sd-0.3185153703262302, 32'sd-0.13672103759897328, 32'sd0.14921744602044903, 32'sd-0.003083649660444622, 32'sd-0.10816221668389141, 32'sd-0.06447523886860025, 32'sd0.12997378075052043, 32'sd-0.10225510082032419, 32'sd0.13347060005251665, 32'sd0.05860022112679505, 32'sd-0.03504328208592132, 32'sd-0.15896880261871224, 32'sd0.10483046207847027, 32'sd-0.045564851777577686, 32'sd-0.12219136694398164, 32'sd0.1257084516856323, 32'sd-0.16673234126078715, 32'sd0.10239609974309526, 32'sd-0.06641544735010096, 32'sd0.21870378859710626, 32'sd-0.18447063745397427, 32'sd-0.24992572684393366, 32'sd0.21965614282655346, 32'sd0.13851419535501486, 32'sd0.056754618432151446, 32'sd-0.01659650985668082, 32'sd-0.17458979331300098, 32'sd0.14486554449881994, 32'sd0.12910126591960405, 32'sd-0.038977867751988284, 32'sd-0.10150450051210358, 32'sd0.12366835960600629, 32'sd-0.0696905776918699, 32'sd-0.03773244731776892, 32'sd0.13111841127994855, 32'sd0.08362459405380619, 32'sd0.10351495789423511, 32'sd0.08137212618740394, 32'sd-0.17965802020670618, 32'sd-0.15094685409772024, 32'sd-0.0417808131866325, 32'sd-0.13357261661816933, 32'sd0.18563358985989853, 32'sd0.06411195656104525},
        '{32'sd0.12184059240536833, 32'sd-0.04659440501946958, 32'sd-0.13795639749166458, 32'sd0.13660713679213973, 32'sd0.02030088769925967, 32'sd0.08434144824251295, 32'sd0.008722780856908353, 32'sd0.02072442762909364, 32'sd-0.014801969025533495, 32'sd0.19184424238001582, 32'sd0.14087452403682277, 32'sd0.12328846175885899, 32'sd0.021401810360676093, 32'sd0.16617755274618493, 32'sd0.21538330159611477, 32'sd-0.04142795580268588, 32'sd0.260325835634789, 32'sd0.00809274866981024, 32'sd-0.011646458027416122, 32'sd0.13389974076678632, 32'sd-0.04954249942846862, 32'sd0.06489207999514018, 32'sd-0.08825444128981064, 32'sd-0.10108038679142467, 32'sd-0.07380216226426377, 32'sd0.08050036427343636, 32'sd0.17209418118725567, 32'sd0.060606633664956444, 32'sd0.024069955128522377, 32'sd0.06449295720006243, 32'sd0.04601413702538994, 32'sd0.1299346398134095, 32'sd0.03443563046865803, 32'sd-0.05666133785760118, 32'sd-0.17179753987505442, 32'sd0.14304948001707918, 32'sd-0.07900877697420872, 32'sd-0.15850384905847367, 32'sd0.08513332258065284, 32'sd0.03245951747857743, 32'sd-0.11797773540202759, 32'sd-0.1429390191329581, 32'sd0.061357682394576396, 32'sd0.155613498819865, 32'sd-0.19027699308384347, 32'sd-0.2551122351400231, 32'sd0.16469770022895724, 32'sd-0.0742824593483843, 32'sd-0.12079289602544557, 32'sd0.07199353628996676, 32'sd-0.21652031049378734, 32'sd0.2545095288059455, 32'sd-0.13933397778987872, 32'sd-0.20786150402174045, 32'sd0.11611774649598812, 32'sd0.06039128125645472, 32'sd-0.055678188942053106, 32'sd-0.13240187157128155, 32'sd0.03658078617049054, 32'sd0.12248432503608239, 32'sd-0.30780429715586016, 32'sd-0.20311917007587593, 32'sd-0.06337870483438318, 32'sd-0.07067127847115871, 32'sd-0.0127490684483825, 32'sd-0.20009745924852662, 32'sd0.19334078448971453, 32'sd0.06568201913948825, 32'sd0.14184246877969292, 32'sd0.09136307306258179, 32'sd-0.06983654664377126, 32'sd0.24954037283878885, 32'sd0.004227827490776201, 32'sd-0.04701344510727686, 32'sd-0.09431833518273486, 32'sd0.13695792058723597, 32'sd-0.029942392651860966, 32'sd0.15432783917173834, 32'sd-0.0023288365621786608, 32'sd0.09515327463964404, 32'sd0.014640302747209158, 32'sd0.011329380096741367, 32'sd0.12010864092114544, 32'sd0.27262390190360025, 32'sd0.1771719414565154, 32'sd-0.021915671334734526, 32'sd0.23409480791932272, 32'sd0.02905860516168416, 32'sd-0.11472666951647749, 32'sd-0.03268906711559755, 32'sd-0.18785097173973242, 32'sd0.05631309653642333, 32'sd0.17933346909271686, 32'sd0.1297699728545596, 32'sd-0.08562906633816239, 32'sd0.06162930745218727, 32'sd0.0978850054821972, 32'sd-0.12092620493318107, 32'sd-0.04636119181567208, 32'sd-0.21794984558498692, 32'sd-0.17090175429138077, 32'sd-0.16127576442759325, 32'sd-0.14792520198691808, 32'sd-0.20267439226113193, 32'sd-0.08618379599539323, 32'sd0.07175386312549156, 32'sd0.20382551832806511, 32'sd-0.10518826093027323, 32'sd-0.24227826371257996, 32'sd0.05943218781490338, 32'sd0.13449852273400212, 32'sd0.16947840869490302, 32'sd0.0890506789725618, 32'sd0.0865312817707955, 32'sd0.03592782215434254, 32'sd-0.07425023964767519, 32'sd0.186936300168394, 32'sd0.08268313125064651, 32'sd-0.0687636963938209, 32'sd-0.08917523411399604, 32'sd0.12885154277083546, 32'sd-0.14543165505495065, 32'sd-0.05478306776040772, 32'sd-0.23359736402102793, 32'sd-0.05148649361504322, 32'sd-0.08262416754886402, 32'sd-0.06064085774754776, 32'sd0.08015312677187011},
        '{32'sd-0.048810686640723404, 32'sd0.30316602473151355, 32'sd0.06076613388622326, 32'sd-0.07608243154499773, 32'sd-0.15196494259773544, 32'sd0.11359941638201966, 32'sd0.08012428264801184, 32'sd0.09268745046920698, 32'sd-0.16464938086977268, 32'sd0.08749709230374365, 32'sd0.043248918480207045, 32'sd0.04646640192904839, 32'sd0.1136989970690003, 32'sd0.26874313822164275, 32'sd0.009941654062665858, 32'sd0.13120533116463654, 32'sd0.17670142220075394, 32'sd0.17722928113870348, 32'sd0.18346898458960786, 32'sd0.23715918402442038, 32'sd0.00562486229589641, 32'sd0.302482844449132, 32'sd0.018825996003005968, 32'sd-0.2094181457918271, 32'sd0.16040447141348732, 32'sd0.023704624395386825, 32'sd0.18557398013173954, 32'sd0.09917122231561898, 32'sd-0.1777017137863153, 32'sd-0.011032354218580146, 32'sd0.1941662158483804, 32'sd0.176276717810828, 32'sd-0.06305258411568455, 32'sd0.07446571033757823, 32'sd-0.023258665395298226, 32'sd0.151571449326486, 32'sd0.014418343320762953, 32'sd-0.018701171214797647, 32'sd0.1563990373378777, 32'sd-0.1149141693925702, 32'sd-0.13031843894679293, 32'sd0.13695897744603894, 32'sd0.05750291679024704, 32'sd0.22319701845529527, 32'sd0.175550831048836, 32'sd-0.0681791121996501, 32'sd-0.10254129254107514, 32'sd-0.11278448609601884, 32'sd-0.07437890816368967, 32'sd-0.029256049171996538, 32'sd0.09675386039691322, 32'sd0.12710498079051596, 32'sd-0.11805156982608944, 32'sd-0.17884757011050517, 32'sd0.03207920701627004, 32'sd-0.0005420665729732017, 32'sd-0.018554418545232505, 32'sd0.12079878231360115, 32'sd0.12963817132292174, 32'sd0.20751714023233528, 32'sd-0.0714816208930994, 32'sd0.03558520681176588, 32'sd0.01522301852966126, 32'sd-0.20960531465282675, 32'sd0.01965543572096313, 32'sd-0.010049532136808419, 32'sd0.0895667818256234, 32'sd-0.16138791608131814, 32'sd0.23784985144802148, 32'sd0.11127371381780354, 32'sd0.055424528887335636, 32'sd0.17031027518910125, 32'sd-0.008315494519085587, 32'sd0.22207316647666386, 32'sd0.09853375842457078, 32'sd-0.07721053679082555, 32'sd-1.6165197607421676e-05, 32'sd0.09399590339508905, 32'sd-0.1488211851529693, 32'sd0.20373553418703974, 32'sd-0.03293274436073556, 32'sd0.010741717818041355, 32'sd0.323586407057261, 32'sd-0.06932344815875306, 32'sd0.00220602543272236, 32'sd-0.04084625244575003, 32'sd-0.03258585021374289, 32'sd0.14215695197057157, 32'sd-0.14415682588397982, 32'sd0.09231574380808025, 32'sd-0.17644248913224067, 32'sd0.03669418307365636, 32'sd-0.08045156216902931, 32'sd-0.12003103844392148, 32'sd0.038287808910250354, 32'sd0.16243023259274916, 32'sd0.0565366225519908, 32'sd-0.09980960172489121, 32'sd0.10663575965072013, 32'sd0.2585273814020687, 32'sd-0.19453791875102952, 32'sd-0.24982057307562217, 32'sd-0.1799665286880313, 32'sd0.09355054699734473, 32'sd-0.17523350183686776, 32'sd0.24436842156887356, 32'sd-0.04199344053042431, 32'sd0.08178599908876309, 32'sd0.15075630183686983, 32'sd-0.003519866139774616, 32'sd-0.14904866914831955, 32'sd-0.05984321091205968, 32'sd0.040822143179412136, 32'sd0.21280513263742357, 32'sd-0.02958561713913562, 32'sd-0.22083721782114948, 32'sd0.18941513198015913, 32'sd0.05628313292565574, 32'sd0.16018633059194248, 32'sd0.10715642451219747, 32'sd-0.05452900502000616, 32'sd-0.21323140386234624, 32'sd0.07729037950573453, 32'sd0.12698742383429976, 32'sd0.10668283732552983, 32'sd0.16163911850895052, 32'sd0.11584612082781054, 32'sd0.08454483362034106},
        '{32'sd-0.04435431675829014, 32'sd-0.02492518162722873, 32'sd-0.0922394893786112, 32'sd-0.30140912451481766, 32'sd-0.1143989512885434, 32'sd-0.07285813980628841, 32'sd0.15784841171855452, 32'sd-0.09197357947136484, 32'sd-0.23221170510261183, 32'sd-0.14466210303907878, 32'sd-8.233644275711522e-05, 32'sd-0.005729840157640575, 32'sd-0.30657430774484395, 32'sd-0.037360363968935675, 32'sd0.06846297829886176, 32'sd0.04110455293826236, 32'sd0.30441855893416875, 32'sd0.0037050653445781664, 32'sd0.03785138752619594, 32'sd0.10996287966230799, 32'sd-0.17379830811628466, 32'sd0.01075905228256752, 32'sd-0.30866769230534463, 32'sd0.14905818106773902, 32'sd-0.13847263695946457, 32'sd0.11144285638318643, 32'sd-0.12833416413744456, 32'sd-0.017028043370235453, 32'sd0.063092866706158, 32'sd0.03689942006333504, 32'sd-0.03882393802055258, 32'sd-0.0893638387655522, 32'sd-0.2622212103399947, 32'sd-0.03885237305959902, 32'sd0.2118968819210948, 32'sd-0.08066485437245247, 32'sd-0.22870331446991227, 32'sd-0.10067987768741954, 32'sd-0.02745286112834222, 32'sd-0.0522705199713724, 32'sd-0.19124707130776147, 32'sd0.06776772640841765, 32'sd0.012878772412932385, 32'sd-0.04826894921712447, 32'sd0.2665253802176805, 32'sd-0.0027466313928897097, 32'sd-0.38936425400626334, 32'sd-0.015615998002984837, 32'sd-0.24039610122583482, 32'sd-0.1486680745198858, 32'sd0.21566053198384963, 32'sd-0.24457679400353988, 32'sd-0.1365724435099573, 32'sd0.040572760879062676, 32'sd0.11530973405934968, 32'sd-0.16813995267704981, 32'sd-0.05319482979389096, 32'sd0.16258155033523022, 32'sd0.01373015682840496, 32'sd-0.06964562038006439, 32'sd0.2290342513506561, 32'sd0.12676096270038179, 32'sd-0.24357787699067765, 32'sd-0.03656435460477994, 32'sd0.18861696704962194, 32'sd-0.09120094673216096, 32'sd0.086635348794744, 32'sd0.01786004838376042, 32'sd-0.03809998705160599, 32'sd-0.1024201363115739, 32'sd0.06481282101529937, 32'sd-0.017742803141125307, 32'sd0.01159475680039052, 32'sd0.1619008324400153, 32'sd-0.08614340105983921, 32'sd0.09320026088040705, 32'sd-0.035972663214762474, 32'sd-0.15567227245516843, 32'sd-0.03889699309258703, 32'sd0.056402139620551794, 32'sd-0.005566170123125166, 32'sd-0.019564434338126983, 32'sd0.11720403313815732, 32'sd-0.10726185051189084, 32'sd-0.020126946162973225, 32'sd0.19698767597867048, 32'sd0.1076183285626391, 32'sd0.2217896878958896, 32'sd-0.11648624275097245, 32'sd-0.14429216591661553, 32'sd0.13933346193408072, 32'sd-0.030723229360192877, 32'sd-0.21570231311631313, 32'sd-0.14823823738410502, 32'sd-0.018914943505470787, 32'sd0.04423124591093855, 32'sd0.037722886169494936, 32'sd-0.20953247966842464, 32'sd-0.004978185920236896, 32'sd0.18597762601578624, 32'sd-0.2661946902094207, 32'sd0.0013225976578255137, 32'sd-0.2334163950205284, 32'sd0.032459817647691507, 32'sd-0.09053973261350104, 32'sd-0.024583893152889467, 32'sd-0.20209710491238744, 32'sd0.05587939242857886, 32'sd0.02587880500943274, 32'sd-0.004770879478872604, 32'sd-0.10615679098986364, 32'sd-0.15870406637717396, 32'sd0.20611341297180003, 32'sd0.18999893350257804, 32'sd-0.068358405612737, 32'sd-0.13007817643278524, 32'sd0.07965597142205393, 32'sd0.08072302873622433, 32'sd0.1270746411726309, 32'sd0.018908909242842067, 32'sd0.014804891372289904, 32'sd-0.03177487695305075, 32'sd0.11855552966923728, 32'sd-0.07408041402627731, 32'sd-0.15828792083646417, 32'sd0.024038824989873163, 32'sd0.08719465947211408, 32'sd0.13882809831815915},
        '{32'sd0.075245076016843, 32'sd-0.03913380891693224, 32'sd0.0465330473866347, 32'sd0.02768990438282041, 32'sd-0.08159554202663742, 32'sd-0.09192659258849822, 32'sd-0.09470581020774604, 32'sd-0.0865726996893167, 32'sd-0.16809694500166053, 32'sd0.1472879447040246, 32'sd-0.017708605986691883, 32'sd0.09831106938527671, 32'sd0.17250152700443266, 32'sd-0.14225757765223818, 32'sd-0.14842883296836437, 32'sd0.11479117426561174, 32'sd0.16365269609820593, 32'sd-0.2704140475629073, 32'sd-0.039895773047398365, 32'sd0.03504848348337571, 32'sd-0.22613488834998108, 32'sd-0.05843378598816249, 32'sd-0.1605234626842765, 32'sd0.013336773035910063, 32'sd-0.14123800884448123, 32'sd-0.12675546503820553, 32'sd0.20187737536777092, 32'sd0.008197154144210699, 32'sd-0.22972329882473597, 32'sd0.10507909796823678, 32'sd0.018810678841259667, 32'sd-0.21452723494026602, 32'sd-0.06590068574025548, 32'sd-0.049522972166009226, 32'sd0.2025253918991844, 32'sd-0.14306616433161132, 32'sd0.20905445866376962, 32'sd-0.12234745531581967, 32'sd0.1268837950676065, 32'sd0.027477067161656765, 32'sd0.15879415785239476, 32'sd0.16594493256619075, 32'sd0.20787463683653126, 32'sd0.040880282120367435, 32'sd0.1898423172564554, 32'sd0.1370635665823767, 32'sd0.24232963739960398, 32'sd0.0014241905767743226, 32'sd0.0910989171539913, 32'sd0.12091568059427138, 32'sd0.0003836495031417332, 32'sd-0.07972739672923558, 32'sd0.05336516095713287, 32'sd0.16043436559667323, 32'sd-0.01746346661744469, 32'sd-0.15467469565718092, 32'sd0.2393639677185007, 32'sd-0.12427101991361668, 32'sd-0.1931498078267209, 32'sd-0.01917373871274713, 32'sd-0.08133231479612144, 32'sd-0.10761083007865149, 32'sd0.11569961239496085, 32'sd0.06033244351693415, 32'sd0.1432257678325645, 32'sd0.07815216028359541, 32'sd0.012583896120981156, 32'sd0.19827283638963636, 32'sd-0.06237672609934741, 32'sd-0.23196442495312058, 32'sd0.06247664934029353, 32'sd0.08883425397332137, 32'sd0.02991075419937694, 32'sd0.09414963439083762, 32'sd0.11347373104909586, 32'sd0.1602686051306, 32'sd0.10752606073825378, 32'sd0.2510830034263254, 32'sd-0.08729106967156583, 32'sd0.1113466695435354, 32'sd-0.21971671205875895, 32'sd-0.017464312243467076, 32'sd0.09250205502446232, 32'sd0.1789300448087912, 32'sd0.10590276642983928, 32'sd-0.1865024909151068, 32'sd-0.11082985456699598, 32'sd-0.25123736952051284, 32'sd-0.09986143503851934, 32'sd0.06282439992534933, 32'sd0.09261827946587216, 32'sd-0.10370972599836707, 32'sd0.0469075613535912, 32'sd0.05722598128549231, 32'sd0.06682718343928985, 32'sd-0.21520402331423877, 32'sd-0.023272910345646287, 32'sd0.13817805821330834, 32'sd0.09756735404495856, 32'sd0.12770356992086435, 32'sd0.057327399012392276, 32'sd0.00010412805582157847, 32'sd-0.12410302767230312, 32'sd-0.08971851855503456, 32'sd-0.1776893332711896, 32'sd-0.07783786851579767, 32'sd-0.20818739635041647, 32'sd0.11170808371803125, 32'sd0.10759128532806721, 32'sd-0.05016570974913993, 32'sd0.19303037270365525, 32'sd-0.14326371733597282, 32'sd-0.04356444798004441, 32'sd0.0656623138325769, 32'sd0.1931360765834376, 32'sd0.1376512945681606, 32'sd-0.17778403794568795, 32'sd0.1695936482763491, 32'sd0.002955124661158645, 32'sd0.03265282394759474, 32'sd0.17648202895995008, 32'sd0.1477970716333417, 32'sd0.047182867754593585, 32'sd-0.2325257042435153, 32'sd0.21292725329481837, 32'sd-0.12238149520427102, 32'sd0.26016490049608787, 32'sd0.051111196404152945},
        '{32'sd-0.09906447219937477, 32'sd-0.07761347458205443, 32'sd-0.19544070083716505, 32'sd0.1505527819209299, 32'sd0.04334716621651655, 32'sd-0.06005712337871036, 32'sd-0.20911288354012764, 32'sd0.16775930353348772, 32'sd0.13617237979700503, 32'sd0.02407184652188252, 32'sd-0.10559601224104362, 32'sd-0.052207664913781975, 32'sd-0.0457642990860882, 32'sd-0.10061998427299111, 32'sd-0.2256430401781246, 32'sd-0.1810307222416693, 32'sd0.1700052389665425, 32'sd-0.23314855483704514, 32'sd0.027486568710227696, 32'sd-0.014898588782961596, 32'sd-0.041038465329919616, 32'sd0.05574244142248325, 32'sd0.11394833452385202, 32'sd0.08878412293437199, 32'sd-0.25946979897652667, 32'sd0.17123514172481413, 32'sd0.03819074667540518, 32'sd-0.2846876867205207, 32'sd0.1226964813488115, 32'sd0.16018171108112644, 32'sd-0.08811715673808893, 32'sd-0.005239818175013342, 32'sd0.12119209361676866, 32'sd0.013549186231488722, 32'sd-0.06402357623819381, 32'sd-0.14458102064754447, 32'sd0.04212622472194155, 32'sd0.07725441931828127, 32'sd0.04283800881459935, 32'sd0.08382809845930043, 32'sd0.05153385534946064, 32'sd0.14180500777541044, 32'sd0.1794069720204979, 32'sd0.08412056765845329, 32'sd-0.009315053873670289, 32'sd0.3024714738128755, 32'sd-0.07113454553442229, 32'sd-0.02312507730763905, 32'sd-0.08126934105226692, 32'sd-0.1251899887540951, 32'sd0.05616717994394306, 32'sd-0.024041573006035738, 32'sd-0.10561726381245512, 32'sd0.15430575357347567, 32'sd-0.122694432950252, 32'sd0.008150025215949933, 32'sd-0.15549463036479744, 32'sd0.023619996811489047, 32'sd0.07715157188200814, 32'sd0.2374566494507654, 32'sd-0.10957473107480957, 32'sd0.15845405001621185, 32'sd0.13749649427905095, 32'sd0.09532753999971612, 32'sd0.05360449631393532, 32'sd0.004236868260017339, 32'sd0.08425011633242313, 32'sd-0.02957708845923808, 32'sd-0.09882633460642433, 32'sd-0.08510998939149533, 32'sd-0.27034771182976275, 32'sd-0.30467008711141236, 32'sd-0.1673462484615944, 32'sd0.18246880525469764, 32'sd-0.09003789903044956, 32'sd0.2406363558399259, 32'sd0.17672104180261336, 32'sd-0.3080581172757816, 32'sd0.22130711069931666, 32'sd-0.0745386790930619, 32'sd-0.018523800329763893, 32'sd0.18291100329167442, 32'sd0.16794887694338773, 32'sd0.12355524963559751, 32'sd0.31749354775055094, 32'sd0.15746361671904902, 32'sd-0.09047107728480959, 32'sd-0.11709460101154057, 32'sd0.060656692514397294, 32'sd0.11598924917558731, 32'sd-0.05016125276262772, 32'sd0.12707693264147385, 32'sd-0.038323992237986736, 32'sd0.06444553867540372, 32'sd0.054917743528422144, 32'sd-0.1230878519557354, 32'sd-0.04271231733479459, 32'sd-0.007919121786674031, 32'sd0.14948171590879894, 32'sd0.2062283540513715, 32'sd-0.12411142431440653, 32'sd-0.1885719606842057, 32'sd0.09663116253588067, 32'sd0.16849202991731846, 32'sd-0.07146928580717186, 32'sd-0.14402700111631775, 32'sd-0.10990781617308866, 32'sd-0.16937310074779818, 32'sd0.10281278701189085, 32'sd0.11295023589464336, 32'sd0.0883386259554079, 32'sd-0.3280219403452036, 32'sd-0.23727298668146146, 32'sd0.18643834870376277, 32'sd-0.03739088549223291, 32'sd-0.19678344533347802, 32'sd0.09011332436599778, 32'sd0.05415469442821297, 32'sd0.04860709832751812, 32'sd0.01860304341248138, 32'sd-0.305202691049943, 32'sd0.08252793737398949, 32'sd-0.030732306496257866, 32'sd-0.12458561244929321, 32'sd-0.2006468389761952, 32'sd-0.21534151365441767, 32'sd-0.07834155650268763, 32'sd0.05277857472698837},
        '{32'sd0.07410876000946774, 32'sd-0.3698238409135545, 32'sd-0.02003742260104424, 32'sd0.20440382959159675, 32'sd0.14818181369683395, 32'sd-0.2751356615459531, 32'sd-0.0454515167795998, 32'sd0.03931237313367676, 32'sd0.15092042032698774, 32'sd-0.01508526287092608, 32'sd-0.07480912584339353, 32'sd0.049900556696270276, 32'sd0.027230794076540086, 32'sd0.11690010876295255, 32'sd0.035347834315609686, 32'sd0.011401827205633663, 32'sd0.02139576087635575, 32'sd0.14985418690199784, 32'sd-0.03035640728805698, 32'sd0.23461534167364262, 32'sd0.1439709536660004, 32'sd-0.0706381342860444, 32'sd-0.019756928425403927, 32'sd0.11401112356749185, 32'sd-0.41867527122015147, 32'sd-0.08957686901565454, 32'sd-0.27638540626610336, 32'sd-0.10605054863922113, 32'sd-0.18486218875322186, 32'sd0.029014943512712752, 32'sd-0.1720131880705656, 32'sd0.08513730261538163, 32'sd-0.07510670467632131, 32'sd0.17720962221303818, 32'sd0.24533261981992655, 32'sd-0.08648185339644043, 32'sd-0.07546926130435276, 32'sd-0.26771377385464035, 32'sd0.14244818768710643, 32'sd0.289826832662894, 32'sd0.059783203315114, 32'sd0.05753172720040969, 32'sd0.18176190220128996, 32'sd-0.2736392701153145, 32'sd0.10573701848794158, 32'sd-0.06477298777751232, 32'sd-0.1402424124985251, 32'sd-0.12221106588418444, 32'sd-0.07230540967321877, 32'sd0.11812231897616403, 32'sd-0.15554517261922618, 32'sd-0.19903717090221373, 32'sd-0.16866404268409974, 32'sd-0.016442178374247197, 32'sd0.09834815639235403, 32'sd0.15198949410891263, 32'sd-0.14825942954856233, 32'sd0.006524286536708208, 32'sd-0.18026417521476082, 32'sd-0.15319493558158373, 32'sd0.21370752065097187, 32'sd0.14492944086909107, 32'sd-0.03620429183136038, 32'sd0.2336614867588597, 32'sd-0.0218649146140083, 32'sd-0.21163702381168092, 32'sd0.005703938667330594, 32'sd0.15327783960163394, 32'sd-0.19915761088338377, 32'sd-0.03999249887980887, 32'sd-0.10476497016722366, 32'sd0.12056655263557096, 32'sd0.28626244887185687, 32'sd0.0548867383372998, 32'sd-0.13777328431940686, 32'sd-0.3430487553651127, 32'sd-0.0674696526952078, 32'sd0.09225366759361789, 32'sd0.13020766922258406, 32'sd0.015639227699514292, 32'sd-0.004302945586581507, 32'sd-0.22557098211079582, 32'sd-0.05463542288481857, 32'sd0.06594203756965902, 32'sd0.04410839719290663, 32'sd-0.0450732231165814, 32'sd-0.02094881802681037, 32'sd-0.1005592534809067, 32'sd-0.0727462021281018, 32'sd-0.19586569076641366, 32'sd-0.13844802911746718, 32'sd-0.07164123245765469, 32'sd0.15869871295664162, 32'sd-0.14593497018768883, 32'sd0.18399763790017454, 32'sd0.12838628632983004, 32'sd-0.04640873820894002, 32'sd0.1669945768963897, 32'sd0.14117277466779118, 32'sd-0.24637971188206237, 32'sd-0.150249976843613, 32'sd0.1467446748028905, 32'sd-0.18253809515521513, 32'sd-0.18638340414436366, 32'sd-0.08951239963800073, 32'sd-0.21300446838055867, 32'sd-0.029673074838750126, 32'sd-0.2518835621555524, 32'sd0.07976244824192158, 32'sd0.25019539786891776, 32'sd0.04698106787411035, 32'sd0.01714780755747424, 32'sd0.313405338995811, 32'sd-0.07134581980470309, 32'sd-0.07270467913731161, 32'sd-0.14170516306745778, 32'sd0.1772259692949172, 32'sd-0.13675103238119293, 32'sd0.0713975566734599, 32'sd0.09263457215012476, 32'sd-0.07369149596161789, 32'sd0.09826248868002295, 32'sd0.10936846228735082, 32'sd0.00443126164607825, 32'sd0.027009424879216055, 32'sd0.0024062929821517206, 32'sd0.09671364509160418, 32'sd0.15099284394407242},
        '{32'sd0.17477522016674352, 32'sd-0.15106286741033131, 32'sd0.02123218388222262, 32'sd0.1456975712548906, 32'sd-0.1413865456320702, 32'sd-0.1018955667481582, 32'sd0.14915619574317573, 32'sd-0.01953568632682688, 32'sd-0.16592770073899568, 32'sd-0.14296019001057522, 32'sd-0.030556708148173267, 32'sd-0.04877597582838003, 32'sd-0.21961314605586787, 32'sd0.09666192855358947, 32'sd0.12895259828016145, 32'sd-0.3534200689492139, 32'sd0.16432272823651228, 32'sd-0.16135012465502516, 32'sd0.00961401366852643, 32'sd0.1496330534520952, 32'sd0.11617274814268701, 32'sd0.023289817547403297, 32'sd-0.06763091465908098, 32'sd-0.008197848628751735, 32'sd-0.17416269973117807, 32'sd0.027182581389673836, 32'sd-0.15327765817018907, 32'sd-0.05605556186611474, 32'sd-0.22305908470902663, 32'sd-0.2977917512026326, 32'sd0.021063645860312143, 32'sd-0.15697664534176978, 32'sd-0.10278588805501489, 32'sd0.004065153726197087, 32'sd0.050390257594099694, 32'sd-0.3243868360186187, 32'sd0.16771025437680243, 32'sd-0.04164938023612343, 32'sd0.046218266230172195, 32'sd0.2912191857147569, 32'sd-0.1018505787336276, 32'sd0.12980312448738593, 32'sd-0.1620710825429281, 32'sd-0.06955444553091886, 32'sd0.19291541065631435, 32'sd0.17348151787298477, 32'sd-0.32737611222489144, 32'sd-0.27122317514325484, 32'sd-0.14530892235457313, 32'sd-0.21197002417063157, 32'sd-0.20154692540725758, 32'sd-0.09992217697757624, 32'sd-0.033399850205374296, 32'sd0.07984293127555364, 32'sd0.3154841134020625, 32'sd-0.11668817709490545, 32'sd0.020443700320952975, 32'sd0.06281231475761416, 32'sd0.15854024079665546, 32'sd0.2109047043601334, 32'sd0.008173964732257677, 32'sd0.1955864992341671, 32'sd0.1008766333563915, 32'sd0.2613257345416747, 32'sd-0.024678195727534793, 32'sd-0.010397483544989126, 32'sd-0.1480777284521407, 32'sd-0.08488719861565025, 32'sd-0.12182604248123406, 32'sd0.06603398231866758, 32'sd0.19258757899272547, 32'sd-0.1812998213841102, 32'sd-0.10364253270077149, 32'sd-0.19209813465465303, 32'sd-0.07495063981655446, 32'sd-0.035079073993159446, 32'sd-0.018725474683167518, 32'sd0.03987767698409049, 32'sd0.08330417793677437, 32'sd0.04650348514715095, 32'sd-0.056746547181734476, 32'sd0.1126215175870737, 32'sd0.21375730560737286, 32'sd-0.11776778175749003, 32'sd0.1249423179332994, 32'sd0.042891779001685656, 32'sd0.11066485289835294, 32'sd0.006100359558601628, 32'sd0.10426749683608187, 32'sd-0.16674561768065732, 32'sd0.21094598215267954, 32'sd0.03382288764465471, 32'sd-0.21523452410118657, 32'sd-0.16401656083149246, 32'sd-0.0789085423445792, 32'sd-0.0050838424202658185, 32'sd-0.19381057121121176, 32'sd0.020283815415296346, 32'sd-0.07790235273125884, 32'sd0.1756309069820054, 32'sd0.03201008238951916, 32'sd-0.043037841603278594, 32'sd-0.1420130758727873, 32'sd0.06523832835198576, 32'sd-0.06301664528008516, 32'sd-0.14405411283463274, 32'sd-0.11568265336314067, 32'sd0.10291748501887055, 32'sd0.11072859412647082, 32'sd-0.08718995681891589, 32'sd0.18291697546402327, 32'sd-0.17673065254506576, 32'sd0.0888324223483673, 32'sd0.1763832124431195, 32'sd-0.07322266501727756, 32'sd0.052802688871767575, 32'sd0.0317402317150562, 32'sd0.26113620785382957, 32'sd0.08525316599144657, 32'sd0.021409176860113278, 32'sd-0.1268784173886004, 32'sd-0.008444476006865556, 32'sd0.03276775317149889, 32'sd-0.15845170413224413, 32'sd-0.13738962671506366, 32'sd-0.09257734087202764, 32'sd-0.10348408565383774, 32'sd-0.009694914562173569},
        '{32'sd-0.017765557196728565, 32'sd0.10951080679153598, 32'sd-0.19676619986268418, 32'sd0.14048328243600366, 32'sd-0.2339625862591353, 32'sd-0.05708091569040154, 32'sd-0.015245574492901542, 32'sd-0.2515859008992347, 32'sd-0.090233702881789, 32'sd0.19781939313404495, 32'sd0.10549515984477355, 32'sd0.05779360665797868, 32'sd0.018425739745139436, 32'sd-0.00645825704183993, 32'sd0.1213121114496166, 32'sd0.197150567107264, 32'sd0.05157954508883906, 32'sd-0.09924468756182589, 32'sd-0.056369932736011256, 32'sd-0.24778263959090174, 32'sd-0.03891972653723818, 32'sd-0.21715680416524688, 32'sd0.08614323641844945, 32'sd-0.03428009460736567, 32'sd0.24330268445414657, 32'sd0.14498875042231196, 32'sd-0.06870169325798926, 32'sd0.14595202209948868, 32'sd-0.08072295583463648, 32'sd-0.07012627958837797, 32'sd0.06031928576555699, 32'sd-0.19292658792197973, 32'sd0.19714304642545596, 32'sd-0.1238520021895875, 32'sd0.23352155187627974, 32'sd-0.117730631227004, 32'sd0.21225655049474387, 32'sd0.11268467767122449, 32'sd0.10877625910797915, 32'sd0.169806039675829, 32'sd0.08501379559303446, 32'sd-0.07463077259273851, 32'sd0.07882084211373323, 32'sd-0.045356470388574315, 32'sd-0.30158704896949484, 32'sd0.1672125489423274, 32'sd0.0850923302978617, 32'sd0.08237015225251813, 32'sd0.1149474550442372, 32'sd-0.20340740880321723, 32'sd-0.006449055787213567, 32'sd-0.03564360671527101, 32'sd0.10899920778008775, 32'sd-0.1310041722356102, 32'sd0.00753244034850818, 32'sd-0.13595132566740073, 32'sd0.1046516098482061, 32'sd0.04617695361673962, 32'sd0.05871930193299951, 32'sd-0.25591202539508223, 32'sd-0.0011182917212472566, 32'sd0.0853293581255235, 32'sd0.05929150708950429, 32'sd-0.11015190933648014, 32'sd-0.07697824087099273, 32'sd0.015845946774903114, 32'sd0.028332664555284843, 32'sd0.20378433656673944, 32'sd-0.18844498558810588, 32'sd0.03990367718224957, 32'sd-0.06292157566363817, 32'sd0.27431220470626944, 32'sd0.3103234800301326, 32'sd-0.18127157587736278, 32'sd0.1566892329909978, 32'sd-0.05625473345535878, 32'sd0.1747345138108729, 32'sd-0.02292501019865844, 32'sd0.06372414843354145, 32'sd-0.1315133964226983, 32'sd-0.2327970559532467, 32'sd0.03667262089214835, 32'sd-0.20318433247555917, 32'sd-0.19466410001011758, 32'sd-0.14115216568407996, 32'sd0.011437246536348493, 32'sd0.0782219410394631, 32'sd-0.02936770965108737, 32'sd0.11766428187810173, 32'sd0.19643897876793426, 32'sd0.035218119934582355, 32'sd0.08647850301182426, 32'sd0.24240973217084227, 32'sd-0.15200776218591636, 32'sd0.12528892192329563, 32'sd0.060506660985970157, 32'sd0.08724945980439427, 32'sd0.09185516937411443, 32'sd0.026275893424788848, 32'sd-0.19270051095846563, 32'sd-0.0026704182565296455, 32'sd-0.07669915849197154, 32'sd-0.08259294331897526, 32'sd-0.004640388523644893, 32'sd0.05674025717587538, 32'sd-0.11565156818682289, 32'sd0.011148615304718732, 32'sd-0.1647560962551378, 32'sd0.004288557818583702, 32'sd0.053942896711885874, 32'sd0.12026423722476674, 32'sd-0.12152733394547603, 32'sd-0.26880912361791204, 32'sd-0.23365609480430818, 32'sd0.005318258018665784, 32'sd0.024172203910285763, 32'sd-0.00527313809152595, 32'sd-0.028043766644311695, 32'sd-0.11378455780823567, 32'sd0.07602517780494529, 32'sd-0.07945165306389174, 32'sd-0.15845956043788406, 32'sd0.10795920265903923, 32'sd-0.12327094758002098, 32'sd0.19518410518717896, 32'sd0.1635516176115474, 32'sd-0.11188084229957812, 32'sd0.1368674064932967},
        '{32'sd0.1166156455072414, 32'sd0.030671042193226004, 32'sd0.03236720374794033, 32'sd0.06611003019536787, 32'sd-0.03789545048057319, 32'sd0.17001805240565748, 32'sd-0.01808534640031825, 32'sd0.2569434452621486, 32'sd0.020241439161634154, 32'sd-0.1311225647032668, 32'sd-0.14841418436950865, 32'sd0.11669774381932074, 32'sd0.16663642646073912, 32'sd-0.17929719658118792, 32'sd-0.056056009775884076, 32'sd-0.07172776818198703, 32'sd-0.01546583068393177, 32'sd0.20393556094367218, 32'sd0.06453717187773046, 32'sd0.0340427700948983, 32'sd0.2910208358060136, 32'sd0.2422373863198954, 32'sd-0.07372277549365587, 32'sd0.04821722484791069, 32'sd0.13338276313995182, 32'sd-0.14198310548826576, 32'sd-0.21254274198764184, 32'sd0.16360522568641384, 32'sd-0.150318559208245, 32'sd-0.18877997164001784, 32'sd-0.0056339228696265465, 32'sd-0.05922280497505796, 32'sd-0.16449126638366596, 32'sd-0.17387731131389142, 32'sd-0.01344134394167502, 32'sd0.1851831017514107, 32'sd-0.00470582411190241, 32'sd0.16329902670535962, 32'sd-0.12007323150704498, 32'sd-0.08823637759265364, 32'sd0.09782799818013717, 32'sd0.0856958982672063, 32'sd-0.05780948045558916, 32'sd0.00798551188846682, 32'sd-0.025733992460653974, 32'sd-0.04902438622097052, 32'sd0.20355551816688, 32'sd-0.1573983017664462, 32'sd-0.013850233408703835, 32'sd0.13545414875705575, 32'sd-0.09663221079701809, 32'sd-0.14730405101428862, 32'sd0.000850598232664304, 32'sd0.1403761101052389, 32'sd-0.06180458411120808, 32'sd-0.09227351830427755, 32'sd0.21642262773969517, 32'sd0.07366787344005588, 32'sd0.03659141133534531, 32'sd-0.21513782093056646, 32'sd-0.10113352218348871, 32'sd-0.13422159778916135, 32'sd-0.2049688923022194, 32'sd0.09871335063533693, 32'sd0.30809233904616123, 32'sd0.03995328921169671, 32'sd-0.130213845248045, 32'sd0.04106365421505669, 32'sd-0.23005370003347342, 32'sd0.045179026559432164, 32'sd-0.07984856170475622, 32'sd0.14101814023199938, 32'sd0.0776373028222917, 32'sd0.192441111034226, 32'sd0.06225107181230641, 32'sd0.059416445909600726, 32'sd-0.02921255644547632, 32'sd0.17397268640067098, 32'sd0.11027731277347465, 32'sd-0.18485485752368805, 32'sd0.12464421702920774, 32'sd-0.037780157526297514, 32'sd0.011606708399937484, 32'sd-0.10223484578477893, 32'sd-0.16668174154643461, 32'sd-0.14803338795339543, 32'sd0.04011915362875131, 32'sd0.24465891886962138, 32'sd-0.07633988655642152, 32'sd-0.10546137023615079, 32'sd-0.10199586007634964, 32'sd-0.2033959008104763, 32'sd-0.24117234566523477, 32'sd0.17147421038555707, 32'sd0.1266001892826685, 32'sd-0.12875146050106212, 32'sd0.030335460600788927, 32'sd0.20728667767228076, 32'sd0.12995236496416374, 32'sd-0.08161235076507281, 32'sd0.09893971582593175, 32'sd-0.06655373932699662, 32'sd0.007115918981789003, 32'sd0.2166646927025192, 32'sd-0.3042729254524271, 32'sd-0.11544409815773626, 32'sd0.12827412329451987, 32'sd0.05492518146321429, 32'sd-0.10779486616075615, 32'sd0.0852640112857219, 32'sd-0.30686457525043054, 32'sd-0.04571714728154185, 32'sd0.17757251754061484, 32'sd-0.004972054898558164, 32'sd-0.11988750156071143, 32'sd0.21352351805629524, 32'sd0.1409211913506407, 32'sd-0.01779786523757261, 32'sd0.08730953082606506, 32'sd-0.25012649026956424, 32'sd0.2592237808829766, 32'sd0.1611411413392977, 32'sd0.07282411812380617, 32'sd0.0414622824794083, 32'sd-0.055295480983781904, 32'sd0.10836026149019633, 32'sd-0.07311508562805509, 32'sd-0.051369139006498456},
        '{32'sd-0.09897381038174684, 32'sd-0.06084022662769187, 32'sd-0.06067324172040819, 32'sd-0.08666087739712129, 32'sd-0.07113757022871009, 32'sd0.09617650817307166, 32'sd-0.15172749353457646, 32'sd-0.1337376221512761, 32'sd-0.03333040629131448, 32'sd0.21337179406009726, 32'sd0.1698732974406922, 32'sd0.051422782479230544, 32'sd0.020493218127828644, 32'sd0.0520736509972999, 32'sd-0.053716014205451156, 32'sd0.09664726340490254, 32'sd-0.0442947961839649, 32'sd-0.13197486660010405, 32'sd-0.18991182091488196, 32'sd0.07952260553737402, 32'sd-0.12217129933124132, 32'sd0.18063835716772178, 32'sd-0.18678647973434534, 32'sd0.04500344101434037, 32'sd-0.16349633743469202, 32'sd0.12592814696504015, 32'sd0.10116209903582032, 32'sd-0.1394749221194745, 32'sd0.16655362071933796, 32'sd-0.17466292773748118, 32'sd-0.00410531497627071, 32'sd0.24863074836759566, 32'sd-0.08252779514283093, 32'sd-0.19868423447669478, 32'sd-0.1484842559885592, 32'sd-0.046440662092525134, 32'sd0.0740107490920701, 32'sd-0.008536468707699946, 32'sd-0.1777939224713827, 32'sd-0.1426214791541076, 32'sd0.13382793791107803, 32'sd-0.1561010457230357, 32'sd-0.29184390919065, 32'sd0.045078017224931134, 32'sd0.09519056083463603, 32'sd0.06018720804145974, 32'sd0.2893201879685878, 32'sd-0.1145315143975961, 32'sd-0.2573545756199081, 32'sd-0.14804873451192296, 32'sd0.2741554739158564, 32'sd0.1451218280140441, 32'sd-0.24531299625455108, 32'sd-0.15192495203528303, 32'sd0.2024042911420158, 32'sd0.0008900002664995216, 32'sd0.09474423131806838, 32'sd0.19968289499352465, 32'sd0.054617452722186786, 32'sd-0.20450457917563608, 32'sd0.18162026108092355, 32'sd-0.006362187819479246, 32'sd-0.15500452051166497, 32'sd-0.005782357660171557, 32'sd-0.026868840684830544, 32'sd-0.05695885092809149, 32'sd0.056138682790178356, 32'sd0.17242739999891563, 32'sd-0.3302957478536988, 32'sd-0.05777998192104742, 32'sd-0.11335533285402133, 32'sd0.12110020679166418, 32'sd0.3069555992997738, 32'sd-0.029460583584273475, 32'sd0.006398333910515985, 32'sd-0.04252100733767392, 32'sd0.13875215192271317, 32'sd-0.004427061774737933, 32'sd0.1656941196625896, 32'sd0.19529110472297018, 32'sd-0.2640129487111787, 32'sd-0.1225010038720604, 32'sd-0.14671614509995426, 32'sd-0.11943706538038694, 32'sd-0.056728897269148454, 32'sd0.18884890662378406, 32'sd-0.1826255792404504, 32'sd0.17646278264679313, 32'sd0.097476119400634, 32'sd-0.029376277161037825, 32'sd0.11181950884230557, 32'sd0.0869374353959709, 32'sd-0.13150344128448022, 32'sd0.047767673202996554, 32'sd0.00465368740386221, 32'sd0.051831432829848846, 32'sd-0.0544916579811813, 32'sd-0.1909841942984574, 32'sd0.09631015301939738, 32'sd0.022907749038912555, 32'sd0.02694824095296076, 32'sd-0.03232527605646129, 32'sd-0.15687786760051783, 32'sd-0.23271643234230413, 32'sd0.08252045176587183, 32'sd-0.08598610159713303, 32'sd-0.005438177574522009, 32'sd0.13136346723432388, 32'sd-0.05778330793785782, 32'sd0.1603799449472058, 32'sd-0.15480834650230493, 32'sd-0.22748067994835944, 32'sd-0.08691785559656856, 32'sd-0.18722421248759105, 32'sd0.05098008073321894, 32'sd0.18913203215383118, 32'sd0.14390954009737167, 32'sd0.10270850891522133, 32'sd0.015165484103972305, 32'sd0.1385706412897554, 32'sd-0.10162080155164953, 32'sd0.111974795282924, 32'sd-0.03421324066090248, 32'sd0.01661778879093637, 32'sd0.034038829485248064, 32'sd0.30419138842475685, 32'sd0.009303889199830101, 32'sd0.13865468847908097},
        '{32'sd0.032608148660147065, 32'sd0.12644712679047776, 32'sd-0.002139523101502016, 32'sd0.10471571546629715, 32'sd-0.15802838487639678, 32'sd-0.19067860197149944, 32'sd-0.013522736716533422, 32'sd-0.23739222180810032, 32'sd-0.16994352273526253, 32'sd-0.10527047278383529, 32'sd0.22454030350628748, 32'sd-0.02182407973744482, 32'sd-0.018313617659144337, 32'sd-0.01168985861670653, 32'sd0.08885142823987825, 32'sd-0.13467618004877732, 32'sd-0.08137190040374832, 32'sd-0.004628396147177128, 32'sd0.027851176223524572, 32'sd-0.048902076402609046, 32'sd-0.3397498782891119, 32'sd0.13066320267658388, 32'sd0.024493597445591805, 32'sd-0.1329525129052451, 32'sd0.03927791074884537, 32'sd0.27151369097550293, 32'sd0.2420141391753665, 32'sd0.21287387034722347, 32'sd0.19082693729893196, 32'sd-0.23838818877400667, 32'sd-0.3139049931015949, 32'sd0.0522397768098166, 32'sd-0.09567483993669618, 32'sd-0.10219641289821392, 32'sd-0.08253324551447429, 32'sd0.18859465227679628, 32'sd-0.25201335862743585, 32'sd-0.10024601423540036, 32'sd0.043867881815725436, 32'sd0.049215918528964626, 32'sd0.04666780136090155, 32'sd-0.011336392095159709, 32'sd-0.042662360688752746, 32'sd0.17630765644623997, 32'sd0.02867465609940094, 32'sd0.22418117269827403, 32'sd-0.003030827608336019, 32'sd0.09626120997214928, 32'sd0.1289312273030922, 32'sd-0.04223425438092452, 32'sd0.05095031836497392, 32'sd0.135401875869459, 32'sd-0.0211437141342836, 32'sd0.22173041495657594, 32'sd-0.006334712468207421, 32'sd0.040644952519364175, 32'sd-0.09721865903551517, 32'sd0.007795922261967962, 32'sd-0.025780113662631308, 32'sd0.21604813449985055, 32'sd0.010193602273538872, 32'sd-0.14415460078434725, 32'sd-0.1582454509611696, 32'sd0.12814637476563884, 32'sd0.054974722812218726, 32'sd0.13133504864017914, 32'sd-0.062487312954939055, 32'sd0.0036951921195134685, 32'sd-0.09148369508531255, 32'sd0.05286570671086057, 32'sd0.11751682616895215, 32'sd-0.1839164906582695, 32'sd-0.2016271673170593, 32'sd-0.16723222962697692, 32'sd-0.1865316958513193, 32'sd0.19737022454620756, 32'sd-0.14427810689233386, 32'sd0.11236237791094147, 32'sd-0.03776375465095972, 32'sd0.027935757372136532, 32'sd-0.02119224733550027, 32'sd-0.03705543222032156, 32'sd0.03622519036053175, 32'sd-0.09790105137528049, 32'sd0.034487689746141, 32'sd-0.019614807138826806, 32'sd0.030594219692364522, 32'sd-0.14038394493095643, 32'sd-0.0960685370669436, 32'sd-0.13512967011776608, 32'sd0.004865358842701544, 32'sd-0.1395943240411702, 32'sd0.28553403191545323, 32'sd0.13199196913134667, 32'sd-0.18473003802499322, 32'sd0.09354414656028118, 32'sd0.1169889740234883, 32'sd-0.02753672114315139, 32'sd-0.005062086112304186, 32'sd-0.16374462558734018, 32'sd0.058332476404228305, 32'sd0.18414754735300007, 32'sd0.15898779802180682, 32'sd-0.002173268233668894, 32'sd-0.17139463016251077, 32'sd-0.14954110606579157, 32'sd0.10891391906925074, 32'sd-0.0738831556003839, 32'sd0.16967501359087045, 32'sd-0.05254432213663226, 32'sd-0.23128917052266448, 32'sd-0.06561257425072735, 32'sd-0.018677588781642884, 32'sd0.06512536197293778, 32'sd0.033340999329053975, 32'sd-0.07237459178701144, 32'sd0.046171073202582805, 32'sd-0.17621688336256933, 32'sd-0.0197100941451455, 32'sd0.06796659397509962, 32'sd0.23224754398767664, 32'sd-0.024929040752347826, 32'sd0.06459810747068262, 32'sd0.038630573757422244, 32'sd-0.15399631163453684, 32'sd0.19382753750352288, 32'sd0.0622740640326304, 32'sd0.05846946812866302},
        '{32'sd-0.21440814547723777, 32'sd-0.08816330847017523, 32'sd0.13532810593871192, 32'sd0.0141933290683429, 32'sd0.07727893495083235, 32'sd0.03902006378284128, 32'sd-0.20239058540010982, 32'sd-0.010084133522422975, 32'sd0.14888484266232707, 32'sd-0.04320867115542393, 32'sd-0.1875302399326801, 32'sd0.008729161390708798, 32'sd-0.18614686510713482, 32'sd0.2034506003519528, 32'sd0.09417275920492137, 32'sd-0.12953348726735242, 32'sd0.043562237315719676, 32'sd0.23748219938405513, 32'sd-0.003853401495799166, 32'sd0.14163685459742412, 32'sd-0.10186411811294549, 32'sd-0.038858762767161145, 32'sd0.3261813491950103, 32'sd-0.02862436248372179, 32'sd0.004008019312311938, 32'sd-0.175232087694959, 32'sd0.18556544662015187, 32'sd0.21932242105339347, 32'sd-0.14205535706948144, 32'sd-0.17229363426506095, 32'sd0.024783099312892114, 32'sd0.11341648619006325, 32'sd-0.06411733697172729, 32'sd0.01047471196433759, 32'sd-0.11796868537418065, 32'sd-0.1783429203754089, 32'sd-0.06108629338206574, 32'sd-0.03989883032087534, 32'sd0.2032037210290366, 32'sd0.07974495828601927, 32'sd-0.2711586995845133, 32'sd0.014847784377038504, 32'sd-0.1857923473424469, 32'sd-0.25088559239349356, 32'sd-0.07855812214217955, 32'sd-0.019146095719636335, 32'sd0.027968205482194853, 32'sd-0.1956942307096106, 32'sd-0.23186769642304433, 32'sd-0.024168550813233134, 32'sd0.012412039227907287, 32'sd0.006467854511431659, 32'sd-0.194933945865031, 32'sd-0.0985946539395919, 32'sd0.32556300089556867, 32'sd-0.14065011481210316, 32'sd-0.07517857028663857, 32'sd0.11699549758684483, 32'sd-0.2604123766751309, 32'sd0.016002368429043554, 32'sd-0.10831366228789287, 32'sd0.02442395481660683, 32'sd-0.20929081491670945, 32'sd0.26712588212808225, 32'sd-0.11275840675883113, 32'sd-0.1634734214508391, 32'sd0.02228482138135916, 32'sd0.11765945859945287, 32'sd-0.1596403830134944, 32'sd-0.01272491620296051, 32'sd-0.19983333472664935, 32'sd-0.1383980426666628, 32'sd-0.03425649986533683, 32'sd-0.13479307834205503, 32'sd0.11043580371243805, 32'sd-0.0035232346428342855, 32'sd0.2037140936076598, 32'sd-0.16566361400039883, 32'sd0.14973227978173076, 32'sd0.08063157674709648, 32'sd0.19584139568655531, 32'sd-0.11703360576308013, 32'sd0.0014175314115618812, 32'sd-0.24472333682862737, 32'sd-0.005570833521997128, 32'sd0.057274992478476186, 32'sd-0.22202125183517152, 32'sd0.07964215488376213, 32'sd0.09051581003710316, 32'sd-0.016097787078476363, 32'sd0.12320769888248573, 32'sd0.11565991922389485, 32'sd0.02462943269389739, 32'sd0.14411756234513814, 32'sd0.02508985383709004, 32'sd0.11671349710230867, 32'sd0.14244978044249784, 32'sd0.005158746977007444, 32'sd-0.05521091673776943, 32'sd0.12200022097290145, 32'sd-0.1292940686586197, 32'sd0.0158295563026853, 32'sd-0.12692475653610913, 32'sd0.24099261239933695, 32'sd-0.04417891272545226, 32'sd-0.22909848547912584, 32'sd0.1543712165174636, 32'sd-0.0016805745088392906, 32'sd0.0548856736857577, 32'sd-0.23820058109084752, 32'sd0.09558939048843339, 32'sd0.04985218284916546, 32'sd-0.01003458340401389, 32'sd0.09018222939255817, 32'sd-0.1262842648529862, 32'sd0.1326280750287815, 32'sd0.10161522556904626, 32'sd0.03766354728405203, 32'sd0.07894969291852773, 32'sd0.016413866457375872, 32'sd0.15388890862301036, 32'sd-0.09795149053738118, 32'sd0.044015778084434506, 32'sd0.06549331605371661, 32'sd-0.15595198944557287, 32'sd0.10948027441403721, 32'sd-0.003100782349872327, 32'sd0.18325658361263203},
        '{32'sd0.17427776029183709, 32'sd-0.04730366521024956, 32'sd-0.14153798428184405, 32'sd0.0054099722474677155, 32'sd-0.04111473342243913, 32'sd-0.12624723795187767, 32'sd0.13547231336266716, 32'sd0.18427928868569132, 32'sd-0.12199247632016637, 32'sd0.2571644023818198, 32'sd0.13939043213833083, 32'sd0.044280462413046895, 32'sd0.07953462383948466, 32'sd-0.17409287646359223, 32'sd0.022999426728484068, 32'sd0.06025516604522789, 32'sd0.08112919743198195, 32'sd-0.13672676552746355, 32'sd0.04286764679028756, 32'sd-0.18998293519540213, 32'sd0.13109861771674294, 32'sd-0.0919559553686443, 32'sd-0.06550959226189391, 32'sd-0.15481980353586827, 32'sd-0.12208802305468426, 32'sd0.23176719042974675, 32'sd0.0028864787696238695, 32'sd-0.15666082092022407, 32'sd0.06097723448280104, 32'sd0.20475133859621855, 32'sd-0.16794286272965286, 32'sd0.03351820373097354, 32'sd0.29042042300549253, 32'sd0.077813947231125, 32'sd0.1945400552657719, 32'sd-0.1284940033630701, 32'sd-0.0024065184377167585, 32'sd0.022646937095289945, 32'sd0.09999711114760328, 32'sd0.04891279296422555, 32'sd0.07762106473260885, 32'sd-0.28107835512763624, 32'sd-0.09210959716887085, 32'sd-0.10806620459535154, 32'sd-0.27442824321198495, 32'sd0.10061923309669268, 32'sd0.30431278768527426, 32'sd-0.15484884736088314, 32'sd0.14487095373534503, 32'sd-0.055390514661649876, 32'sd0.020120601196286773, 32'sd0.009414305324789396, 32'sd-0.16776409360386083, 32'sd-0.19619808240946296, 32'sd-0.07325709356946931, 32'sd0.05400902196209524, 32'sd0.15317553849967097, 32'sd0.21987559038685187, 32'sd-0.12114669637246911, 32'sd0.003055404772346801, 32'sd-0.10297258012119767, 32'sd-0.19988410172643978, 32'sd-0.007261735381430783, 32'sd0.19132480729261814, 32'sd-0.07026284671675963, 32'sd0.13309340666147135, 32'sd0.07894456076990107, 32'sd0.07735874206093586, 32'sd0.16994592958735583, 32'sd-0.02557985693746206, 32'sd0.20806432889457321, 32'sd0.07399593038653264, 32'sd-0.031421481806911886, 32'sd-0.036430500528750305, 32'sd-0.13886488124329452, 32'sd0.15224457369524869, 32'sd0.1028556595775953, 32'sd0.14365687403106958, 32'sd0.027828014033367758, 32'sd0.08700152598996029, 32'sd0.022444888725190706, 32'sd0.1470378839011447, 32'sd0.06305658346855626, 32'sd0.09590170519926297, 32'sd0.1120300645478333, 32'sd-0.14401675600666278, 32'sd0.04440162912038194, 32'sd0.13291940690514914, 32'sd0.15241985771257727, 32'sd-0.1982915716647499, 32'sd0.027117328223052278, 32'sd0.13522358252583155, 32'sd-0.036907175079300074, 32'sd-0.2235187015327861, 32'sd0.19746511547660547, 32'sd-0.16817786095367382, 32'sd-0.1507473194460933, 32'sd-0.030889470903214734, 32'sd-0.16646166726329448, 32'sd0.14785730152171903, 32'sd-0.17863429534458405, 32'sd-0.00581717279351792, 32'sd0.0761682032145257, 32'sd0.01498135973784299, 32'sd-0.0522889480498049, 32'sd0.21304746816384829, 32'sd-0.02973991596704607, 32'sd-0.09066491521105605, 32'sd-0.07059232775874778, 32'sd0.03274090124167261, 32'sd0.17379986695534005, 32'sd-0.02638603250627813, 32'sd0.11841556628747882, 32'sd0.036940833325852906, 32'sd0.10906867773743043, 32'sd0.13869560947338425, 32'sd0.03869666342393116, 32'sd0.019507855230934883, 32'sd-0.12365422705658555, 32'sd0.012472698141733246, 32'sd-0.190140069633184, 32'sd0.021868332466769357, 32'sd-0.14009840219536254, 32'sd-0.03286734595249763, 32'sd-0.03236768557136613, 32'sd0.1606141063674938, 32'sd-0.16907151713108684, 32'sd0.07310394242877195},
        '{32'sd0.1344062732527156, 32'sd-0.2807265404664669, 32'sd-0.149239789728396, 32'sd-0.04476020382459342, 32'sd-0.21297537615456558, 32'sd0.02065460946910614, 32'sd-0.002692260465915971, 32'sd0.14040489927434266, 32'sd0.012946165835830538, 32'sd-0.1886893945279961, 32'sd0.17912238943443015, 32'sd0.2889316155247691, 32'sd-0.11414732085290374, 32'sd-0.02291862435830981, 32'sd-0.04274166366649112, 32'sd-0.1567968208470461, 32'sd0.06768863771298153, 32'sd0.033699234275384626, 32'sd-0.17701629551559467, 32'sd0.05396587540347072, 32'sd-0.1254572324326435, 32'sd0.22563385199785435, 32'sd-0.04071601258132112, 32'sd0.1857120020813286, 32'sd0.13198447989847106, 32'sd-0.02780030299346581, 32'sd-0.2375030225007118, 32'sd0.01630011791624968, 32'sd-0.02665216154828147, 32'sd0.03839744940892835, 32'sd0.20043028230417234, 32'sd0.21200418071372534, 32'sd-0.3270620406405551, 32'sd0.1380815357818819, 32'sd-0.09262332919173824, 32'sd-0.0576900061704379, 32'sd-0.051150213854605366, 32'sd0.09686721915233776, 32'sd-0.13668815500804976, 32'sd-0.01812008665875239, 32'sd0.019584890851857682, 32'sd0.15511541815165908, 32'sd-0.2763012213532772, 32'sd-0.15422494247051635, 32'sd0.05262067480208087, 32'sd-0.1926783308117408, 32'sd0.08648345000849676, 32'sd-0.28523026791754635, 32'sd-0.19029126930840534, 32'sd-0.11179598187829308, 32'sd0.14722190906419524, 32'sd-0.2957096283544982, 32'sd0.08032926416770646, 32'sd-0.09389690898366385, 32'sd0.018116767486525555, 32'sd-0.05439351289809288, 32'sd-0.043953121286817214, 32'sd0.14669164540015606, 32'sd-0.10823197995422414, 32'sd-0.007091471190994125, 32'sd0.006313790279686311, 32'sd0.18079804938991528, 32'sd-0.01643509134624753, 32'sd0.00905563238891073, 32'sd-0.13594641105730923, 32'sd-0.1440155437561408, 32'sd0.2388045252328544, 32'sd-0.1535845935093721, 32'sd-0.3347291725933474, 32'sd-0.009030669117986025, 32'sd-0.0318409033181796, 32'sd-0.08034997902296312, 32'sd0.20814435104001197, 32'sd-0.05121943678392994, 32'sd0.2801192940929916, 32'sd-0.12192615459851612, 32'sd-0.11510079304733924, 32'sd-0.03960194726032223, 32'sd-0.02014642150535119, 32'sd-0.03872645214158462, 32'sd0.20862915618655417, 32'sd-0.00026901526426692816, 32'sd-0.08181890542113313, 32'sd0.11709273956668342, 32'sd0.12992675769841372, 32'sd0.053882048526999245, 32'sd0.15475792400678604, 32'sd0.008488124992004027, 32'sd0.025883262243795294, 32'sd0.018478848867683074, 32'sd-0.041163509548221504, 32'sd0.1543435489455145, 32'sd-0.2692214734724338, 32'sd-0.07515151118869759, 32'sd0.11655631705377024, 32'sd0.25784551498976205, 32'sd0.32475580186247877, 32'sd0.21719550278333719, 32'sd0.17893891258421665, 32'sd-0.14532048104104295, 32'sd0.038270978183546994, 32'sd-0.05498903075391017, 32'sd-0.3045688594976327, 32'sd-0.16994478805068244, 32'sd-0.2340473466489249, 32'sd-0.07983568327861898, 32'sd-0.0814492125665835, 32'sd0.232751326381849, 32'sd0.029769140778056615, 32'sd-0.008158133266276468, 32'sd-0.16659339157674755, 32'sd0.06731283056685326, 32'sd-0.06226416333514665, 32'sd0.03608791192302576, 32'sd-0.1663405036046435, 32'sd-0.09613082832788014, 32'sd-0.01700226216953005, 32'sd-0.21185437618575353, 32'sd-0.014227072165565473, 32'sd0.1181142829363174, 32'sd0.1564883588001413, 32'sd0.31264852955689515, 32'sd0.13980085732065053, 32'sd0.1177167736231725, 32'sd0.015598491606627091, 32'sd0.207789747234398, 32'sd0.058357019411662346, 32'sd-0.11373395771358981},
        '{32'sd0.03319715986295908, 32'sd-0.0249870148448237, 32'sd-0.1656956979504203, 32'sd0.08496104836823858, 32'sd0.1285839375826741, 32'sd0.005169722594168021, 32'sd0.18100131154866636, 32'sd0.022444926864506342, 32'sd0.1804233841055862, 32'sd-0.063179669160769, 32'sd0.05252889727687598, 32'sd0.16153740591214244, 32'sd0.03221130371920357, 32'sd0.12039633104504277, 32'sd0.06573955790572497, 32'sd-0.11029091301653957, 32'sd-0.17216579153152764, 32'sd-0.09534364544138152, 32'sd0.05797633960783885, 32'sd-0.11725754106483625, 32'sd0.08303834751663007, 32'sd-0.15742556823348203, 32'sd0.04222834053202231, 32'sd0.1332314848246722, 32'sd-0.015153537644505971, 32'sd-0.022754617260733523, 32'sd-0.1366214364720412, 32'sd-0.11978377220186354, 32'sd-0.24113424970167413, 32'sd0.17602302841259765, 32'sd0.11369843470360894, 32'sd0.04208475535242838, 32'sd-0.21480021382027187, 32'sd0.15897418864978194, 32'sd-0.022566342856555295, 32'sd-0.28281235759556356, 32'sd-0.04997548507337088, 32'sd-0.22280958630183914, 32'sd-0.2540033500524764, 32'sd-0.13579320198766714, 32'sd0.053623813660116926, 32'sd0.09109501857575267, 32'sd-0.18894375443845243, 32'sd-0.0009005974788150295, 32'sd0.24363888985788332, 32'sd0.08958437588202298, 32'sd0.043961238740653406, 32'sd-0.1327481511528921, 32'sd0.15102302297180098, 32'sd0.013441986008718975, 32'sd0.19501098814517306, 32'sd-0.04109728185415032, 32'sd-0.01362160876323096, 32'sd-0.17711552542096903, 32'sd0.06792788318380959, 32'sd0.25326588935166267, 32'sd0.0333243146260672, 32'sd0.16287028322261124, 32'sd0.017673786854285202, 32'sd-0.11650096861016017, 32'sd0.0900136624841589, 32'sd-0.10831396370851641, 32'sd0.13897656304269598, 32'sd0.2453365009530888, 32'sd-0.08665286308577645, 32'sd-0.24172605870036135, 32'sd-0.11369181303728595, 32'sd0.08164225133059905, 32'sd-0.2999220539019343, 32'sd-0.007280755695330744, 32'sd0.08134896646087302, 32'sd0.20906101522348106, 32'sd-0.1788996912032405, 32'sd-0.2454454894192372, 32'sd0.04751866112523066, 32'sd-0.08639691762165473, 32'sd-0.22400690005267643, 32'sd0.02111389765772568, 32'sd0.06346480733663491, 32'sd-0.03259969276816138, 32'sd0.003857016724174051, 32'sd-0.22679957489246122, 32'sd-0.00028588405386472174, 32'sd-0.0533000877017824, 32'sd0.08784527224797606, 32'sd-0.20484580472937633, 32'sd-0.020967363317447966, 32'sd-0.11050990694389036, 32'sd0.11448304987969894, 32'sd0.08647723599690474, 32'sd0.21708780573243944, 32'sd-0.04577378554205169, 32'sd-0.23150862173345194, 32'sd0.10657952192018083, 32'sd0.20303686642429314, 32'sd0.031209428582677803, 32'sd0.06250351852126719, 32'sd-0.04230677146260889, 32'sd-0.017400711159039642, 32'sd-0.07655282400188576, 32'sd0.034535713408615214, 32'sd0.1323271500616306, 32'sd0.01872826226260034, 32'sd-0.01156711623130615, 32'sd-0.1321446028985208, 32'sd-0.05852100096086049, 32'sd0.0979035472774862, 32'sd0.08803861722683995, 32'sd-0.08510691978962182, 32'sd-0.17792561623844205, 32'sd-0.16943696855365908, 32'sd0.10872718407865431, 32'sd0.1664745854175826, 32'sd-0.19045380617581617, 32'sd-0.20429710333000023, 32'sd0.07826403655496586, 32'sd0.09182420304275984, 32'sd0.12271652647996471, 32'sd0.10514685626539227, 32'sd0.013264928334801375, 32'sd0.13893436855345018, 32'sd0.13359844385671157, 32'sd-0.08673697786594295, 32'sd-0.10598720894803597, 32'sd-0.01745777018167216, 32'sd-0.13163220361120756, 32'sd-0.1638268307532464, 32'sd0.026875821030738753},
        '{32'sd0.003997760973058812, 32'sd-0.2385881783525356, 32'sd-0.039711466049929714, 32'sd0.23779600863866387, 32'sd0.14994620938698447, 32'sd-0.013680303209889675, 32'sd0.03684217807739801, 32'sd-0.1384272369310956, 32'sd0.15949234900724554, 32'sd-0.0829791795285938, 32'sd0.1669030540044314, 32'sd0.008158654769578296, 32'sd0.2710547351333943, 32'sd-0.163815808276029, 32'sd-0.026325317130666888, 32'sd-0.1391666226322576, 32'sd-0.16767452372691985, 32'sd0.1852544157094373, 32'sd0.06975231973240584, 32'sd0.06012892858152177, 32'sd0.15841602119366816, 32'sd-0.07431439301445841, 32'sd-0.10021074253501067, 32'sd0.0908965482399107, 32'sd-0.06352237361490033, 32'sd-0.11500623257393897, 32'sd-0.0029004621499938263, 32'sd0.033495345270998386, 32'sd-0.051354997282774865, 32'sd0.009616724209669776, 32'sd-0.11364690667564475, 32'sd0.2303389708980729, 32'sd-0.035060248793774375, 32'sd0.11396883521739543, 32'sd-0.12865041895072338, 32'sd0.11671129774539415, 32'sd0.17430540703288783, 32'sd0.09993572951402266, 32'sd-0.09967641078812019, 32'sd0.0897302353798514, 32'sd-0.12396750260173015, 32'sd0.2893762445250082, 32'sd0.09615797016093061, 32'sd0.035019605726625505, 32'sd-0.08249955395337111, 32'sd-0.03883534737396073, 32'sd0.30872360095410145, 32'sd-0.17276490271642198, 32'sd0.009953875501506988, 32'sd0.03500345974037458, 32'sd0.29194468668792223, 32'sd-0.1289578179305301, 32'sd-0.13830037166273054, 32'sd0.03127504062507924, 32'sd0.2288712577115965, 32'sd0.02621924970573503, 32'sd0.15463469175083192, 32'sd-0.15319408559510433, 32'sd-0.2349706925243499, 32'sd0.07796654429579304, 32'sd0.20474345318240356, 32'sd-0.08717935176395407, 32'sd0.09089451393476937, 32'sd0.03594845171750557, 32'sd-0.01962405978714288, 32'sd0.057183710341799227, 32'sd0.08880606912624364, 32'sd0.10650570606340748, 32'sd-0.17383017039279827, 32'sd-0.21787942125867543, 32'sd-0.03080980237267175, 32'sd0.16005931645470256, 32'sd-0.09114185976479748, 32'sd0.21525989693018588, 32'sd-0.15565275604606918, 32'sd-0.08582758760012328, 32'sd0.11153300419332154, 32'sd0.09539858050229626, 32'sd0.110131875872962, 32'sd0.18098699691050874, 32'sd-0.11193349590507987, 32'sd-0.12199761476182487, 32'sd0.0350518781759074, 32'sd-0.0295235422661975, 32'sd0.11481446600017899, 32'sd-0.0325186786975364, 32'sd-0.3630356356712235, 32'sd-0.034231529781677414, 32'sd0.021059181183936713, 32'sd0.13342748724420508, 32'sd0.138906276264849, 32'sd-0.027650665812301356, 32'sd-0.08071797813067993, 32'sd0.1362476247802839, 32'sd-0.09572746084517153, 32'sd-0.12985483850661753, 32'sd-0.1110563617826304, 32'sd-0.07358480784074292, 32'sd-0.2003214423019196, 32'sd-0.003471828789722784, 32'sd-0.13359843685732975, 32'sd0.020422825693345813, 32'sd0.11429006724475975, 32'sd0.19267399506641475, 32'sd-0.12666576325669748, 32'sd0.08884778657449326, 32'sd0.22721875222654792, 32'sd0.21021810433592458, 32'sd-0.10418128635446519, 32'sd-0.16434189258888843, 32'sd-0.0329781489082229, 32'sd0.13357170388686462, 32'sd0.03611447708964321, 32'sd0.11322011829965639, 32'sd0.10935081288716551, 32'sd-0.10728039319897645, 32'sd-0.13217562322852874, 32'sd0.03827922194278158, 32'sd0.18995877613386247, 32'sd-0.039023689343346185, 32'sd-0.08439245620079437, 32'sd-0.16387767432771244, 32'sd-0.029148051306837314, 32'sd-0.08181754585936966, 32'sd0.19989465332939993, 32'sd0.12008197360091105, 32'sd-0.18352435439270015, 32'sd0.26418981192949564},
        '{32'sd0.15466193084152902, 32'sd-0.038657294542217335, 32'sd-0.10866785914644095, 32'sd-0.10289814159315544, 32'sd-0.1400854003519296, 32'sd-0.11226706839455329, 32'sd-0.08420385109208418, 32'sd-0.08778700053496619, 32'sd0.1410859598319578, 32'sd0.1583245482080205, 32'sd-0.05451086555113936, 32'sd-0.06852610653535142, 32'sd0.0987466822131482, 32'sd0.1414353446752335, 32'sd-0.1999718712782384, 32'sd-0.13699471906522132, 32'sd0.12084163498368207, 32'sd-0.0348995652981345, 32'sd0.039072758917431505, 32'sd0.09126939109845784, 32'sd-0.119437822170637, 32'sd-0.11951165009049874, 32'sd0.13604519536531196, 32'sd-0.18818790105709265, 32'sd0.19952165242629433, 32'sd0.26234313252614677, 32'sd-0.09237323484779733, 32'sd0.2050593288171868, 32'sd-0.07745313323085429, 32'sd0.08370226899920447, 32'sd-0.064672118475612, 32'sd-0.08059330754481422, 32'sd-0.055991177415251246, 32'sd0.1017261620607236, 32'sd0.12663791183924983, 32'sd0.08121990123563282, 32'sd0.19966492552439574, 32'sd-0.016582985073768448, 32'sd0.022663627316130638, 32'sd-0.13422637744093538, 32'sd0.1604941892917845, 32'sd-0.07497313882580144, 32'sd0.16284115144281297, 32'sd-0.0035357132501766656, 32'sd-0.14050548254584103, 32'sd0.005615988358840999, 32'sd0.16868078079276294, 32'sd-0.11733588030176081, 32'sd0.06387392499385827, 32'sd-0.17960683141892436, 32'sd0.22558744623640664, 32'sd-0.10924856147475077, 32'sd-0.2056774214130603, 32'sd0.1460976996342364, 32'sd-0.1633360109623518, 32'sd0.23880861212468937, 32'sd0.18512833064462647, 32'sd-0.010437605405314212, 32'sd-0.1729693801723595, 32'sd-0.150663322672929, 32'sd0.1134545378786027, 32'sd-0.034367632292678356, 32'sd0.10114705892468366, 32'sd0.24659236744782212, 32'sd-0.1528387336107561, 32'sd0.021961617138232737, 32'sd-0.019209428063915856, 32'sd0.27895683010175476, 32'sd-0.021016059725384943, 32'sd-0.11857674100555424, 32'sd0.21676457659008078, 32'sd0.11026988950617929, 32'sd0.00041304879325403755, 32'sd0.06506835133083838, 32'sd0.027503896293798152, 32'sd0.20993850153916235, 32'sd-0.049162870461489046, 32'sd0.2952802793778513, 32'sd-0.003137532075605499, 32'sd0.1980867211732877, 32'sd-0.26181366900530906, 32'sd-0.16357925066400755, 32'sd-0.02497979705061576, 32'sd0.04502871198905001, 32'sd-0.045589937003301585, 32'sd-0.1351124651213755, 32'sd-0.294185471725719, 32'sd0.26744123265828224, 32'sd0.03771812174680923, 32'sd-0.16185735100079063, 32'sd0.15448819854849793, 32'sd-0.06502320460997987, 32'sd0.13255932604264026, 32'sd0.005212586371713884, 32'sd-0.1942195576435657, 32'sd0.14518030144699484, 32'sd-0.09484074061588542, 32'sd-0.15568129926010343, 32'sd-0.06848941862171623, 32'sd-0.02294104335128638, 32'sd0.11497725795304747, 32'sd0.20607636724491651, 32'sd0.018875955066276724, 32'sd0.13038616459707905, 32'sd0.09165921064434919, 32'sd0.19859923471565433, 32'sd0.08004457992820528, 32'sd0.09109954320760254, 32'sd-0.07822769835149963, 32'sd-0.05421585121394671, 32'sd-0.08945351576627218, 32'sd-0.2102545409916184, 32'sd0.019769672856265415, 32'sd-0.0025411133940472118, 32'sd0.18169729993164194, 32'sd-0.048623393062150785, 32'sd-0.222072380373704, 32'sd0.024015732458105333, 32'sd0.01211451409492182, 32'sd-0.2366548614174754, 32'sd0.10935018742231739, 32'sd0.07315496627579156, 32'sd0.1602879493901526, 32'sd0.1139875843210631, 32'sd0.22987542155791843, 32'sd-0.1841680653120654, 32'sd-0.2473978894907377, 32'sd-0.04649865009195916},
        '{32'sd-0.08679218703083094, 32'sd-0.3218149159575613, 32'sd-0.1892363723586986, 32'sd0.06600125971689515, 32'sd-0.1738186830334092, 32'sd-0.2031567928485625, 32'sd0.13809070387415118, 32'sd-0.08835270942881719, 32'sd-0.10180811487264456, 32'sd0.028724007541878455, 32'sd0.031037691797652128, 32'sd-0.18481117891187182, 32'sd0.17001258819904747, 32'sd-0.13489992175697263, 32'sd0.08164330615165177, 32'sd0.0432793936730288, 32'sd0.004104799907066397, 32'sd-0.18947905904708298, 32'sd0.1617594630401737, 32'sd-0.13393145857112732, 32'sd-0.13076636901523134, 32'sd-0.06422438894572663, 32'sd0.14235338279933088, 32'sd0.04102329012185829, 32'sd-0.1616787993178984, 32'sd0.016527380184062253, 32'sd0.16284799604609018, 32'sd-0.03786911708533535, 32'sd-0.1408081478019141, 32'sd0.011581342167334092, 32'sd0.08728588220211722, 32'sd-0.0804022108389328, 32'sd-0.0022959990415363433, 32'sd0.2408549128899696, 32'sd-0.06818601126069855, 32'sd0.02966281130817754, 32'sd0.0967260298798828, 32'sd0.16752864483818228, 32'sd0.17544104389651685, 32'sd0.060246616456828744, 32'sd-0.23234360649644226, 32'sd0.1738044972750159, 32'sd-0.1328595868729051, 32'sd-0.1690982922642479, 32'sd-0.09841125699555833, 32'sd0.18510028786836874, 32'sd0.036874471170249806, 32'sd-0.21271630802504138, 32'sd-0.29160427006677164, 32'sd4.827597389318026e-06, 32'sd0.09169664538562455, 32'sd0.19857741221207603, 32'sd-0.08600011007817311, 32'sd0.1352434509305901, 32'sd0.05377120240743788, 32'sd0.12277455051473073, 32'sd0.05789442580286315, 32'sd-0.08121879643553956, 32'sd-0.10458837067264734, 32'sd0.1236294578495571, 32'sd0.04221230242699225, 32'sd-0.016762323957819254, 32'sd-0.07672796792382885, 32'sd-0.01747632341195648, 32'sd0.08563729124920404, 32'sd0.1695566387697578, 32'sd0.08447599234028653, 32'sd-0.01142596500233442, 32'sd-0.21421902026588188, 32'sd0.12619893822224315, 32'sd-0.12423518512595653, 32'sd0.08524556098456951, 32'sd0.14457140531269197, 32'sd0.19957337664935743, 32'sd-0.14934331927448397, 32'sd-0.27539740472901253, 32'sd0.07754913061055536, 32'sd0.021913906884894495, 32'sd0.03404912547365202, 32'sd0.1679936635455524, 32'sd-0.09215656064460377, 32'sd-0.23705967923306762, 32'sd-0.15211872614738006, 32'sd0.1200846641911072, 32'sd-0.06271245717254595, 32'sd-0.05066356194247324, 32'sd0.20817618891643586, 32'sd0.008639511842444818, 32'sd-0.03404691816921676, 32'sd-0.04359444336335733, 32'sd0.2085436206084848, 32'sd0.20415909178893896, 32'sd0.07522808455966096, 32'sd-0.02758405468300828, 32'sd-0.10147340887320906, 32'sd0.12865724459200595, 32'sd-0.19088557761697533, 32'sd-0.12440743723526872, 32'sd-0.03330388588428059, 32'sd-0.10173737359954907, 32'sd-0.1278734302406381, 32'sd-0.006663796787395241, 32'sd0.1961596988152304, 32'sd-0.14605270305575477, 32'sd0.07323460000970589, 32'sd-0.38224038226505697, 32'sd0.09584865150548061, 32'sd0.141002891634121, 32'sd-0.017245181703793553, 32'sd-0.0023559937261692166, 32'sd0.01574298101423646, 32'sd0.1277675534532548, 32'sd0.028522542026596265, 32'sd0.03916873207438904, 32'sd-0.06318969133352435, 32'sd-0.09998286779494193, 32'sd0.17613594696110202, 32'sd-0.06305394946727266, 32'sd-0.018739270566249897, 32'sd-0.012333716230033286, 32'sd0.22372375337816122, 32'sd-0.06418638239715378, 32'sd0.02945841762278687, 32'sd0.12381999506551566, 32'sd0.05350695648907752, 32'sd0.12906598481099657, 32'sd-0.11458360114557545, 32'sd0.14099671489705234},
        '{32'sd-0.016636507481339206, 32'sd-0.04633524279689837, 32'sd0.021810219965829204, 32'sd-0.08348182287765679, 32'sd-0.13283590373952425, 32'sd0.0936641123991048, 32'sd-0.06880101613785854, 32'sd0.20691695081174402, 32'sd0.05393447161785732, 32'sd-0.13061103681509978, 32'sd0.04674565687775391, 32'sd0.017093902355335394, 32'sd0.08249236184373022, 32'sd-0.14868495526651956, 32'sd-0.24422214839672476, 32'sd0.014262666591085138, 32'sd-0.1419489908214194, 32'sd0.14662600102934797, 32'sd0.01947716665188046, 32'sd-0.18751788597214764, 32'sd0.0009605573007942909, 32'sd-0.022328652032553693, 32'sd-0.11089726453801263, 32'sd-0.16304990259567329, 32'sd0.20119534214788662, 32'sd0.13000817431067166, 32'sd-0.06902103360721872, 32'sd0.1411402658262089, 32'sd-0.1057502265876063, 32'sd-0.00453559033686577, 32'sd-0.2156568955175056, 32'sd0.22123590036090088, 32'sd0.027734978870627255, 32'sd-0.05084121743436033, 32'sd0.01921836316148364, 32'sd0.04486435051817433, 32'sd-0.05935554915730559, 32'sd0.14403860978669428, 32'sd0.1307762666894679, 32'sd-0.14973462370556823, 32'sd0.14057316014209642, 32'sd0.022417936648673347, 32'sd-0.1426903967442653, 32'sd-0.21698944879868085, 32'sd0.069829023944445, 32'sd-0.19579822610314718, 32'sd-0.167183722106913, 32'sd0.10874861278990676, 32'sd0.08365984473363518, 32'sd-0.020602654653172552, 32'sd-0.1259669090167919, 32'sd0.16081578346088557, 32'sd-0.13440516172419215, 32'sd0.12472527290006793, 32'sd0.022906536515554566, 32'sd0.03580962524205443, 32'sd-0.2202916704392171, 32'sd-0.21693118555123, 32'sd-0.016172632616893553, 32'sd-0.1170701715882897, 32'sd-0.01429122192972885, 32'sd0.20271650892017312, 32'sd-0.1216192595277624, 32'sd-0.05177061710900441, 32'sd0.00651258595917468, 32'sd0.16379065649397195, 32'sd0.22335852096392841, 32'sd0.02923991677597809, 32'sd-0.06650720334610569, 32'sd0.0906096751529754, 32'sd-0.04460186532049124, 32'sd-0.03534527472884239, 32'sd-0.001224285588635893, 32'sd0.13416480789916357, 32'sd-0.07936619838212487, 32'sd0.03048294926762162, 32'sd0.12887685165035223, 32'sd-0.012115481422482534, 32'sd-0.008241404956363075, 32'sd-0.12957921512248508, 32'sd0.1238936756763765, 32'sd0.1554791597600114, 32'sd0.003724179095693642, 32'sd-0.03382248672692214, 32'sd-0.27044630561474664, 32'sd0.19059861803183983, 32'sd-0.15085213575874562, 32'sd0.2103940054597304, 32'sd0.07612846410906858, 32'sd0.020563791992130123, 32'sd0.07666681881019911, 32'sd0.08484280816225552, 32'sd-0.07330920777983288, 32'sd0.23286955259062966, 32'sd0.04194131486714543, 32'sd0.020389663224990105, 32'sd-0.02140217584632533, 32'sd0.05107879294387051, 32'sd-0.18684771660590982, 32'sd0.1235635957043746, 32'sd0.11632969085540397, 32'sd0.1322598341680441, 32'sd0.024574753067680356, 32'sd-0.0005392558042160326, 32'sd-0.2007964072738052, 32'sd-0.035783233528406164, 32'sd0.0730429314719996, 32'sd0.08968498232303239, 32'sd0.10775331542263292, 32'sd0.041241762795751105, 32'sd-0.28547315944258783, 32'sd0.07313404176771325, 32'sd-0.054227414521937425, 32'sd0.007198530843829299, 32'sd0.1474327673299957, 32'sd0.010792644394978313, 32'sd-0.08963431493176854, 32'sd-0.12492063912281143, 32'sd-0.017503064257877444, 32'sd-0.11977495942206487, 32'sd-0.11798697653017569, 32'sd0.09040898548769535, 32'sd0.18080010208735814, 32'sd0.19074488995806463, 32'sd-0.07444579110656405, 32'sd0.21536615116105173, 32'sd-0.07596346410891601, 32'sd0.0021148339606450292},
        '{32'sd-0.22072355006933164, 32'sd0.03063007139992219, 32'sd0.03996022013466825, 32'sd0.024937698828081948, 32'sd-0.14477996446735641, 32'sd0.07719600364814347, 32'sd0.21407957498851626, 32'sd0.12496644482603844, 32'sd0.12400274574942717, 32'sd-0.005962962493282746, 32'sd0.1293434912340724, 32'sd-0.07442958858191481, 32'sd0.043399025019893185, 32'sd0.05879214722099536, 32'sd0.022988169115871423, 32'sd0.18739740555783027, 32'sd0.03627337225646896, 32'sd-0.2431104947342569, 32'sd0.01478659298921751, 32'sd0.022768831077419144, 32'sd-0.017103443471147887, 32'sd-0.1925514094422687, 32'sd-0.2770008037518238, 32'sd0.14809384111501261, 32'sd-0.0281553120308806, 32'sd-0.004174957069727683, 32'sd-0.13762031760088303, 32'sd-0.005069032321532831, 32'sd-0.015481249888078901, 32'sd0.15167010619179352, 32'sd0.19412482382675575, 32'sd-0.06003866448010182, 32'sd-0.07962867394800444, 32'sd0.0888143434908902, 32'sd-0.06605794385829813, 32'sd-0.048982083347244854, 32'sd0.05815301311066872, 32'sd-0.11345218468625251, 32'sd0.19404240377238743, 32'sd0.13236425849832634, 32'sd0.07818031486972161, 32'sd-0.18763260949314914, 32'sd0.22625878888333267, 32'sd0.04438080693071635, 32'sd0.0785262138425694, 32'sd0.14832757133616167, 32'sd0.2548883933683947, 32'sd0.039936760065422676, 32'sd0.19902883068757238, 32'sd0.044305700947205935, 32'sd0.025942005256727164, 32'sd-0.17673581495689777, 32'sd0.02379574117734792, 32'sd-0.2483642148698798, 32'sd0.026334175035864844, 32'sd-0.02776249390709588, 32'sd-0.1311457330208745, 32'sd-0.20126169848223652, 32'sd-0.07709914281841652, 32'sd-0.11168929583518585, 32'sd0.14678552179758214, 32'sd-0.0910173922103542, 32'sd-0.16379199372261163, 32'sd0.11146989332540462, 32'sd0.026247033849810617, 32'sd-0.009260625817160919, 32'sd0.06140725435904536, 32'sd0.09432931432829242, 32'sd0.04049464732077002, 32'sd0.17190520582604502, 32'sd-0.23778041885080714, 32'sd-0.06721303530729553, 32'sd0.1876240154848762, 32'sd0.08974531528549487, 32'sd-0.16619527240138457, 32'sd0.17978200481497483, 32'sd0.13909602501209622, 32'sd0.16934980683536108, 32'sd0.18039774186964294, 32'sd-0.2643139635535237, 32'sd-0.030208875896929586, 32'sd0.06777959984323557, 32'sd0.07384081890223666, 32'sd-0.03283421073348796, 32'sd0.16417426775836677, 32'sd-0.05899520075347552, 32'sd-0.00871261844225818, 32'sd-0.23498228699693768, 32'sd0.1724845621301364, 32'sd0.2176300343918476, 32'sd0.12593597406817614, 32'sd0.22959980797542848, 32'sd0.0869728408901416, 32'sd-0.1481962310707547, 32'sd0.18314301262795674, 32'sd-0.27731816577730917, 32'sd-0.13525515026212726, 32'sd-0.01642493247608684, 32'sd-0.12811807538102557, 32'sd0.11745778455488999, 32'sd-0.10579139214540767, 32'sd-0.12824038121971165, 32'sd0.05831527021904912, 32'sd-0.1647812756585539, 32'sd0.05072251973885085, 32'sd-0.14200627253922776, 32'sd0.06213288976642456, 32'sd-0.06726265886975102, 32'sd0.14062034719607253, 32'sd-0.12445496344371364, 32'sd-0.06828013404753665, 32'sd0.11177613438594643, 32'sd-0.19044111471785805, 32'sd0.026137224646658262, 32'sd-0.01956623579094946, 32'sd0.2625870412140608, 32'sd-0.09405154717059282, 32'sd0.15799021481466244, 32'sd-0.23816835170458647, 32'sd0.25648186824372515, 32'sd-0.20052602615320705, 32'sd-0.08440231052332575, 32'sd0.15203087025526238, 32'sd-0.090601498445812, 32'sd-0.11631983664974563, 32'sd-0.3201891667979139, 32'sd0.18334065351508924, 32'sd0.223673620373357},
        '{32'sd-0.15687413641467315, 32'sd0.1716683105038971, 32'sd-0.2821262073637795, 32'sd0.1687575111290954, 32'sd0.00011944353008413235, 32'sd-0.1482428902122782, 32'sd-0.13282241827439076, 32'sd0.09821727779949684, 32'sd-0.06887583007097163, 32'sd-0.22038319151960725, 32'sd-0.04494464612633592, 32'sd0.0458409114067568, 32'sd0.0748245771745071, 32'sd-0.08549560006500778, 32'sd-0.052469683183512965, 32'sd-0.005589823057534229, 32'sd0.12856364492618721, 32'sd0.03287202137639879, 32'sd-0.159933412488862, 32'sd-0.09182046737759429, 32'sd-0.06774850642578545, 32'sd-0.029816443376298244, 32'sd-0.29177980427054406, 32'sd-0.04499266453306565, 32'sd-0.0922764750412707, 32'sd0.165790554196379, 32'sd0.17871916404023228, 32'sd-0.14226170651121997, 32'sd-0.16322737900704626, 32'sd0.27074596115270533, 32'sd-0.04006216268852176, 32'sd-0.14487814817750005, 32'sd-0.10198186876303225, 32'sd0.030512544855206478, 32'sd0.016142910954334445, 32'sd-0.0845254209967076, 32'sd0.047970314762149545, 32'sd0.1271404966620138, 32'sd-0.18028484079944398, 32'sd0.11462283719412113, 32'sd-0.09599762607914372, 32'sd0.14200825044690954, 32'sd0.10904932926589524, 32'sd-0.17614690858302243, 32'sd-0.15169396810234106, 32'sd0.12645931081474773, 32'sd0.21588329249199037, 32'sd0.19920232445152336, 32'sd0.02165691699320026, 32'sd0.0730480626352739, 32'sd0.24841030688547464, 32'sd-0.036267002230994175, 32'sd-0.021857237689357656, 32'sd-0.07345291997232029, 32'sd-0.1210980960294639, 32'sd-0.13133396360459765, 32'sd-0.10909240032476768, 32'sd-0.00012539261871766184, 32'sd0.0630269430954957, 32'sd0.0643529264020495, 32'sd0.14089116851054748, 32'sd-0.08727584097889987, 32'sd0.2574639539879219, 32'sd0.0480758239914688, 32'sd-0.22724598816336872, 32'sd-0.09847298600579765, 32'sd0.2634755704146238, 32'sd0.16956344762592196, 32'sd0.01938721384143976, 32'sd0.0373239582301266, 32'sd-0.15997081546659714, 32'sd-0.3195377809568443, 32'sd-0.1320633590876512, 32'sd-0.17324895156039535, 32'sd0.12551509387218895, 32'sd0.2674577906685584, 32'sd0.23604878595580225, 32'sd-0.0986390905206508, 32'sd-0.12099860496791824, 32'sd-0.016621141490508525, 32'sd0.26981111034037564, 32'sd0.03533437725313455, 32'sd0.04692486035693594, 32'sd0.04393459451450639, 32'sd0.033693034252018056, 32'sd-0.08646081615764463, 32'sd-0.04306844579779664, 32'sd0.12000325713115717, 32'sd-0.12924201897433904, 32'sd-0.23151601505409064, 32'sd-0.061200864262995834, 32'sd0.024726327174255897, 32'sd-0.05173680455925406, 32'sd-0.16101823777890076, 32'sd-0.25376124580865567, 32'sd-0.11256518417858777, 32'sd0.0875581081025133, 32'sd0.19571016321351628, 32'sd-0.05853334485067712, 32'sd0.08111674461765561, 32'sd-0.10570856462087588, 32'sd0.1717072469086274, 32'sd0.06771451668137779, 32'sd-0.10822417873512576, 32'sd-0.28347575369559913, 32'sd0.005052050887069204, 32'sd-0.02304078475236996, 32'sd0.030276937034911234, 32'sd-0.1633791516748131, 32'sd0.14030218379341486, 32'sd0.05274027744443807, 32'sd0.17097811922021572, 32'sd0.261262519611406, 32'sd-0.0064994587839434246, 32'sd-0.012502458657646863, 32'sd0.026136033455676957, 32'sd0.07690392883792341, 32'sd-0.13161657780105826, 32'sd0.17645932585252544, 32'sd0.10168750671921088, 32'sd-0.0879163528670056, 32'sd-0.07850668069875816, 32'sd-0.16789525149469042, 32'sd-0.16514805704891933, 32'sd-0.22840361994027847, 32'sd0.050373221544291885, 32'sd0.11845276274978832, 32'sd-0.1060346311567523},
        '{32'sd-0.20459805547621673, 32'sd0.03686809285436891, 32'sd-0.03983317402008428, 32'sd0.013310174049742917, 32'sd0.2064778902802806, 32'sd0.18571394575835112, 32'sd-0.20370615976774345, 32'sd0.17396006506896036, 32'sd-0.08399228199507953, 32'sd0.0014612239243658933, 32'sd0.017516150580407102, 32'sd0.023870204352282598, 32'sd0.03614034425698562, 32'sd-0.031474367642616644, 32'sd-0.08085425285320827, 32'sd0.14279952928152945, 32'sd0.15759435692266394, 32'sd-0.11147606031175485, 32'sd-0.18586128943943886, 32'sd0.02399224054891829, 32'sd0.08216785353351909, 32'sd0.021858693889512747, 32'sd0.09460324024070574, 32'sd0.16664924362204828, 32'sd0.15377439886642308, 32'sd0.16021446441748743, 32'sd0.16034877557402544, 32'sd-0.06545630368620764, 32'sd0.07040087198627949, 32'sd-0.19967435857773466, 32'sd-0.27044488255270044, 32'sd-0.11226782922292286, 32'sd-0.0006908363534758546, 32'sd-0.19781154985721547, 32'sd-0.0013109181881145737, 32'sd0.13106217030081374, 32'sd0.0019402894479556424, 32'sd-0.07982337481446042, 32'sd-0.0052451451291401505, 32'sd0.18902167037536677, 32'sd-0.0585527916698931, 32'sd0.07453984871254686, 32'sd-0.08548319432606868, 32'sd-0.18883159642516376, 32'sd-0.11096262245899435, 32'sd0.01241715232515298, 32'sd0.1973736142943307, 32'sd0.08507753392603971, 32'sd-0.16667591538662244, 32'sd0.05304906733670193, 32'sd0.05350974291651983, 32'sd0.1921042673512485, 32'sd-0.2630743327377476, 32'sd0.1739141058291024, 32'sd-0.2587700286440895, 32'sd-0.0698566298118272, 32'sd-0.12452799422740254, 32'sd-0.047938860301748355, 32'sd-0.04114541237662392, 32'sd-0.07107621270827934, 32'sd0.24099947823139153, 32'sd0.04587035612870187, 32'sd0.03600022558638028, 32'sd0.1991530687204354, 32'sd0.08836248378411182, 32'sd0.23772542568784122, 32'sd-0.1308595814800292, 32'sd-0.03140523662751128, 32'sd0.019887599279893708, 32'sd-0.23966377361379063, 32'sd0.22393450570665985, 32'sd0.012976392863248193, 32'sd-0.10744922905167198, 32'sd0.15428023004619773, 32'sd-0.33259122370207017, 32'sd-0.1592377435707381, 32'sd-0.12836244652932785, 32'sd0.010827849883337596, 32'sd0.17470706210450246, 32'sd-0.033635345862919316, 32'sd-0.1504108689849499, 32'sd0.035926610171642906, 32'sd0.175842787460699, 32'sd-0.02366402935094129, 32'sd-0.0030517382319928607, 32'sd-0.2867473866546143, 32'sd0.002543047686006723, 32'sd-0.030548206137845018, 32'sd0.07886330713025448, 32'sd-0.05888963222317233, 32'sd-0.12789010796812758, 32'sd-0.17016781426208788, 32'sd0.029259115738778565, 32'sd-0.04005154727878438, 32'sd0.07586144624342403, 32'sd0.06802335515614422, 32'sd-0.24231578355880337, 32'sd-0.06388010519442963, 32'sd0.1367341229796265, 32'sd-0.028566578466872133, 32'sd-0.08594008545751186, 32'sd-0.11856443317123595, 32'sd0.22130766427202278, 32'sd-0.17923172295035733, 32'sd-0.04618164884726324, 32'sd-0.19162192044493445, 32'sd0.17982984233755578, 32'sd-0.02264218319845754, 32'sd0.031614362995678005, 32'sd-0.11611584726177164, 32'sd0.016281719929007916, 32'sd0.006913720933607551, 32'sd-0.12832115050724005, 32'sd-0.09746104776703961, 32'sd0.10552133351028475, 32'sd0.2173529086263801, 32'sd-0.1434331094259635, 32'sd-0.11395866238797778, 32'sd0.1366145440075855, 32'sd-0.1022852252968789, 32'sd0.11856839794747497, 32'sd-0.14391751743328993, 32'sd0.09746082910315097, 32'sd-0.16849516706768713, 32'sd0.10556158281353542, 32'sd0.09046812295205849, 32'sd-0.06195935441441833, 32'sd-0.01289704527315687},
        '{32'sd0.023354934046391856, 32'sd-0.16547612512294768, 32'sd-0.24365796915754295, 32'sd0.22860360293856147, 32'sd0.14088807099673456, 32'sd0.16404497908362614, 32'sd-0.0767331695674038, 32'sd0.12883709901183815, 32'sd-0.0649037762200725, 32'sd0.0780974154606826, 32'sd0.14250242611819355, 32'sd0.20235431968825163, 32'sd0.06487592684271132, 32'sd-0.020871086312460947, 32'sd-0.053309024620040106, 32'sd-0.19807486967825114, 32'sd-0.08090479913484908, 32'sd-0.1120261243582066, 32'sd-0.027460257603908023, 32'sd-0.11683068860921557, 32'sd-0.10691844932840913, 32'sd0.12705630227119658, 32'sd-0.24302928090721754, 32'sd-0.02338007482041414, 32'sd-0.03994901670113094, 32'sd0.18992084209203727, 32'sd-0.27312408451670706, 32'sd0.02404317589140097, 32'sd0.0944286136357898, 32'sd0.12678745167567107, 32'sd-0.02508048062915415, 32'sd0.008011968806426652, 32'sd-0.20973890675271348, 32'sd-0.01502044781753129, 32'sd0.11412199015638101, 32'sd0.0023857710003154487, 32'sd0.06094214948584991, 32'sd0.07161190204221389, 32'sd-0.28962823582465097, 32'sd-0.11746585499342808, 32'sd0.28679809534930023, 32'sd0.08976259540646327, 32'sd0.10471835627615832, 32'sd0.16127857464580772, 32'sd0.17692908926985826, 32'sd-0.15194507141079736, 32'sd-0.03573716425967286, 32'sd-0.027751251819632967, 32'sd0.005128702862101022, 32'sd-0.15799060767867848, 32'sd0.2116085925942215, 32'sd0.05389437789777536, 32'sd0.09976214315812212, 32'sd0.16601166714550128, 32'sd0.22115160836062786, 32'sd0.041571392488109114, 32'sd-0.13364828730152117, 32'sd0.14028770744862482, 32'sd-0.06887735687321052, 32'sd0.058971144227095804, 32'sd0.16132532464476199, 32'sd0.08144428955910266, 32'sd-0.0034293684377986232, 32'sd0.13669396281332677, 32'sd0.02711512157303165, 32'sd-0.23278063096718793, 32'sd0.050094425158296624, 32'sd0.10138044259458873, 32'sd-0.2234516222790647, 32'sd0.09204127313121438, 32'sd0.021426375221990694, 32'sd0.20378155190657, 32'sd0.06965460937098335, 32'sd-0.10454631809721922, 32'sd0.20581239738415727, 32'sd0.2023894443761455, 32'sd0.019306396975601624, 32'sd-0.09548505674247112, 32'sd0.17859554436134104, 32'sd0.11390787171584026, 32'sd-0.08168465156692178, 32'sd-0.14604028222177676, 32'sd0.06763742611888088, 32'sd-0.04617859293378375, 32'sd0.18909353466202186, 32'sd-0.1848206708752074, 32'sd0.05070520103192055, 32'sd-0.04860748123725151, 32'sd0.10997626763752776, 32'sd-0.053606286611297564, 32'sd0.028205259279537327, 32'sd0.15657222113274147, 32'sd0.014877934133409182, 32'sd0.17135562385956918, 32'sd0.008423889141561332, 32'sd-0.13174582896655535, 32'sd0.03960143411534101, 32'sd0.2231717435170918, 32'sd-0.13570322640709925, 32'sd0.09007064360313119, 32'sd0.006684922746216748, 32'sd-0.06271100369715908, 32'sd-0.17815660348219536, 32'sd0.07222176995297276, 32'sd-0.07366875042084839, 32'sd-0.10150858258958058, 32'sd0.032078414666994605, 32'sd0.0890651003266496, 32'sd-0.1388318958882096, 32'sd0.14340710470578974, 32'sd-0.23189974329650556, 32'sd0.027656772959539368, 32'sd0.08133206895543532, 32'sd0.0036646650601933088, 32'sd0.08093436089747778, 32'sd0.06740269916356308, 32'sd-0.15757446381271442, 32'sd0.016651554798380735, 32'sd0.17307574878795767, 32'sd-0.2847857399648499, 32'sd0.23922201698008788, 32'sd0.05275786708790555, 32'sd-0.0008305068478419769, 32'sd-0.06184773988033394, 32'sd0.19846893312934635, 32'sd0.11331474141349787, 32'sd-0.05441392768471086, 32'sd0.23229143254404128},
        '{32'sd0.19957882070448513, 32'sd0.188573958799683, 32'sd0.018292789616168065, 32'sd-0.10631259173114972, 32'sd-0.2335971958573098, 32'sd-0.028324512802442442, 32'sd0.08956046643686977, 32'sd0.17429918088449886, 32'sd-0.19567803169506265, 32'sd0.09517670758234659, 32'sd-0.13571738720585777, 32'sd0.03181965011531294, 32'sd-0.03930585939527679, 32'sd0.09403806595959542, 32'sd-0.13115211732931442, 32'sd-0.21211029559607494, 32'sd0.22247833014397814, 32'sd-0.1435471987420549, 32'sd0.07104546194482352, 32'sd0.043979245905681585, 32'sd-0.07502566751615772, 32'sd-0.050278373500956826, 32'sd0.1590828987943834, 32'sd0.0877891502193956, 32'sd0.10388347334138018, 32'sd0.20892885902416808, 32'sd-0.09509226176344597, 32'sd-0.00242769692206774, 32'sd-0.033587835740963655, 32'sd0.1264342295841027, 32'sd-0.1350650125267338, 32'sd-0.17526453808078993, 32'sd0.07069424855030015, 32'sd-0.09333850527930507, 32'sd0.03175028089340656, 32'sd-0.07989390590670141, 32'sd0.20471221246194643, 32'sd-0.08157584655904589, 32'sd0.05183466518190193, 32'sd0.07908061249325125, 32'sd0.14014981890955452, 32'sd0.09312566230862093, 32'sd0.05955185144201261, 32'sd0.1676186657112304, 32'sd-0.22943245108739857, 32'sd-0.007305718643546213, 32'sd-0.02850465795469988, 32'sd-0.012870845286029954, 32'sd-0.04318989005357899, 32'sd-0.10419758735276596, 32'sd0.1581068498057455, 32'sd0.07605633338854645, 32'sd0.007745432559767992, 32'sd0.06126554445571624, 32'sd-0.16725201187396638, 32'sd-0.13913211001635084, 32'sd0.21582454001472673, 32'sd0.0073706561790613115, 32'sd-0.20710876828782418, 32'sd0.11931787971088685, 32'sd0.141570181568889, 32'sd0.005488501433230094, 32'sd0.08761417734810054, 32'sd0.12260570152964959, 32'sd0.06275537009060529, 32'sd-0.1362120779708451, 32'sd-0.022357047052908915, 32'sd-0.09076744960182992, 32'sd0.15854836101260752, 32'sd-0.0402675073094199, 32'sd0.1882175731488963, 32'sd0.018760766857943607, 32'sd0.06459201073407032, 32'sd0.20394241548397676, 32'sd-0.24917782007416395, 32'sd0.17215513197987647, 32'sd-0.1354218196803868, 32'sd-0.04224469739223546, 32'sd0.09055587139509291, 32'sd0.06563765707193613, 32'sd0.024235665700770074, 32'sd0.0737964807129064, 32'sd0.1984943738837591, 32'sd0.09924951762972443, 32'sd-0.07814053493233591, 32'sd0.2132453689645352, 32'sd0.041361829183932323, 32'sd0.1883983338236044, 32'sd0.25822944203401366, 32'sd-0.17171623713830855, 32'sd-0.1778729741547792, 32'sd-0.04699182313327886, 32'sd-0.06803648247428627, 32'sd0.04756816809263584, 32'sd-0.12475802097029821, 32'sd-0.1603164555288956, 32'sd-0.05925454435906845, 32'sd-0.18384091517143458, 32'sd0.23717285354022913, 32'sd0.021230602558234085, 32'sd0.15949532068959604, 32'sd0.15552020387643897, 32'sd-0.10286523170428717, 32'sd-0.05110073479533353, 32'sd-0.036676199123150864, 32'sd0.14310982381666842, 32'sd0.19722356896671997, 32'sd-0.09625552712029142, 32'sd-0.17317829047374814, 32'sd0.1959954955436475, 32'sd0.15594275531947063, 32'sd-0.1625218343775577, 32'sd0.042119152972885536, 32'sd0.26949350638185093, 32'sd0.012350989097385285, 32'sd0.07378253924206334, 32'sd0.055020586991307095, 32'sd0.045158115912044425, 32'sd0.021188946094376822, 32'sd0.22717508373226905, 32'sd-0.049904670198718734, 32'sd-0.24967031538073786, 32'sd-0.0855505562053657, 32'sd0.03569228258535158, 32'sd0.1035837380897336, 32'sd0.1081588693672126, 32'sd-0.05082386271941911, 32'sd-0.11972151596949648},
        '{32'sd0.04489204008821181, 32'sd0.06321153329132925, 32'sd0.036814767535486154, 32'sd0.15149644763989983, 32'sd0.04119239276134772, 32'sd-0.15800736573247898, 32'sd0.1408176292586471, 32'sd-0.22119141769098197, 32'sd0.11460979980064055, 32'sd-0.015869575196320856, 32'sd-0.17758457188975466, 32'sd-0.07882790951747272, 32'sd-0.17155673453890327, 32'sd-0.23367230666069266, 32'sd0.24034034657103545, 32'sd0.007203052169612635, 32'sd0.10156195244473369, 32'sd0.05053009932338358, 32'sd-0.08435958561449934, 32'sd0.03627391165912896, 32'sd0.10834783574715898, 32'sd-0.17797941738906775, 32'sd0.04037489278287394, 32'sd0.1352101527359879, 32'sd0.08260568407884926, 32'sd-0.007687060026101563, 32'sd-0.1467289781919873, 32'sd-0.10234340884092936, 32'sd0.04244685058150538, 32'sd0.19030791114963366, 32'sd-0.11819801392685729, 32'sd-0.2532800705382981, 32'sd0.17048625721374983, 32'sd0.1645338571037118, 32'sd0.15854163240705615, 32'sd0.01870638094079028, 32'sd0.07819100045658586, 32'sd-0.03436583472482865, 32'sd-0.0628535244371508, 32'sd-0.14558877662824685, 32'sd-0.18399432999517212, 32'sd-0.08389020877695165, 32'sd0.033982235949948876, 32'sd0.14175758560752616, 32'sd-0.03878699034292576, 32'sd-0.12404374943837898, 32'sd0.1794985048476441, 32'sd-0.18713697368795165, 32'sd0.12218742138307433, 32'sd0.1449215802455263, 32'sd-0.10125176452524468, 32'sd-0.1365687507153109, 32'sd0.09459153495369846, 32'sd0.10941048416877476, 32'sd-0.2306963614952352, 32'sd-0.1561122013273054, 32'sd0.17287158577579873, 32'sd-0.15468767128945857, 32'sd0.05981334230589349, 32'sd-0.18731619337245142, 32'sd0.2737053778691333, 32'sd0.02083962723098283, 32'sd-0.24315904049408965, 32'sd0.0957404526653762, 32'sd-0.04155383969580856, 32'sd-0.04351017885043817, 32'sd0.050731383439245006, 32'sd0.08076312732277147, 32'sd0.14371588397474683, 32'sd0.02328153706624373, 32'sd-0.15247409055376568, 32'sd0.01915200974057291, 32'sd0.10399642817326897, 32'sd0.1811720727156482, 32'sd-0.27555844593566686, 32'sd-0.07835735255143293, 32'sd0.10584869207402836, 32'sd-0.03987021448109773, 32'sd0.12635610736567665, 32'sd0.16536434799312455, 32'sd0.07482679187857413, 32'sd-0.10538564790666881, 32'sd0.10140553450841114, 32'sd-0.12029085625334439, 32'sd0.08619700304713214, 32'sd0.10165002985507542, 32'sd0.0006110460624616766, 32'sd-0.09028277411048215, 32'sd0.16785065027214843, 32'sd0.2953820724397227, 32'sd0.12810531864979902, 32'sd0.21030300453373102, 32'sd0.19233003654140074, 32'sd-0.07005456886126257, 32'sd0.18836579935904754, 32'sd-0.2031973417352104, 32'sd-0.05370864805161598, 32'sd-0.2580417872252115, 32'sd-0.058688121372475, 32'sd-0.032658426115362044, 32'sd0.04053611361020106, 32'sd-0.10631092088936325, 32'sd0.16853541701786956, 32'sd-0.0027762478341145105, 32'sd0.1660873470086815, 32'sd0.015731707522738565, 32'sd0.1605871785018592, 32'sd-0.1559993366539345, 32'sd0.04650626330984964, 32'sd-0.0919879823404852, 32'sd0.11995987277686604, 32'sd-0.1746609139172506, 32'sd-0.32662540847425997, 32'sd0.035004009530335736, 32'sd0.18627778740407286, 32'sd0.05951062884324996, 32'sd-0.21406702281756387, 32'sd0.058160503500705264, 32'sd-0.11616641410673084, 32'sd0.06535574993994624, 32'sd-0.09905451759302789, 32'sd0.05266283483442194, 32'sd0.13542096139290488, 32'sd0.0126384155116866, 32'sd-0.09063995209152496, 32'sd-0.3253460818835353, 32'sd0.29070462261628954, 32'sd0.24035786153257652},
        '{32'sd0.07948060045062083, 32'sd0.03549056905413019, 32'sd-0.06499710962291497, 32'sd0.0825227618111894, 32'sd0.14725997727491927, 32'sd-0.020050730651349612, 32'sd0.10243914582830843, 32'sd0.04731014889600568, 32'sd0.02419461298357209, 32'sd-0.10781930938619821, 32'sd0.11012161394342239, 32'sd0.19312337266211727, 32'sd-0.06770986338258471, 32'sd0.165657238942166, 32'sd0.08864162572527436, 32'sd-0.20836034458107142, 32'sd-0.20631747828318073, 32'sd-0.016072415828211378, 32'sd0.06898960917872587, 32'sd-0.18372259975414315, 32'sd-0.0052215606812700335, 32'sd-0.032133753102013336, 32'sd0.18226582824085752, 32'sd-0.06585570446552937, 32'sd0.16518470060662685, 32'sd0.17180160778860157, 32'sd-0.017273412095902406, 32'sd-0.01999998944225605, 32'sd0.02138072019331587, 32'sd0.09426630056819435, 32'sd-0.0810303468926168, 32'sd-0.16538831135264628, 32'sd0.07324203804308342, 32'sd-0.01698970283413757, 32'sd0.0073212776653755664, 32'sd0.006404327121660691, 32'sd-0.009109973291634543, 32'sd0.0686319867290351, 32'sd0.132688457658724, 32'sd0.15775791701733965, 32'sd0.020080622693213222, 32'sd0.1282890163086601, 32'sd0.08521084061881148, 32'sd0.22512907226267542, 32'sd0.29558114057611556, 32'sd-0.1770781926229478, 32'sd-0.13392027177341195, 32'sd0.12711681919863313, 32'sd0.22003765981150733, 32'sd-0.17000426136694757, 32'sd-0.19572089384090843, 32'sd0.29867570276375743, 32'sd-0.16592784856017012, 32'sd-0.2167470083590448, 32'sd0.0354027909147847, 32'sd-0.0020886005812265226, 32'sd-0.0910238888114475, 32'sd0.09671861883688555, 32'sd0.06789907443917936, 32'sd0.11577632578989894, 32'sd-0.22256326372703905, 32'sd-0.2327351306503852, 32'sd-0.1597516192753705, 32'sd0.09062525149200155, 32'sd-0.04429749322594803, 32'sd-0.03279844471461577, 32'sd-0.02564685176119449, 32'sd-0.052647683418192766, 32'sd0.22480300122711877, 32'sd0.026481707258722523, 32'sd-0.1495475627189743, 32'sd0.026616309570949067, 32'sd-0.07555505746939814, 32'sd-0.20733640549262697, 32'sd-0.24191909751135693, 32'sd0.026025095988566553, 32'sd-0.15194970245408299, 32'sd-0.08344922063698053, 32'sd-0.008106479272139817, 32'sd-0.12159712073220255, 32'sd-0.033603847202187447, 32'sd0.035344300796368855, 32'sd-0.06597033967353033, 32'sd0.1839602318490557, 32'sd0.12955927015243882, 32'sd-0.21085355610799328, 32'sd-0.12214908331303492, 32'sd0.16286479425944708, 32'sd-0.225449965041543, 32'sd0.2512278678388468, 32'sd-0.24791980971073677, 32'sd-0.09608932286945657, 32'sd0.02523083069218559, 32'sd0.19650336271941837, 32'sd0.06150124242450493, 32'sd0.10354700441782046, 32'sd0.10796907927823869, 32'sd-0.10630626527285547, 32'sd0.15390051603213126, 32'sd0.24785112968861275, 32'sd0.2038635384499901, 32'sd-0.038882985366916284, 32'sd-0.10647808603960678, 32'sd-0.09523259429193676, 32'sd0.15078285032686067, 32'sd-0.1305727590831742, 32'sd-0.07536990297069078, 32'sd-0.15081873577479765, 32'sd0.15782606800359902, 32'sd-0.006349385502318879, 32'sd-0.12993416877775185, 32'sd-0.2270947211305039, 32'sd0.1982779519209749, 32'sd-0.2646551585389858, 32'sd0.1872889548204997, 32'sd-0.11677573105979476, 32'sd0.216596685441995, 32'sd0.16018174896174892, 32'sd-0.04273281608555754, 32'sd0.20881240345486227, 32'sd0.13579611030557845, 32'sd-0.13294009253835767, 32'sd-0.2589318673253605, 32'sd-0.2631306392605117, 32'sd0.010394119590047383, 32'sd-0.09095157047747285, 32'sd0.28281869066460574, 32'sd0.04935212990081167},
        '{32'sd0.12014938410879922, 32'sd0.04932860962902338, 32'sd-0.15082583963569848, 32'sd-0.0717414255919569, 32'sd0.20493810053550515, 32'sd-0.06672108969079582, 32'sd-0.15322093600236505, 32'sd0.12812641856922607, 32'sd0.11349663453414015, 32'sd-0.15617929451781618, 32'sd0.0012498013533932993, 32'sd0.165933611512451, 32'sd0.08482939232078718, 32'sd0.09185471374194941, 32'sd-0.00273695828679684, 32'sd0.10761580949573422, 32'sd0.10887421495046941, 32'sd-0.07317851992971919, 32'sd-0.23785851248600642, 32'sd0.07184919012237742, 32'sd-0.027409052035325582, 32'sd0.05341926254579673, 32'sd0.24157745784466503, 32'sd0.19244291737899916, 32'sd0.10000484380319692, 32'sd0.08665499936854286, 32'sd-0.25717012314244875, 32'sd0.09058564814770428, 32'sd-0.02980840481186106, 32'sd-0.009057578302275155, 32'sd-0.18024484409736008, 32'sd0.04999320230562195, 32'sd-0.2866905566857385, 32'sd-0.11801639160907795, 32'sd-0.017930894503913285, 32'sd0.17162435584379473, 32'sd-0.15068087708189562, 32'sd-0.13826054656212808, 32'sd-0.059630841592491546, 32'sd0.2296181264745369, 32'sd-0.12115921761289661, 32'sd0.20968145325085233, 32'sd0.14215096139017605, 32'sd0.24484033469704433, 32'sd0.23486933367291962, 32'sd0.12901624437265863, 32'sd-0.19326073907113525, 32'sd0.1362114120067544, 32'sd0.08647347164136462, 32'sd-0.14585642473294272, 32'sd-0.024511530314990735, 32'sd-0.05551522901577837, 32'sd0.09970921178696282, 32'sd0.062077264107735404, 32'sd0.11339664465560137, 32'sd0.0096676330047342, 32'sd-0.1675304811377109, 32'sd0.019294778787817966, 32'sd0.07158669356291526, 32'sd0.08990118681010509, 32'sd-0.21192235401957243, 32'sd-0.10582112466242367, 32'sd0.14003210977437242, 32'sd0.005426283593371047, 32'sd0.22941422348436477, 32'sd0.08576854023545256, 32'sd0.16244092850670738, 32'sd-0.17473193803083054, 32'sd0.12438504786600538, 32'sd-0.19623690471995806, 32'sd0.06840962944079293, 32'sd-0.17895000173064496, 32'sd0.006083249791912483, 32'sd-0.07623006134608526, 32'sd0.0162811083133658, 32'sd0.17251114698986345, 32'sd-0.016860857629140268, 32'sd0.02555787997436995, 32'sd0.18001358365803946, 32'sd-0.07035339389288325, 32'sd-0.1251223092749688, 32'sd-0.13062211414031882, 32'sd0.09286476847872963, 32'sd0.06172015165681298, 32'sd-0.06653626463007882, 32'sd-0.05552076461012273, 32'sd-0.22381917603978677, 32'sd-0.02315564606212353, 32'sd-0.0753493849273143, 32'sd0.06591519976924017, 32'sd-0.19215577000967662, 32'sd-0.18339855220247825, 32'sd-0.002510671899543802, 32'sd0.021893926779355, 32'sd-0.0966558832778744, 32'sd-0.1167557016252092, 32'sd0.10342238780288829, 32'sd-0.15867422890415953, 32'sd-0.05777666495004992, 32'sd0.041495439509152375, 32'sd0.08894434450947343, 32'sd-0.08616467227319477, 32'sd-0.0005838844487558936, 32'sd0.011232295863204733, 32'sd-0.10172436258567548, 32'sd-0.05964545455225842, 32'sd-0.18125394390821306, 32'sd0.07749782664126084, 32'sd-0.1775674077279996, 32'sd0.15170973257677606, 32'sd-0.3204933775228891, 32'sd-0.2275782438331933, 32'sd-0.10220646345977843, 32'sd-0.05982891768282157, 32'sd0.015066991491260335, 32'sd-0.07613760341236936, 32'sd-0.0634409125427506, 32'sd-0.20687743904249517, 32'sd-0.04186699896156766, 32'sd-0.07412620166336395, 32'sd0.07726235901533016, 32'sd0.192684346220247, 32'sd0.1605609730110833, 32'sd-0.1630857436839159, 32'sd0.016717220674309745, 32'sd-0.08207115824311761, 32'sd-0.1794207240732346, 32'sd-0.06724934477612489},
        '{32'sd0.03767418061751362, 32'sd0.13793351869409812, 32'sd-0.1294847068781104, 32'sd0.190046490856709, 32'sd0.09115737817435315, 32'sd-0.1357256860516767, 32'sd0.1686088285892474, 32'sd0.1221459919316296, 32'sd-0.06604141890253667, 32'sd0.07703261711534401, 32'sd-0.00804520362327565, 32'sd-0.06859317589672052, 32'sd0.062056912667864526, 32'sd-0.10595009467980927, 32'sd-0.0423851933702375, 32'sd0.1511943155780066, 32'sd0.12473219389765003, 32'sd0.0702705228066766, 32'sd0.13912813968502338, 32'sd0.0314688795305918, 32'sd0.025926731821058507, 32'sd-0.13334861587293684, 32'sd0.051575566058873826, 32'sd0.015696637518281622, 32'sd0.005873725529142223, 32'sd0.08660593657970073, 32'sd0.2637661887255913, 32'sd-0.023591416364600885, 32'sd0.07235708789216079, 32'sd-0.2512029600669146, 32'sd-0.029577910565110912, 32'sd-0.02881826171876247, 32'sd0.08475152423186352, 32'sd-0.11920933863623034, 32'sd0.1314276434037686, 32'sd0.07661031830174274, 32'sd-0.11000635973377827, 32'sd0.022695418760057963, 32'sd0.09914017159784415, 32'sd-0.12048502334131361, 32'sd0.14496625874635757, 32'sd-0.16018587821646485, 32'sd-0.14307328905255906, 32'sd0.11373433415077447, 32'sd-0.13263128742867078, 32'sd-0.061712079451541925, 32'sd-0.002539286181892642, 32'sd-0.17242989480934082, 32'sd-0.1992414758839117, 32'sd0.09993617798322253, 32'sd-0.012450934552050753, 32'sd0.14468611969969014, 32'sd0.02255343200209056, 32'sd0.17690372471587784, 32'sd-0.18846930536021103, 32'sd-0.009526530665014594, 32'sd0.06984739423238431, 32'sd0.06772154895026412, 32'sd0.11285489332486226, 32'sd0.017750404398156568, 32'sd0.0500874021896763, 32'sd-0.11268334660825627, 32'sd-0.05142635196703549, 32'sd-0.06503295959068474, 32'sd-0.1440185665899517, 32'sd-0.10393639609604083, 32'sd0.03553999207668482, 32'sd0.12958662480342997, 32'sd-0.13851616836917038, 32'sd0.2309820611186802, 32'sd0.0025054365726466196, 32'sd0.12630506955873147, 32'sd0.10927877902073238, 32'sd0.11568316520999297, 32'sd0.12019026330142475, 32'sd0.10634823881204654, 32'sd-0.025851873010458014, 32'sd0.26974934239885673, 32'sd-0.16362382836509912, 32'sd-0.09226980994538893, 32'sd0.002383248022730273, 32'sd0.1933909755708495, 32'sd-0.04064023911183129, 32'sd0.17637118838578247, 32'sd0.03591419466712381, 32'sd-0.14003722850821154, 32'sd0.25104219040476305, 32'sd-0.06340441490340903, 32'sd-0.0831770256150869, 32'sd-0.19909805623637442, 32'sd-0.024527305494520972, 32'sd-0.008618673898929131, 32'sd0.16889721348917147, 32'sd-0.3452318972626937, 32'sd0.22483523422116417, 32'sd-0.13115197974143256, 32'sd0.026773360558324716, 32'sd-0.06221903318103917, 32'sd-0.03646221039033936, 32'sd-0.20520606582199474, 32'sd0.15180157783445938, 32'sd-0.03325095227585232, 32'sd0.2170554511541219, 32'sd-0.044303413331203266, 32'sd-0.11663252755810816, 32'sd0.05942875888366986, 32'sd-0.021579383233362448, 32'sd-0.2976059226097414, 32'sd-0.05993605491827463, 32'sd0.01865230963317486, 32'sd0.151177563111496, 32'sd0.12623666643874668, 32'sd0.10500127573616297, 32'sd-0.07417993600512811, 32'sd0.18884870564781484, 32'sd0.08792879612383743, 32'sd0.030194023668151347, 32'sd-0.004995569856921846, 32'sd0.004280135825709375, 32'sd-0.006876587237063991, 32'sd0.12557903302542497, 32'sd0.22910482536421004, 32'sd-0.06511895170175656, 32'sd0.07762772143490139, 32'sd-0.16559908613110505, 32'sd0.20629982095536006, 32'sd-0.12078631541178789, 32'sd0.027160327650558126},
        '{32'sd-0.061487752161402176, 32'sd0.20629667847658023, 32'sd0.11878149468770006, 32'sd-0.01651299027568884, 32'sd0.054701350178707434, 32'sd-0.15262095866177108, 32'sd-0.16497727186293623, 32'sd-0.0365605987048468, 32'sd0.08742833733142033, 32'sd-0.05897831642669954, 32'sd-0.1191352324744369, 32'sd-0.12208174150945053, 32'sd-0.1243454536347622, 32'sd0.009997624491697218, 32'sd0.2039890693162466, 32'sd-0.03993291074907355, 32'sd-0.17524548695423764, 32'sd0.1262841627147397, 32'sd0.27071584135926163, 32'sd0.10273754615753228, 32'sd-0.019868434992507115, 32'sd-0.238356650694711, 32'sd0.015441891805168724, 32'sd0.08737629474903018, 32'sd-0.18457554853272828, 32'sd-0.13037129236117007, 32'sd0.019712122839342275, 32'sd0.062417815641715196, 32'sd-0.08421340828430493, 32'sd-0.20471959148756236, 32'sd-0.00022951940617967572, 32'sd-0.041289393324056185, 32'sd0.1634873252434407, 32'sd-0.0673696080976015, 32'sd-0.02090523314411254, 32'sd0.011555828294713008, 32'sd0.10048412243020381, 32'sd-0.0727320215290728, 32'sd0.10708453143945564, 32'sd0.0724986281120085, 32'sd-0.29329576875400665, 32'sd-0.025536751888671202, 32'sd0.19012456028345637, 32'sd0.08452838426907186, 32'sd0.16053494599335344, 32'sd0.09727948118621957, 32'sd-0.08352822660453961, 32'sd-0.11156937071939717, 32'sd0.17070992787023942, 32'sd0.18017930949152228, 32'sd-0.14951387573090613, 32'sd0.004804944353738089, 32'sd-0.12076786899087312, 32'sd-0.015132887539525852, 32'sd-0.004577962138970363, 32'sd-0.18301642193307643, 32'sd-0.11232364574752078, 32'sd-0.2614524640243119, 32'sd0.13579274869109376, 32'sd0.12936252021894143, 32'sd0.1979592721601317, 32'sd0.26501472081863275, 32'sd0.13513669041721127, 32'sd0.1412877614721289, 32'sd0.01829487768899927, 32'sd0.11849444541239232, 32'sd-0.06822883700265316, 32'sd0.006409626637432239, 32'sd0.13144863213909275, 32'sd-0.006288611480758653, 32'sd0.04532787478409133, 32'sd0.14168412785845969, 32'sd-0.16391718475502579, 32'sd-0.09333878041619965, 32'sd0.03497582394378468, 32'sd0.1988631909392496, 32'sd0.06291880961053353, 32'sd-0.016505389053154858, 32'sd0.1595932144473026, 32'sd-0.17257630747133504, 32'sd-0.17742540209968402, 32'sd-0.06751452827351759, 32'sd0.027768176199404953, 32'sd-0.07352735293360807, 32'sd0.157320756474332, 32'sd0.060454250930343734, 32'sd0.1518081078130619, 32'sd-0.17376292688730244, 32'sd0.024963382673338433, 32'sd0.1859327846004493, 32'sd0.07102992077162616, 32'sd-0.04617794535243129, 32'sd0.15316027859597334, 32'sd0.061001735131458984, 32'sd-0.1916364992007709, 32'sd0.1434288492850735, 32'sd-0.17864169227344412, 32'sd-0.16597250677228975, 32'sd-0.10249069655031115, 32'sd0.035658397774956024, 32'sd0.12415504461302408, 32'sd-0.002112206568292452, 32'sd0.038387939555432224, 32'sd0.029406050425182684, 32'sd0.1579828908745032, 32'sd0.03462241475700448, 32'sd-0.05300292667123728, 32'sd0.16631210469417643, 32'sd0.0928906537837347, 32'sd-0.13412650970310575, 32'sd0.14236413174098994, 32'sd0.08726033152649171, 32'sd-0.2302269347548079, 32'sd0.048184499248079625, 32'sd0.08619998540501903, 32'sd0.04289807326469431, 32'sd-0.13715145714611576, 32'sd0.29551545587107375, 32'sd-0.18162362307815555, 32'sd0.1882195099175742, 32'sd-0.11641360756413809, 32'sd-0.03587121125637819, 32'sd0.15825001011379736, 32'sd0.13570663537906852, 32'sd0.051675599482621674, 32'sd-0.18795700830046128, 32'sd0.12468207147057157, 32'sd0.10830033797014728},
        '{32'sd-0.03785864685877041, 32'sd-0.017611517864506532, 32'sd-0.10309387341881088, 32'sd0.09085820528148714, 32'sd-0.19862726870357064, 32'sd0.008986385539074453, 32'sd0.08441842926552837, 32'sd0.020579492611168503, 32'sd-0.07461761739731163, 32'sd0.20318047875198128, 32'sd0.07252506215647654, 32'sd0.12218968094368561, 32'sd0.13733437691810887, 32'sd-0.09987567172611747, 32'sd-0.02246637626466572, 32'sd0.0584763578069982, 32'sd0.145034260462878, 32'sd0.18737879132224647, 32'sd0.09120118846646455, 32'sd-0.07937001914638545, 32'sd-0.31708663301251433, 32'sd0.006092934428170983, 32'sd-0.1268113762695405, 32'sd0.09794979467601585, 32'sd0.07421418020422872, 32'sd0.01577737291632841, 32'sd0.01288988238316038, 32'sd-0.061761807589370804, 32'sd-0.133429800028395, 32'sd0.09755826215239782, 32'sd0.176140764374631, 32'sd0.18797980525942815, 32'sd-0.030910637254192585, 32'sd0.16294229634282065, 32'sd0.10292963958465627, 32'sd0.13859800815619222, 32'sd-0.13994452573525779, 32'sd-0.28049971505139626, 32'sd0.174387576404345, 32'sd-0.06332128643916934, 32'sd0.07266722054546722, 32'sd-0.24005070817956592, 32'sd0.016260421522699763, 32'sd-0.05530145298210593, 32'sd0.1567238139905398, 32'sd-0.23419313761486588, 32'sd-0.018406067531294826, 32'sd0.05576618980325146, 32'sd-0.26637717945550576, 32'sd0.011254554968846458, 32'sd0.06765462458879629, 32'sd-0.04702776712814812, 32'sd0.1843459428915762, 32'sd-0.1686186713442151, 32'sd-0.2147789543713049, 32'sd-0.03507702909678854, 32'sd-0.21980231966538977, 32'sd-0.0026901608488094147, 32'sd0.08172987682240297, 32'sd0.28529945119608807, 32'sd0.09728993183708294, 32'sd0.1427860011291047, 32'sd0.07057737738589664, 32'sd-0.25659331982160055, 32'sd-0.2998235610056939, 32'sd-0.18076255198390828, 32'sd0.10157507598643871, 32'sd0.043022961530404566, 32'sd-0.03533167866996781, 32'sd-0.15081885187848323, 32'sd0.11713122683677865, 32'sd-0.24201271600988639, 32'sd-0.09740618581189567, 32'sd-0.17435574995607725, 32'sd0.08451525569722498, 32'sd-0.19337876252131295, 32'sd-0.03105166568909, 32'sd-0.08078918964773553, 32'sd-0.30607073647333694, 32'sd0.021492365978621853, 32'sd-0.15930202471104576, 32'sd0.09624255609214563, 32'sd0.3005835210246125, 32'sd-0.07623683087803769, 32'sd0.09661895298209901, 32'sd0.0698367743035846, 32'sd0.1791757503848116, 32'sd-0.11890729585049781, 32'sd0.11844908770084206, 32'sd-0.17034918378264632, 32'sd0.08029682868905123, 32'sd-0.08847265924045257, 32'sd0.08218973625012099, 32'sd-0.16547733355140218, 32'sd-0.16854800802063244, 32'sd-0.09119039369942847, 32'sd0.19013155420016403, 32'sd0.1937949095346858, 32'sd-0.19153408806116337, 32'sd-0.09793194288653478, 32'sd-0.023122075141871014, 32'sd-0.17896709570924832, 32'sd0.04731889423275159, 32'sd0.04162733693484299, 32'sd0.11024005355666826, 32'sd0.2098255666185538, 32'sd0.2790309483285033, 32'sd0.03280272909013115, 32'sd-0.20505338890548003, 32'sd0.11255738589537026, 32'sd0.11948189849303678, 32'sd0.05070265078603257, 32'sd0.19888281153067042, 32'sd0.0228836497113379, 32'sd-0.02487565355164403, 32'sd0.125102768654253, 32'sd-0.09640150740822875, 32'sd0.13265469682992087, 32'sd-0.11420634944604317, 32'sd0.06689004571128446, 32'sd-0.02903044463536759, 32'sd0.08011949080274106, 32'sd-0.01092810266139501, 32'sd0.1267570474356569, 32'sd0.037485500137908016, 32'sd-0.08329414639100871, 32'sd-0.1486918797952588, 32'sd-0.04496950706941584},
        '{32'sd0.04229688878948161, 32'sd-0.10289145124912642, 32'sd-0.12311946524411334, 32'sd0.07189580790167083, 32'sd-0.16166664909633374, 32'sd-0.06223322509979736, 32'sd-0.12557900952180118, 32'sd0.18493193105485484, 32'sd0.052748643524560254, 32'sd0.13652980711763604, 32'sd0.03247614520365451, 32'sd-0.09140055403175215, 32'sd0.24257278509880975, 32'sd0.15075598216021954, 32'sd-0.09749649014371531, 32'sd0.076797748599309, 32'sd-0.2076119378016595, 32'sd-0.12016770835265213, 32'sd-0.26643622234230663, 32'sd0.0448094498836833, 32'sd-0.12753440123443593, 32'sd0.12039362563240928, 32'sd-0.15112778935129642, 32'sd-0.020332571871647435, 32'sd-0.1812954278359428, 32'sd-0.060698223737654905, 32'sd0.07412519893280299, 32'sd0.15042082847641136, 32'sd-0.2103591620156475, 32'sd-0.12862914938807962, 32'sd-0.11939241171231427, 32'sd-0.16649256804526488, 32'sd0.15000073082182938, 32'sd-0.020619969638060846, 32'sd0.1396239568465699, 32'sd-0.22739220097306276, 32'sd0.006789966812198402, 32'sd-0.02695507359065622, 32'sd0.060381123467955454, 32'sd-0.11954162159357043, 32'sd0.16683384903765217, 32'sd-0.09157664168735112, 32'sd0.1971103485940297, 32'sd0.15669275281969813, 32'sd-0.03778145185384493, 32'sd0.0908608154676893, 32'sd0.1202021546648212, 32'sd0.01318531903270879, 32'sd0.020506142315263324, 32'sd-0.0845326970854913, 32'sd0.2127220568859425, 32'sd0.056292182081839864, 32'sd-0.06816735517765567, 32'sd-0.09221747167585079, 32'sd0.05199057494004364, 32'sd0.01773949730956253, 32'sd0.10093212385133897, 32'sd0.13472448836037323, 32'sd-0.08701523206343695, 32'sd0.129847816770839, 32'sd-0.08489309990878344, 32'sd0.10855803012441193, 32'sd-0.09023319857625582, 32'sd0.09044104586112375, 32'sd-0.008178119980811109, 32'sd0.0036293050551400594, 32'sd0.11551139991204196, 32'sd-0.03255284227798406, 32'sd-0.008617544395907988, 32'sd-0.1694301037086018, 32'sd-0.03545912619776243, 32'sd0.004048228714442293, 32'sd-0.003935659358432236, 32'sd0.0517762554073604, 32'sd-0.14312206424266125, 32'sd-0.18085832671884322, 32'sd-0.06692367976472044, 32'sd0.2523492228854565, 32'sd-0.05602962471583271, 32'sd0.21609741523350964, 32'sd-0.015599618411378068, 32'sd-0.25314086701926447, 32'sd-0.15530899132699874, 32'sd0.0009259737318651582, 32'sd0.15012769536677834, 32'sd-0.14523857400679652, 32'sd-0.22724113220423378, 32'sd0.007816835913344802, 32'sd-0.10475689142338028, 32'sd0.09163900969067466, 32'sd0.16276398846993456, 32'sd0.021874752230202264, 32'sd-0.044749987330539254, 32'sd0.04332313306629593, 32'sd-0.05745242549329063, 32'sd0.20497304784572098, 32'sd-0.1483223667423531, 32'sd0.05861149959690669, 32'sd0.1732886747416771, 32'sd-0.0524960883795452, 32'sd0.18023768278003713, 32'sd-0.027189450692148624, 32'sd-0.10705187969437863, 32'sd0.006272436962310423, 32'sd0.1418627679568822, 32'sd-0.22245499480414727, 32'sd-0.04455515037827374, 32'sd-0.05471923143564089, 32'sd0.19257225495138164, 32'sd0.13816837001364124, 32'sd0.046738259927839226, 32'sd0.19402595962716468, 32'sd0.13876697431826118, 32'sd-0.04906475977004714, 32'sd0.15251565894487448, 32'sd0.037345358515821374, 32'sd-0.08821758854830797, 32'sd0.16955231257763417, 32'sd-0.1277085069443808, 32'sd-0.13884372754420413, 32'sd0.20671041603589627, 32'sd0.05121322472645607, 32'sd-0.06381628414438184, 32'sd-0.07830875878017307, 32'sd0.23456897965124213, 32'sd0.14706625466169732, 32'sd0.24449248989617886, 32'sd-0.0817626819691335},
        '{32'sd0.20477042729452297, 32'sd-0.2143241816061529, 32'sd-0.12278054378798166, 32'sd-0.021241598350680863, 32'sd0.06596645307419016, 32'sd-0.023462822774853613, 32'sd0.05218360781927266, 32'sd0.009593490516741281, 32'sd-0.24497645054723888, 32'sd-0.031895884981886904, 32'sd0.06544907015793065, 32'sd-0.19609726837329433, 32'sd0.15325460923366027, 32'sd-0.13969573810408356, 32'sd-0.07764179292941571, 32'sd0.11664054873253538, 32'sd-0.03671902714858169, 32'sd-0.1541038654528207, 32'sd-0.23227777836080168, 32'sd0.024493187117079523, 32'sd0.10516152969355638, 32'sd0.09845818364070232, 32'sd-0.05557337788860788, 32'sd0.10670660078783019, 32'sd-0.11161770368091109, 32'sd0.1234397844383107, 32'sd0.12669231862988775, 32'sd-0.12335082912568439, 32'sd-0.13153493522704607, 32'sd-0.2151611801320954, 32'sd-0.16747815365144048, 32'sd-0.159228344565437, 32'sd0.11279569265474496, 32'sd0.16246433422984072, 32'sd-0.1188970698649798, 32'sd0.15770144540978925, 32'sd0.22807089552285478, 32'sd0.1890529596446082, 32'sd-0.11967545971324473, 32'sd-0.0019290262354016575, 32'sd0.20612836072790003, 32'sd0.07704874767715703, 32'sd0.08512105369018826, 32'sd-0.293750756978361, 32'sd-0.10425533952647117, 32'sd0.2237477933233786, 32'sd-0.04360252137887331, 32'sd0.17347876160657383, 32'sd0.09264822696107038, 32'sd0.03982562242990089, 32'sd0.11398665773082461, 32'sd-0.04624763200065574, 32'sd0.08044213118156966, 32'sd0.09284392776477833, 32'sd-0.033169220561846784, 32'sd0.0352050794799816, 32'sd-0.030873563338263046, 32'sd-0.18199462651591394, 32'sd-0.03984825826888406, 32'sd0.107577105135214, 32'sd-0.12806128292130053, 32'sd0.1700467503956382, 32'sd0.11407901693090826, 32'sd0.1533789989155347, 32'sd-0.155758039723773, 32'sd0.05168993452441588, 32'sd-0.08339068429126263, 32'sd0.061030593356206815, 32'sd-0.021537024716444968, 32'sd-0.06806253732836455, 32'sd0.1687320899330858, 32'sd0.06803875820599148, 32'sd0.16965647542346562, 32'sd-0.0881040549221905, 32'sd0.07951225742318957, 32'sd0.02773384213791223, 32'sd-0.13479429252461447, 32'sd-0.03809005243071693, 32'sd-0.06766249875253702, 32'sd-0.13486368664762463, 32'sd0.04889472745319166, 32'sd-0.1395350155396432, 32'sd-0.01046883022183714, 32'sd0.1423168476277267, 32'sd0.10639317372520259, 32'sd-0.022047504096078904, 32'sd-0.23828434201089027, 32'sd0.1409468798895029, 32'sd0.18303957860198433, 32'sd-0.21969649972374883, 32'sd0.17783580518073785, 32'sd0.22700796519613317, 32'sd-0.13850676395803851, 32'sd-0.13173857570516437, 32'sd-0.13008499107557783, 32'sd-0.052956710710560774, 32'sd0.026953277106140452, 32'sd0.05182267650960927, 32'sd-0.05180339626299026, 32'sd0.05525006931042079, 32'sd-0.04861742465534763, 32'sd0.1347809413971752, 32'sd0.0267038987619384, 32'sd0.1478936688584105, 32'sd-0.03937570185271132, 32'sd-0.08633662339463755, 32'sd0.10219367869316655, 32'sd-0.10354995727798694, 32'sd0.16232958508527523, 32'sd-0.03068677459366145, 32'sd0.19594817861995892, 32'sd0.19130894775254811, 32'sd-0.2446784270518513, 32'sd0.15903971412568363, 32'sd0.09941218370441753, 32'sd-0.11209618562653482, 32'sd0.050231451608683426, 32'sd0.09451561139271221, 32'sd0.04496142317785813, 32'sd0.12948997816233507, 32'sd0.14200102127891992, 32'sd0.09195744934096037, 32'sd-0.11778415135457919, 32'sd0.24136696851233005, 32'sd0.2312841868970587, 32'sd0.17102552440496874, 32'sd0.04499876267881313, 32'sd-0.018079643671169276},
        '{32'sd0.2210269911149397, 32'sd0.1093833613648068, 32'sd-0.09432618532815762, 32'sd-0.19212072995506946, 32'sd-0.11960800507912231, 32'sd0.10932106763605445, 32'sd0.006963988180058412, 32'sd0.02049446346998514, 32'sd-0.09000451797571225, 32'sd0.050553309338016, 32'sd0.01901863325721113, 32'sd0.14547145735841557, 32'sd0.005381927606630004, 32'sd-0.05926182548533494, 32'sd-0.0487563794652234, 32'sd-0.20121726890722255, 32'sd0.13906810879326711, 32'sd-0.010112709394106231, 32'sd0.07130964655293279, 32'sd0.17347203728607904, 32'sd0.2358837389030382, 32'sd-0.06040643146532121, 32'sd0.14434783229249834, 32'sd-0.15287782281355375, 32'sd-0.19982301581227913, 32'sd-0.09283174111688884, 32'sd0.1798838880315068, 32'sd0.20496247439148546, 32'sd0.026631750114829687, 32'sd-0.0343042193581078, 32'sd0.14898732135505102, 32'sd-0.05790563621001795, 32'sd0.10264751183979767, 32'sd-0.1856853453447989, 32'sd-0.215510488121492, 32'sd-0.018266808135832948, 32'sd-0.049950306758813554, 32'sd0.01699446876183349, 32'sd0.14153600989453433, 32'sd-0.07353798085346942, 32'sd0.02917993546248014, 32'sd0.07505318046122578, 32'sd0.15801381005186982, 32'sd-0.245452442314309, 32'sd0.07535805498576724, 32'sd-0.016980864756378295, 32'sd-0.09988700541133085, 32'sd0.13509661097923753, 32'sd0.11906520558617374, 32'sd0.07268253494065666, 32'sd-0.2199468921279914, 32'sd-0.09873302484866993, 32'sd-0.05527334897955501, 32'sd0.0683261126604434, 32'sd-0.09343121867635834, 32'sd-0.1818272154348172, 32'sd-0.0984781507192796, 32'sd-0.13134984548779238, 32'sd-0.07793586404117694, 32'sd0.20615562673501833, 32'sd-0.02689844784551789, 32'sd-0.09814953855143294, 32'sd0.12081914035741449, 32'sd0.13697547849959057, 32'sd0.21415934117454732, 32'sd-0.2433862737676833, 32'sd-0.06490221029467551, 32'sd-0.07681701048514165, 32'sd0.1800866146790647, 32'sd0.12022086703305833, 32'sd-0.13858653650403258, 32'sd0.07268681847733392, 32'sd-0.4520659150867844, 32'sd0.08637509038996244, 32'sd-0.1926033787934993, 32'sd-0.23485697321544027, 32'sd-0.14729255028718086, 32'sd0.033233247872615855, 32'sd-0.20587553919030913, 32'sd-0.1851024554396939, 32'sd-0.1030109995884965, 32'sd0.18175498969440124, 32'sd-0.11568791844881071, 32'sd-0.16700002685794924, 32'sd-0.09153683516725776, 32'sd-0.034905536826197577, 32'sd0.24459992225247765, 32'sd0.044351207108204324, 32'sd-0.022213683455456816, 32'sd-0.08852394439621446, 32'sd0.09101322792478611, 32'sd-0.168223991326496, 32'sd-0.2177141378038605, 32'sd0.07434108753977253, 32'sd0.02504756642423279, 32'sd-0.0742715234493012, 32'sd-0.22428655841944747, 32'sd0.21756368674840135, 32'sd0.16686742456050718, 32'sd0.1319794526830404, 32'sd0.14348551724682845, 32'sd-0.0924866958126697, 32'sd-0.10183874756908855, 32'sd0.09510859154663594, 32'sd0.18346122923962846, 32'sd-0.05722054661831769, 32'sd0.03986565924233801, 32'sd0.08053776368961574, 32'sd0.17822871094928955, 32'sd-0.02225558619418041, 32'sd-0.1445309845760371, 32'sd0.2692472558584905, 32'sd0.023325025292718488, 32'sd-0.06764135881256741, 32'sd-0.20150678774397715, 32'sd0.015943397584005814, 32'sd0.12115524765168925, 32'sd-0.14171754388723562, 32'sd0.28522225570179505, 32'sd0.12183733639318262, 32'sd0.21968955741798535, 32'sd0.1458641588134154, 32'sd0.006013425008356948, 32'sd-0.20617049999453801, 32'sd-0.3133599220595369, 32'sd0.0003895306731147529, 32'sd0.21327399456278046, 32'sd-0.10795196318942357},
        '{32'sd0.07580577364909441, 32'sd0.05427182155008132, 32'sd-0.0816321894819817, 32'sd-0.04336411710553221, 32'sd0.1803777457637192, 32'sd0.17629707409655745, 32'sd-0.005964758141487546, 32'sd-0.08731155735141541, 32'sd-0.14226944887431622, 32'sd-0.15245494014899724, 32'sd-0.054220104163398376, 32'sd0.16802384303270998, 32'sd-0.22773400531340282, 32'sd0.10704855340608845, 32'sd0.11976774550582077, 32'sd0.01653819116856033, 32'sd-0.055356691237418716, 32'sd-0.11105241563147521, 32'sd0.05598198431594394, 32'sd0.2010429853379043, 32'sd0.03533618839586426, 32'sd-0.06314068567337151, 32'sd0.12410161626360845, 32'sd0.02289716336708766, 32'sd0.15471348228867685, 32'sd-0.03065848211034378, 32'sd-0.20655933919349975, 32'sd-0.1564503527951901, 32'sd0.2468031905507024, 32'sd-0.08361138769812737, 32'sd0.14321918574229175, 32'sd-0.08703378270296895, 32'sd-0.26146788311754504, 32'sd-0.014835193828004757, 32'sd0.18588485460797097, 32'sd-0.05325353528123396, 32'sd-0.022902317673248525, 32'sd-0.003210350753264396, 32'sd-0.12496234775278359, 32'sd0.19085094468329594, 32'sd-0.09527850031509588, 32'sd-0.04792101965821149, 32'sd0.17870859701360922, 32'sd-0.015351904382235007, 32'sd-0.17453467160384933, 32'sd0.1356640392048944, 32'sd-0.21219039479121868, 32'sd0.26737758561111974, 32'sd-0.21374710136083475, 32'sd-0.0681049188484165, 32'sd-0.034407602888075116, 32'sd0.005067554986294894, 32'sd0.17634647736171077, 32'sd-0.04081771939131186, 32'sd0.14045139486709207, 32'sd-0.15679593337801323, 32'sd0.08588852269884935, 32'sd-0.10785231313298446, 32'sd0.12620378996644596, 32'sd0.06137345636886117, 32'sd0.12216960770634017, 32'sd-0.010602307838075496, 32'sd-0.18381027140948122, 32'sd-0.16867441529399035, 32'sd0.07382307384397707, 32'sd0.1963778674901868, 32'sd0.10560823880539925, 32'sd-0.051705222852971015, 32'sd0.13735214210178487, 32'sd0.10488540850837151, 32'sd0.014959639378675543, 32'sd-0.12937315176033434, 32'sd-0.0752494982018406, 32'sd-0.11841661178075513, 32'sd0.16309806230652396, 32'sd0.20551499676624468, 32'sd0.17480404202104896, 32'sd-0.039484802051380066, 32'sd-0.0018232836821584773, 32'sd-0.2034704709738547, 32'sd0.0013903531874489919, 32'sd0.03945793304921321, 32'sd-0.0027957807634187374, 32'sd-0.11944068918966941, 32'sd0.16736662690336127, 32'sd0.14072086343110177, 32'sd0.1726954464649812, 32'sd0.025669362205343063, 32'sd-0.03784821618480507, 32'sd-0.06237039145366265, 32'sd-0.2051967177613115, 32'sd-0.17175485128235093, 32'sd-0.10232754073562783, 32'sd0.0976157643395648, 32'sd0.12240143893315386, 32'sd0.0068971173132159076, 32'sd0.0648624206372317, 32'sd0.12599792074785435, 32'sd-0.08562410187507025, 32'sd-0.02027433225781481, 32'sd0.16006953485457392, 32'sd0.0570940184129271, 32'sd-0.08630182782972307, 32'sd0.053384068783280315, 32'sd0.08950697855665557, 32'sd-0.17119614765188962, 32'sd-0.085773987660819, 32'sd0.044645470287949546, 32'sd0.10540290238991004, 32'sd0.1782645810688376, 32'sd0.02354315304890684, 32'sd-0.239667908470478, 32'sd-0.0059576917806464765, 32'sd0.08373681853913029, 32'sd0.1957461617071722, 32'sd0.09857314248680643, 32'sd-0.005419460540950046, 32'sd0.3002591920509713, 32'sd0.19777668215259775, 32'sd-0.05147633962964592, 32'sd-0.04993643660371822, 32'sd0.15911623696448096, 32'sd-0.15355384921953566, 32'sd-0.024133564969347154, 32'sd-0.09661317979460682, 32'sd-0.046697970658987495, 32'sd-0.0682949991562442, 32'sd0.1704079791248041},
        '{32'sd0.11722801849163494, 32'sd-0.16375767795720206, 32'sd0.09968562586790526, 32'sd-0.1345534142963603, 32'sd0.21659048454264476, 32'sd-0.2779893934996315, 32'sd-0.16192394526835924, 32'sd-0.05873879225694935, 32'sd-0.120267452317842, 32'sd-0.22188753221863075, 32'sd-0.08266983625705841, 32'sd0.10676841125478088, 32'sd-0.11516553483851381, 32'sd-0.02824851922307541, 32'sd-0.06634282483357473, 32'sd-0.04233737599287937, 32'sd-0.07021739096587198, 32'sd0.14836125722417154, 32'sd-0.05019332600797847, 32'sd-0.011889515445226843, 32'sd0.00632494402883105, 32'sd0.12832508715601681, 32'sd0.0970177539447595, 32'sd-0.021247716908247866, 32'sd0.02675094420901577, 32'sd-0.14410397743538217, 32'sd-0.16101270588893182, 32'sd-0.10517897503003096, 32'sd-0.014115645666806152, 32'sd0.028698246007017682, 32'sd0.1165885748202589, 32'sd0.2391899000189136, 32'sd-0.05444615091626422, 32'sd0.07199780967797312, 32'sd-0.04001406700625005, 32'sd0.047749663883072835, 32'sd-0.24356103334463994, 32'sd-0.12064869144160746, 32'sd-0.16904506213958634, 32'sd0.18185969946038508, 32'sd0.1504729333760725, 32'sd0.06067048194627167, 32'sd-0.09118140765073894, 32'sd-0.034522840497066005, 32'sd-0.2148408649839936, 32'sd0.13440030386917726, 32'sd-0.09676747101322981, 32'sd-0.03541548971493434, 32'sd0.24460735557911842, 32'sd0.1349190709389482, 32'sd-0.1344973170896673, 32'sd-0.14304673551608313, 32'sd-0.09740008304999814, 32'sd0.08397593649724841, 32'sd-0.04335295416721404, 32'sd-0.24477004054974363, 32'sd-0.1255641696757753, 32'sd-0.24139882806665405, 32'sd0.17992085069599217, 32'sd-0.10344595515831777, 32'sd-0.2357063541843794, 32'sd0.013402878825834099, 32'sd-0.06752518035842162, 32'sd-0.05014024307313153, 32'sd-0.059460389008901625, 32'sd0.0686792217286218, 32'sd0.1142586395569708, 32'sd-0.06220657885017272, 32'sd0.09527359165491203, 32'sd-0.015390458918289026, 32'sd0.10053380948992698, 32'sd0.05018429751835063, 32'sd-0.03378478272952041, 32'sd-0.11346722979122545, 32'sd-0.01078371089619042, 32'sd0.0922906987117759, 32'sd0.1328748077033083, 32'sd0.02261826325748204, 32'sd0.14307194124571154, 32'sd0.15117617696420618, 32'sd0.15857862040347837, 32'sd-0.06278875353695688, 32'sd0.10033238527663486, 32'sd0.04914895368217769, 32'sd-0.17622189899248905, 32'sd0.16161669064118345, 32'sd-0.17420907087761228, 32'sd-0.21360523909191803, 32'sd-0.1206682715471106, 32'sd0.0903165859592079, 32'sd-0.0930033877922161, 32'sd-0.16711663452558634, 32'sd-0.08952863078117247, 32'sd-0.12039114082256153, 32'sd-0.07742321406846735, 32'sd-0.17747226749354403, 32'sd-0.03321347056496153, 32'sd0.12215078970575954, 32'sd0.01006409293793662, 32'sd0.023721146368173403, 32'sd-0.03788622214986656, 32'sd-0.1421248515133502, 32'sd0.13819320326111992, 32'sd-0.06397027056638367, 32'sd0.049895255957289185, 32'sd0.14734696294728483, 32'sd0.0006138849998503816, 32'sd0.07144166378565238, 32'sd-0.11260109644927488, 32'sd-0.1119231239627378, 32'sd-0.0015926573336751233, 32'sd-0.06883465419153609, 32'sd0.2951764409395066, 32'sd-0.045972683664529154, 32'sd0.023068354146884615, 32'sd-0.13620574102517682, 32'sd-0.07645966227429522, 32'sd-0.061345668166528464, 32'sd0.10050076424238329, 32'sd-0.32994217354806327, 32'sd-0.13466929683890513, 32'sd0.0821875449408527, 32'sd-0.19117102974495953, 32'sd-0.2506539534220104, 32'sd-0.10276860626649922, 32'sd-0.0918450889523844, 32'sd0.09019819292649005, 32'sd0.13851934418193074},
        '{32'sd0.07134620535772977, 32'sd0.20619349774689835, 32'sd0.003976890844238708, 32'sd-0.11279173318778392, 32'sd-0.016384998812577777, 32'sd-0.22415090782912708, 32'sd0.1562633917550526, 32'sd0.13978671046480465, 32'sd-0.12791262246912524, 32'sd-0.22583112120685997, 32'sd-0.10120826775813943, 32'sd0.09381693075405387, 32'sd0.07308246808762485, 32'sd0.1884970558433879, 32'sd0.1288647111117054, 32'sd0.018681877956590626, 32'sd-0.01916690685842788, 32'sd0.021917632399109675, 32'sd-0.19638607210440023, 32'sd0.06392570573663466, 32'sd0.04209964542910054, 32'sd0.10756852699923165, 32'sd0.023213663665229443, 32'sd0.12035875751779394, 32'sd-0.18714802061001165, 32'sd-0.15858704114104485, 32'sd0.11840217048309495, 32'sd-0.055811962470280356, 32'sd-0.3812463141357382, 32'sd-0.08584654568397627, 32'sd0.05809734299916545, 32'sd-0.10959078863162346, 32'sd0.03799297951599059, 32'sd-0.0962280902416583, 32'sd-0.13870550346992555, 32'sd-0.17926049345537998, 32'sd0.23550726402574382, 32'sd-0.18194378917410384, 32'sd0.11301299075594368, 32'sd0.11844187633134055, 32'sd0.0018940591992815407, 32'sd0.08325701522193404, 32'sd-0.14047309615621753, 32'sd0.07957034494138088, 32'sd-0.03477079067434378, 32'sd0.18774582598895964, 32'sd0.055173444115686025, 32'sd0.06116541796995841, 32'sd-0.08138743372706336, 32'sd-0.14392229590254427, 32'sd0.270071159792913, 32'sd-0.05022479361492982, 32'sd-0.13809601158256696, 32'sd-0.19181877107826725, 32'sd0.001608424358553625, 32'sd0.04469675575679817, 32'sd-0.12442827119366345, 32'sd-0.01738457695174485, 32'sd-0.08300685012193176, 32'sd-0.11915491893065838, 32'sd0.08056556089331601, 32'sd-0.02710451679253849, 32'sd0.0028677168391980945, 32'sd-0.02722985227592142, 32'sd0.10438391152551663, 32'sd-0.1443448518568865, 32'sd-0.11197959196331672, 32'sd-0.24294222315397565, 32'sd0.15492323686213144, 32'sd0.0019138546326288382, 32'sd0.1126670220357947, 32'sd0.14966161622849994, 32'sd0.15387032635587045, 32'sd0.15723303778000516, 32'sd-0.014835915800943206, 32'sd-0.18259156444852237, 32'sd0.1591062308737139, 32'sd0.06835717614328493, 32'sd0.0216586156048679, 32'sd-0.14536427979221742, 32'sd-0.05495530868222657, 32'sd0.11122849319250559, 32'sd0.13602081000913072, 32'sd0.08126178153165012, 32'sd0.16771837024790612, 32'sd-0.012545623793774264, 32'sd-0.04399513079937559, 32'sd-0.02205373383243324, 32'sd0.19314155972980285, 32'sd-0.12226440223492749, 32'sd0.12872756376793631, 32'sd0.16232687541319502, 32'sd-0.20967304658135952, 32'sd0.11394795728227715, 32'sd0.007875158097116168, 32'sd0.04961108435228645, 32'sd-0.15517011423092822, 32'sd0.0811874278328062, 32'sd-0.22364176748243964, 32'sd0.172978618818451, 32'sd-0.1287133991722643, 32'sd0.024420375137332393, 32'sd-0.11613962901898957, 32'sd0.09478535737382952, 32'sd-0.16002622341324954, 32'sd0.15744505194241196, 32'sd0.23990441765554113, 32'sd0.16805568773349538, 32'sd0.09363922056074253, 32'sd0.03480396743904506, 32'sd0.0700908472335954, 32'sd0.08108883392618854, 32'sd0.15575231757835292, 32'sd-0.08594160098171724, 32'sd0.0027634846054287146, 32'sd0.06713181356055734, 32'sd0.0767667872111465, 32'sd-0.24432820587516413, 32'sd0.06587909950885662, 32'sd0.247984720378706, 32'sd0.14308993984035787, 32'sd0.07978171227548825, 32'sd-0.257810872787439, 32'sd-0.021353647419773455, 32'sd0.047667542092554735, 32'sd-0.011622253872532197, 32'sd0.12440078115561107, 32'sd0.04479821225775515},
        '{32'sd-0.14358927313987455, 32'sd0.15004718286215402, 32'sd-0.1083073573040616, 32'sd0.0775949737555797, 32'sd-0.19916676288487328, 32'sd-0.18530660668852503, 32'sd-0.16286924524298696, 32'sd-0.21677843393406504, 32'sd0.06748502305135642, 32'sd0.2393183543475962, 32'sd0.08072663609239122, 32'sd0.19010328587427855, 32'sd0.13795248996962114, 32'sd0.0021016272769636157, 32'sd0.044756523446303605, 32'sd0.13518074445954587, 32'sd-0.20525630299189687, 32'sd-0.1999457248431527, 32'sd-0.015920132839292125, 32'sd-0.17404948687019856, 32'sd0.19263216474907216, 32'sd-0.141157372540458, 32'sd0.017976892698272386, 32'sd0.15423386403369618, 32'sd-0.09796733612175655, 32'sd-0.15263495957279766, 32'sd0.09537228974647284, 32'sd-0.09346679235065863, 32'sd0.23169156555996706, 32'sd0.14679951029213134, 32'sd-0.03762646744070617, 32'sd0.03291021052755558, 32'sd-0.1190232231463067, 32'sd-0.27136382597610675, 32'sd0.03564622100152204, 32'sd-0.02534059070812695, 32'sd-0.09226507249554326, 32'sd0.2481836405147952, 32'sd0.15506618638141015, 32'sd-0.04558325630102996, 32'sd-0.043152780551372574, 32'sd-0.17580680788702857, 32'sd-0.12975240213463685, 32'sd-0.0008703492813487804, 32'sd-0.000872333889030602, 32'sd0.15590437017625544, 32'sd0.3857217558936134, 32'sd-0.14826730217681786, 32'sd0.07473347328447404, 32'sd0.07755461129091411, 32'sd0.08809698041202968, 32'sd-0.2300404860191383, 32'sd-0.17689784050446178, 32'sd-0.043979658156686315, 32'sd-0.17423538128671595, 32'sd-0.16695994688496946, 32'sd0.17856441384979096, 32'sd0.04460685578854826, 32'sd0.11087703518971569, 32'sd-0.04225318202149157, 32'sd-0.0868598648696154, 32'sd0.062088953243450914, 32'sd0.03669427602876091, 32'sd0.12391757510961252, 32'sd-0.0691309659418636, 32'sd0.227518476131562, 32'sd-0.028912954724249533, 32'sd-0.04294122647668666, 32'sd-0.08698776187074322, 32'sd0.17984020824773284, 32'sd0.03458077431280889, 32'sd-0.05184825338545161, 32'sd0.2022502259116901, 32'sd-0.034933605809503915, 32'sd0.08151469803101909, 32'sd-0.10262439886629135, 32'sd-0.09776439073100873, 32'sd0.023901461133025118, 32'sd0.13377600595891925, 32'sd0.09612513425132953, 32'sd0.12090850826308712, 32'sd0.004498421911593788, 32'sd0.05057230442220217, 32'sd-0.29144111346538154, 32'sd-0.12429495624173358, 32'sd0.00840237328765869, 32'sd-0.03596473482656049, 32'sd0.05277731481199685, 32'sd-0.020334470867774585, 32'sd0.21041186229126063, 32'sd0.031162958632929342, 32'sd0.0015473470832326262, 32'sd-0.06871242483827607, 32'sd-0.16054082124910904, 32'sd0.23216374675623885, 32'sd-0.04827071187919016, 32'sd0.13019913072882394, 32'sd-0.17466755648447999, 32'sd0.01602799498671485, 32'sd0.1463850815250699, 32'sd0.18796744604788773, 32'sd0.0028905041699472823, 32'sd0.10328766177895733, 32'sd-0.059793769917016334, 32'sd0.21141145616582005, 32'sd-0.11810111145767313, 32'sd0.11731853139737032, 32'sd0.08598164797344222, 32'sd-0.23347335862528437, 32'sd0.11563820570446236, 32'sd0.14546993594030733, 32'sd-0.0830659717431911, 32'sd-0.019512390172488465, 32'sd-0.2554025262407493, 32'sd0.23062037178914127, 32'sd0.14787830320863674, 32'sd-0.22086116541751516, 32'sd0.2040410618306137, 32'sd0.006868344550945439, 32'sd-0.03611088188820081, 32'sd0.05571277209556439, 32'sd-0.19030062216644666, 32'sd-0.12675982359721646, 32'sd0.18953305095460185, 32'sd0.24820622295839986, 32'sd0.196974760825856, 32'sd0.03345550187970904, 32'sd0.167017706192906},
        '{32'sd-0.28060352399131444, 32'sd0.12417947469271177, 32'sd-0.12707641048460652, 32'sd0.14886923942757663, 32'sd-0.11245640985616036, 32'sd0.1381276386283418, 32'sd0.07080500612647322, 32'sd-0.09039036848051565, 32'sd-0.27142315517467996, 32'sd0.19057927854461496, 32'sd0.12152350342688933, 32'sd0.11477662876216985, 32'sd0.021618921900815005, 32'sd-0.11751769701238585, 32'sd0.034034158772163946, 32'sd-0.07830763610223589, 32'sd0.23014450832139424, 32'sd0.03572891054570344, 32'sd0.0035791424432308374, 32'sd-0.15758848276465898, 32'sd-0.19258903833554752, 32'sd-0.12503131299352882, 32'sd-0.26034851101875917, 32'sd0.005602749875050994, 32'sd0.17260210694666686, 32'sd0.14311629707274456, 32'sd0.05427374932307467, 32'sd-0.006742632727328567, 32'sd0.16506110312920952, 32'sd0.005360681605095413, 32'sd-0.09066375788239142, 32'sd0.14198607130901583, 32'sd-0.19568660171755756, 32'sd-0.01507561685979377, 32'sd0.1042377822279837, 32'sd-0.12892465279642992, 32'sd-0.24148844261011618, 32'sd0.13693508875589336, 32'sd-0.02473907057524971, 32'sd-0.2135964053428479, 32'sd0.004997461746834049, 32'sd-0.1186472401848023, 32'sd0.12905195986755183, 32'sd-0.10189838949708292, 32'sd-0.006655776135732462, 32'sd0.10467550098499626, 32'sd-0.20746826335285606, 32'sd-0.22344282122650405, 32'sd0.13011052777849547, 32'sd0.11387037134514931, 32'sd0.17046033493205262, 32'sd-0.1581229615923504, 32'sd0.0929395040786425, 32'sd0.040124532082694266, 32'sd0.13230144582919426, 32'sd-0.055338963643893416, 32'sd0.06678356092015615, 32'sd0.016627481839161698, 32'sd0.10186792860743638, 32'sd0.15262364615091967, 32'sd0.039169856367944865, 32'sd0.06719295112127308, 32'sd0.005667515391520679, 32'sd-0.07271132606064587, 32'sd0.01653256431886297, 32'sd-0.10415745008488132, 32'sd-0.14272595616522804, 32'sd0.03227587104696612, 32'sd0.04994648608922568, 32'sd0.13819376865261995, 32'sd0.1498942436831875, 32'sd-0.021977182146924203, 32'sd-0.08021963129435823, 32'sd-0.15577052121929344, 32'sd-0.05117347472703564, 32'sd0.11235902421995117, 32'sd-0.08328562129745083, 32'sd0.1624066081421054, 32'sd0.1989047566976893, 32'sd-0.050292378699927164, 32'sd-0.28144534114476977, 32'sd0.15632193471000205, 32'sd0.0895006187930222, 32'sd-0.2532301143184229, 32'sd0.20012327049797646, 32'sd-0.06562097191861821, 32'sd0.023308615771860275, 32'sd-0.024325638160697403, 32'sd0.015960189031938188, 32'sd-0.05602914739673578, 32'sd-0.13113637864930314, 32'sd0.06281044169136472, 32'sd-0.06799133390662539, 32'sd0.07521044952940423, 32'sd-0.03069118606948221, 32'sd-0.10610562039690097, 32'sd-0.1510579110868751, 32'sd-0.050678768418030935, 32'sd-0.033466451260479535, 32'sd-0.12149219823005368, 32'sd0.2114283835827421, 32'sd0.23877687093509006, 32'sd9.477552098358142e-05, 32'sd-0.24341529532162567, 32'sd-0.08766109074979807, 32'sd0.0048960548449841585, 32'sd-0.05597693702353088, 32'sd-0.1480173524444814, 32'sd-0.11690355345740204, 32'sd-0.15032600319927353, 32'sd0.1475544633451618, 32'sd-0.14202311294577058, 32'sd-0.15587775153590416, 32'sd-0.12499507953063554, 32'sd0.29467749834521695, 32'sd0.02664607295205598, 32'sd-0.0868786594845831, 32'sd-0.125319571129878, 32'sd0.06051407337252278, 32'sd-0.09336585100975547, 32'sd0.19117291584623786, 32'sd0.13523096208695096, 32'sd0.02994427226680538, 32'sd0.057747757420162006, 32'sd-0.012021980259177454, 32'sd0.04778959880537285, 32'sd0.0632392832416153, 32'sd0.09123551678715987},
        '{32'sd0.07031778092140042, 32'sd0.18288309356000945, 32'sd0.010012807937408589, 32'sd-0.02450005946546817, 32'sd0.23334043441722999, 32'sd0.2607357508034505, 32'sd-0.24286826409532053, 32'sd0.12601183020359263, 32'sd-0.09730953919734582, 32'sd0.10517984253451615, 32'sd0.052755658167937, 32'sd-0.036932169110684344, 32'sd0.029733914292463567, 32'sd-0.024417343510648906, 32'sd-0.07966886739898064, 32'sd-0.031226853344183188, 32'sd-0.07673625952870451, 32'sd-0.05915505221572816, 32'sd0.19818600361214717, 32'sd0.17004705495158035, 32'sd0.15256879218475888, 32'sd0.3459419050372023, 32'sd-0.0921409234871891, 32'sd0.1514600874821296, 32'sd-0.04167192063800042, 32'sd-0.06644996948171746, 32'sd-0.22285830270504342, 32'sd-0.2286289938859232, 32'sd-0.024735607770752302, 32'sd-0.0023354589211402933, 32'sd0.16361156099917876, 32'sd-0.11640713091034213, 32'sd-0.2995816265853071, 32'sd-0.050508697032672134, 32'sd0.07582636154431603, 32'sd0.1639050573942141, 32'sd0.07252716833090858, 32'sd-0.06124237354579071, 32'sd-0.24903183129309978, 32'sd-0.02866920134349755, 32'sd0.20957683841792332, 32'sd0.01773962851455979, 32'sd-0.16610935895653534, 32'sd0.00040396678674146463, 32'sd0.14436718736829077, 32'sd0.02792170657469366, 32'sd-0.1260249194592859, 32'sd0.10975704141603522, 32'sd0.003430865478650884, 32'sd0.15161432137270273, 32'sd0.20860257872097193, 32'sd-0.06448900323300806, 32'sd-0.032347022827974664, 32'sd-0.10503224418424809, 32'sd0.20567045779772275, 32'sd-0.13261701706101106, 32'sd-0.20607211077218357, 32'sd0.028717278793064172, 32'sd-0.01891982216910501, 32'sd0.16036692426769109, 32'sd-0.023769422311196792, 32'sd-0.0008008912141207589, 32'sd0.09184397950251519, 32'sd0.05505069479609141, 32'sd0.1550818707177843, 32'sd-0.1459143384298852, 32'sd-0.09517278179596483, 32'sd0.09305879979036266, 32'sd-0.08599847136332656, 32'sd0.10086745727297006, 32'sd-0.07085792046947943, 32'sd-0.13096998415480707, 32'sd0.08676516564421075, 32'sd-0.022472272178670684, 32'sd-0.05604945340362922, 32'sd-0.05147881893759971, 32'sd-0.173503815285886, 32'sd-0.03229493327049398, 32'sd0.15823139055849653, 32'sd0.05019498253962665, 32'sd-0.16406533059032816, 32'sd0.2072137441277403, 32'sd0.04201926387157047, 32'sd-0.03985796997197329, 32'sd0.01889085132987703, 32'sd0.02974355004995665, 32'sd-0.15043382621799703, 32'sd0.1452201620391728, 32'sd-0.0845362716196719, 32'sd-0.04160685086311638, 32'sd0.00782595093513723, 32'sd0.09366881243225182, 32'sd0.011885895761888941, 32'sd0.12603559072032355, 32'sd0.06291566777958653, 32'sd0.04703634600673222, 32'sd0.1665950173049541, 32'sd0.007283168627034632, 32'sd0.027432877032167336, 32'sd-0.15555423494900444, 32'sd0.19056950604741496, 32'sd0.10494210738408419, 32'sd-0.011127189512204866, 32'sd0.15303982080798806, 32'sd-0.1114852522610415, 32'sd0.16547264940061432, 32'sd0.09998893307125059, 32'sd-0.1326635122216051, 32'sd-0.034179305440814635, 32'sd0.08199907231476096, 32'sd0.09064161692570705, 32'sd-0.17084565740079002, 32'sd0.1566399382874324, 32'sd0.08826485046355105, 32'sd0.0153282723177789, 32'sd-0.21558449026847407, 32'sd0.23242614827973507, 32'sd0.012873772022212385, 32'sd0.020432899954622843, 32'sd-0.24690037206090454, 32'sd-0.07352112132318356, 32'sd0.12347822302610656, 32'sd0.11948127389292207, 32'sd0.0706761976379465, 32'sd0.11368593638686052, 32'sd0.24349411381765115, 32'sd-0.21736536517470031, 32'sd0.20125050684448356},
        '{32'sd0.09622275035460186, 32'sd0.0989015983907257, 32'sd0.0274072873550073, 32'sd0.1747653657294963, 32'sd0.1929818276251525, 32'sd0.0819086763022143, 32'sd-0.1875681690616536, 32'sd0.020609319356444365, 32'sd-0.10484259216390002, 32'sd0.09918208472813413, 32'sd-0.09428977881342457, 32'sd0.06981969214566425, 32'sd0.052578675792374865, 32'sd0.14965912073804133, 32'sd0.15244912954273257, 32'sd-0.11889534230631679, 32'sd-0.045950304321757486, 32'sd-0.007078688409665773, 32'sd0.2121040506605987, 32'sd0.09719661246027893, 32'sd0.008082835039396902, 32'sd0.19987555141711216, 32'sd0.12895320608696112, 32'sd0.11409764027709975, 32'sd-0.17385209742517255, 32'sd0.011546837978808008, 32'sd0.09037179394728401, 32'sd0.1386522047328418, 32'sd0.002137580893616131, 32'sd-0.23142259397999906, 32'sd-0.16612376233072773, 32'sd-0.06090865434099867, 32'sd0.09296776197316448, 32'sd-0.023251473599535586, 32'sd0.03157738248236455, 32'sd0.15790643116667144, 32'sd0.12822937525487932, 32'sd0.008662576803423506, 32'sd0.002006234291497846, 32'sd0.1963104095309515, 32'sd0.07239236868764039, 32'sd0.288061866568895, 32'sd0.15745886408751741, 32'sd-0.10943023521913313, 32'sd0.11301501362111194, 32'sd0.16899306248806584, 32'sd-0.3687290474182163, 32'sd0.22018953259945068, 32'sd-0.2426012726979581, 32'sd-0.16033955037259878, 32'sd-0.07925224314803607, 32'sd0.11288379450162662, 32'sd0.2165629977312835, 32'sd0.20099152183885005, 32'sd-0.058324760711319375, 32'sd-0.2692604781814382, 32'sd-0.06969850722052333, 32'sd-0.0945442388612388, 32'sd0.026575117371058672, 32'sd0.10984372829429037, 32'sd0.017447944624418003, 32'sd-0.021256604643855766, 32'sd0.05443212094491789, 32'sd0.052923622241606225, 32'sd0.09088373948397635, 32'sd-0.049154192639836905, 32'sd-0.1835902984958824, 32'sd0.042462688501523835, 32'sd0.1379100732505748, 32'sd0.2171361506306081, 32'sd-0.15440289822114728, 32'sd-0.28771888670446716, 32'sd-0.3409165437621842, 32'sd0.21385294457338366, 32'sd-0.26193181971733254, 32'sd-0.14849211024907083, 32'sd-0.23425081371713874, 32'sd-0.3331149616636346, 32'sd0.09594352570496917, 32'sd-0.11657980769585922, 32'sd0.042838510298660155, 32'sd0.0035977829732220176, 32'sd0.22374011229528773, 32'sd0.17651968909144164, 32'sd0.08126410191720025, 32'sd0.002959847312359741, 32'sd0.028037331829882575, 32'sd-0.12168094678370031, 32'sd0.1094034741568874, 32'sd0.008958352111850114, 32'sd-0.11563866229514763, 32'sd0.11941470964289035, 32'sd-0.17848426512891416, 32'sd0.24234546188966305, 32'sd-0.17105304378276312, 32'sd0.019917638274225883, 32'sd-0.06378088303515428, 32'sd0.11836638451605028, 32'sd-0.06708013243891775, 32'sd0.07490981437759542, 32'sd0.11368678582136825, 32'sd0.17334081287001973, 32'sd-0.06774921882261734, 32'sd0.1507781277150729, 32'sd-0.03738046723209661, 32'sd0.09035239615124153, 32'sd0.12092707056852389, 32'sd-0.14234291308384506, 32'sd-0.10046428811918576, 32'sd0.09918514725910248, 32'sd0.03564478714414918, 32'sd0.044905432077442374, 32'sd0.11729321110468913, 32'sd0.171820399948776, 32'sd-0.017675049140548217, 32'sd-0.1579732010569796, 32'sd0.13555071492685838, 32'sd-0.04756871935472286, 32'sd-0.09729746837715826, 32'sd0.11894274037252034, 32'sd0.04032560384463974, 32'sd-0.11106256366524336, 32'sd-0.09361480178691248, 32'sd-0.007305921590897141, 32'sd-0.07091264893359459, 32'sd0.1867623101384058, 32'sd0.20034207025558265, 32'sd-0.27944361829868836},
        '{32'sd-0.2109440536953244, 32'sd0.1131540658533114, 32'sd0.08120512292017938, 32'sd-0.08925070764819092, 32'sd-0.105174521191839, 32'sd0.15380376355028272, 32'sd0.04907146203301149, 32'sd0.1865383742283977, 32'sd-0.10053071575109869, 32'sd0.032308131923862025, 32'sd-0.20666105210866506, 32'sd-0.005723750231900902, 32'sd-0.10192256041667448, 32'sd-0.07603104362939067, 32'sd0.024724651240668492, 32'sd0.1351608173549326, 32'sd-0.162661944184012, 32'sd0.03440356340227308, 32'sd0.12085477943073289, 32'sd-0.0004382320386726242, 32'sd0.061899890091833616, 32'sd-0.01952823555437891, 32'sd0.10438570385589406, 32'sd-0.020872286078977568, 32'sd0.2858256228549075, 32'sd0.19659093155126486, 32'sd0.03534683636301718, 32'sd-0.12439123675949147, 32'sd-0.04977951656670517, 32'sd0.10380563204216277, 32'sd0.02818310333925888, 32'sd-0.20800264042596242, 32'sd-0.06959823447455281, 32'sd-0.14167187762336922, 32'sd-0.25773754339775573, 32'sd-0.0403605132465846, 32'sd-0.02832691758017165, 32'sd-0.19311681370108733, 32'sd0.1011548430983189, 32'sd-0.09099788142463104, 32'sd-0.03969857083312229, 32'sd-0.14204741485542846, 32'sd0.02257678036730265, 32'sd0.11014451524993062, 32'sd0.10959169569234493, 32'sd0.051253871053211, 32'sd0.011536752884684651, 32'sd0.20844624358803543, 32'sd0.04799720080130814, 32'sd0.05164497921302737, 32'sd-0.1296942708719476, 32'sd0.19574669045111823, 32'sd-0.058757715403335325, 32'sd-0.2786629633684859, 32'sd0.0024749847925067125, 32'sd0.27212226726886884, 32'sd-0.017602525815329423, 32'sd-0.050511204750833795, 32'sd0.15273353053274655, 32'sd-0.07414293178027036, 32'sd0.046210351024978544, 32'sd0.037379920440790824, 32'sd-0.22202624217709183, 32'sd-0.04554191294282993, 32'sd-0.09856855461854615, 32'sd0.007332512652958293, 32'sd-0.13286001772622894, 32'sd-0.24238742325692217, 32'sd-0.14674359960058378, 32'sd-0.22937406374236174, 32'sd0.08488530635561016, 32'sd0.045410680905975165, 32'sd-0.2284830708725665, 32'sd0.08204404998544408, 32'sd0.0927746208574383, 32'sd0.03299180902452843, 32'sd0.12590780341677327, 32'sd0.146188942200448, 32'sd-0.13126498153910376, 32'sd0.03697399987384998, 32'sd-0.27836300847015705, 32'sd0.03077175532505945, 32'sd0.12586984193716663, 32'sd0.06902042064794375, 32'sd0.05103133982183184, 32'sd-0.10365223663880795, 32'sd0.12397279278493098, 32'sd0.08704275551419603, 32'sd-0.2154573646281536, 32'sd0.16034405002387764, 32'sd-0.14800067237836517, 32'sd-0.028829535560628984, 32'sd0.05355502970555418, 32'sd-0.12774727738769034, 32'sd-0.22877649306903344, 32'sd-0.06457865704134719, 32'sd0.02087464381918811, 32'sd0.04748593960354255, 32'sd0.13099368060901936, 32'sd0.2196644434416415, 32'sd-0.08663411808709488, 32'sd-0.2086141287863504, 32'sd0.005470353235499036, 32'sd0.10474159941545126, 32'sd0.1334101100292218, 32'sd-0.10747593544444912, 32'sd0.14032919517957917, 32'sd0.11839985184592175, 32'sd0.04876296872287191, 32'sd-0.0004268103821981214, 32'sd0.07525560870553333, 32'sd0.17959893481913206, 32'sd0.14604174547675206, 32'sd-0.07559720569763824, 32'sd-0.20560570544291193, 32'sd-0.18670365419917043, 32'sd0.021215785470658454, 32'sd0.044765337777297284, 32'sd-0.004244247987735969, 32'sd0.24173062109920074, 32'sd0.10876172969512451, 32'sd0.20322683770226485, 32'sd-0.013134727938882746, 32'sd-0.15243042461279147, 32'sd-0.12824008278870358, 32'sd-0.13863938040998325, 32'sd0.14772589076352588, 32'sd0.0903088618679276},
        '{32'sd-0.07970118350998003, 32'sd-0.33005920816281004, 32'sd-0.06257478999077294, 32'sd0.21543435496681315, 32'sd0.08769307891743808, 32'sd0.06541634443449063, 32'sd-0.2914059154780329, 32'sd0.031657432120697, 32'sd0.20745542082952273, 32'sd-0.1586789959104216, 32'sd0.20114826214175743, 32'sd0.09111238897142275, 32'sd0.05606192264731042, 32'sd0.06654335326405465, 32'sd0.2318755625442408, 32'sd-0.0269450782048776, 32'sd0.2253370901746971, 32'sd0.13136951163514674, 32'sd0.020426814698416288, 32'sd0.16849810022015094, 32'sd0.02384410033104802, 32'sd0.11602587707561182, 32'sd0.0567113638554174, 32'sd-0.11485464462827545, 32'sd-0.020475849820432546, 32'sd-0.01691003029788059, 32'sd-0.031167143393738158, 32'sd-0.1120404990022284, 32'sd-0.1539900717675326, 32'sd0.08814592378787466, 32'sd0.29186428112598806, 32'sd0.04178180398356914, 32'sd-0.10041338828064188, 32'sd0.06291024464304865, 32'sd0.1813883721449228, 32'sd0.05644183484687994, 32'sd-0.17702181267690906, 32'sd-0.10787115841181838, 32'sd-0.19725149978043477, 32'sd0.18998232676227123, 32'sd0.05315490849499655, 32'sd0.06768131921595295, 32'sd-0.20796917226188408, 32'sd-0.026065758462882286, 32'sd-0.26968084502086304, 32'sd0.008236956159487926, 32'sd-0.07008322145799678, 32'sd-0.10560281485260425, 32'sd-0.131875443159628, 32'sd-0.16208817684782356, 32'sd-0.0808001034244683, 32'sd-0.04403813557993255, 32'sd-0.20721692630766253, 32'sd0.028587286655040362, 32'sd0.09856757197239584, 32'sd0.008506167041451696, 32'sd-0.15621258586994966, 32'sd-0.11173822806399814, 32'sd-0.2204231222254799, 32'sd0.12298354906707631, 32'sd-0.07033121009916966, 32'sd-0.1684579391894589, 32'sd0.11621659332786052, 32'sd0.14298947402480722, 32'sd-0.10126446217008177, 32'sd-0.08571287574258772, 32'sd0.2123528490257841, 32'sd-0.08848950988051361, 32'sd0.06235817760931684, 32'sd0.03782163558151918, 32'sd0.037531594585639136, 32'sd0.1627393409169993, 32'sd0.12399563496520169, 32'sd-0.0546754043011156, 32'sd0.18720937298888743, 32'sd0.06697761570332389, 32'sd-0.2197418171644131, 32'sd-0.012916217199210765, 32'sd-0.06800301684563154, 32'sd0.0957696934488929, 32'sd-0.10730060528066335, 32'sd-0.01845219503073271, 32'sd0.041477953325286115, 32'sd0.06447952867268256, 32'sd0.20207168425517116, 32'sd-0.2523611420623791, 32'sd-0.0551824351319944, 32'sd-0.1438161019870377, 32'sd-0.07388537615545235, 32'sd0.014281984878202396, 32'sd-0.12211643658433155, 32'sd0.058982815315855766, 32'sd0.0221508571854184, 32'sd0.13907228803032579, 32'sd-0.06690574149035565, 32'sd-0.16334601819472522, 32'sd0.018290514672246502, 32'sd0.13988876071768552, 32'sd0.1776633845751381, 32'sd-0.135978255380106, 32'sd0.0490137875910931, 32'sd0.1024153582644868, 32'sd-0.16179898279326857, 32'sd-0.019867561390379297, 32'sd-0.007165774241815675, 32'sd-0.3263535164173051, 32'sd-0.10805335836773255, 32'sd0.02214803258432132, 32'sd0.12114749972853865, 32'sd0.07173058977669255, 32'sd-0.15591069861628296, 32'sd-0.02069774003305199, 32'sd0.29437842359846544, 32'sd-0.3104444023573949, 32'sd-0.08537573753780298, 32'sd-0.10250798949147777, 32'sd0.13539808643658327, 32'sd-0.07819454075848152, 32'sd-0.010671853464635308, 32'sd0.11621109779434684, 32'sd0.11171881391271574, 32'sd0.14061865990116887, 32'sd0.1457732817472897, 32'sd-0.15109431462556622, 32'sd0.1065633187151967, 32'sd-0.06646853036690868, 32'sd-0.07965567128294264, 32'sd-0.0025473809121106298},
        '{32'sd0.1379680201229344, 32'sd-0.01665361360140971, 32'sd-0.15881869744030794, 32'sd0.3020436758736437, 32'sd0.2855729714518669, 32'sd-0.042473942370534326, 32'sd-0.12058010170279111, 32'sd-0.0338032246327929, 32'sd0.05218101023882166, 32'sd0.06117188239567652, 32'sd-0.021890137834160096, 32'sd-0.20094354285298036, 32'sd-0.07509378975370307, 32'sd-0.10330616145154779, 32'sd-0.19757392349780495, 32'sd-0.29165398801593045, 32'sd-0.26412807393135274, 32'sd0.02094465017563116, 32'sd-0.006483120290416099, 32'sd-0.1391199974493507, 32'sd0.1698891134935016, 32'sd0.06761047545864592, 32'sd0.22399911191944188, 32'sd-0.030406584931722765, 32'sd0.1303260001153635, 32'sd0.169707922064674, 32'sd0.10813807088333563, 32'sd-0.045846660025566165, 32'sd0.1047468138884961, 32'sd-0.417977359300505, 32'sd-0.05858899789689028, 32'sd0.12063886177065544, 32'sd-0.18710511638793298, 32'sd-0.04012781945611129, 32'sd-0.09318160160615031, 32'sd-0.1155541134374352, 32'sd0.216665634068524, 32'sd-0.21084696833328795, 32'sd0.004484733938516001, 32'sd0.06267781674158408, 32'sd0.027757551797123116, 32'sd-0.026940962825667877, 32'sd-0.024572864897960806, 32'sd-0.39076538068836153, 32'sd-0.10755836339851299, 32'sd-0.08416779769855026, 32'sd-0.2676473513474088, 32'sd0.047318039048049244, 32'sd0.03479486284336962, 32'sd0.18251137041037563, 32'sd-0.09293083605882017, 32'sd0.1857843336792958, 32'sd-0.04345085201333627, 32'sd0.21710494641412756, 32'sd-0.15970009944133853, 32'sd-0.07067972150011988, 32'sd-0.17493831687826275, 32'sd-0.18290888515994455, 32'sd-0.22707784554245553, 32'sd0.16355626876258375, 32'sd0.019454979803170323, 32'sd-0.008855659445240817, 32'sd-0.016391013129331642, 32'sd0.08505007053223451, 32'sd0.04170106491445916, 32'sd0.030618102072828366, 32'sd0.09835252270433797, 32'sd-0.013589451221857509, 32'sd-0.18223041462528006, 32'sd-0.022924617130231924, 32'sd-0.1002033164915474, 32'sd0.047152878715272885, 32'sd-0.22609280926947786, 32'sd-0.17624125192527348, 32'sd-0.2504942543492804, 32'sd0.26088853736265355, 32'sd0.002648716595624415, 32'sd-0.12067266701655886, 32'sd0.08466846887867334, 32'sd-0.03649592181762685, 32'sd-0.013524417858882134, 32'sd0.13271583392988404, 32'sd-0.10080254262830325, 32'sd-0.08575432094449893, 32'sd0.0838824650449486, 32'sd0.04677221443813097, 32'sd-0.18532602728194753, 32'sd-0.03129345358310142, 32'sd0.05335310693136388, 32'sd-0.32507332962402563, 32'sd0.1021583403072421, 32'sd-0.2182052027088327, 32'sd0.15211365475174837, 32'sd0.2027899382034827, 32'sd-0.06520388226361089, 32'sd0.10016652941286629, 32'sd0.013844953227173067, 32'sd0.14406530586541103, 32'sd0.03391836979844638, 32'sd-0.14852884660445398, 32'sd0.1812879138991943, 32'sd0.10696613038371927, 32'sd0.09045297857920817, 32'sd0.12478480219927056, 32'sd0.19726515421340027, 32'sd-0.06304736416521195, 32'sd-0.006517254609768282, 32'sd0.041100270173920116, 32'sd0.12345257237395965, 32'sd0.025843485311468746, 32'sd0.21706368782405602, 32'sd0.15226220592979187, 32'sd0.02381505541946743, 32'sd0.14749965189545822, 32'sd-0.22557913644870403, 32'sd0.06548708962203913, 32'sd0.04021750780670664, 32'sd0.13366228193516655, 32'sd-0.17546622469575848, 32'sd-0.09485020654757445, 32'sd-0.10713542174517089, 32'sd-0.07702471364882489, 32'sd-0.2340076574806151, 32'sd0.09606966777033929, 32'sd-0.03458876818630513, 32'sd0.09277578216096216, 32'sd-0.1647012171835572, 32'sd-0.22003264904626768},
        '{32'sd-0.014146025808691171, 32'sd0.2085314406351501, 32'sd-0.04289619009825946, 32'sd-0.17208843807219487, 32'sd-0.18649448014743986, 32'sd-0.14335964457911687, 32'sd0.1050439994688072, 32'sd0.21481559750278068, 32'sd0.06675321261027564, 32'sd0.037093477199397665, 32'sd-0.03840501593346974, 32'sd-0.07674162384159447, 32'sd-0.06406148779454025, 32'sd0.16296294196847894, 32'sd0.13485837767359357, 32'sd-0.029458228194640994, 32'sd-0.02713975896497556, 32'sd0.17899790093120316, 32'sd-0.06995961817787485, 32'sd0.0952894035083338, 32'sd-0.05067102085040421, 32'sd0.13889319873282385, 32'sd0.23479915460792278, 32'sd0.16336901520790773, 32'sd0.1642061767203883, 32'sd0.149896113646204, 32'sd-0.07373359631436735, 32'sd0.1101061211352278, 32'sd0.04037954533955882, 32'sd-0.004325577476361552, 32'sd0.08495835806588341, 32'sd0.1264846556287592, 32'sd-0.03330046050883115, 32'sd0.024360965958151338, 32'sd-0.07136238416578572, 32'sd0.038183040922046205, 32'sd-0.07247950310269402, 32'sd0.20394971087905425, 32'sd0.11564749716430472, 32'sd0.09163119906529552, 32'sd-0.22836707223873323, 32'sd-0.3086432471181124, 32'sd-0.16150625442383137, 32'sd-0.08579643720931537, 32'sd-0.314397271982058, 32'sd-0.11702754105871606, 32'sd0.16602248039581813, 32'sd0.11584231349422398, 32'sd-0.1161823050732022, 32'sd-0.14847860273931587, 32'sd0.11957167196340299, 32'sd-0.09872388339775719, 32'sd-0.15506489883596467, 32'sd0.06707246164488109, 32'sd0.38033765503898825, 32'sd-0.013772079934819641, 32'sd0.12420414153443374, 32'sd-0.023170603803359505, 32'sd0.10986314424520971, 32'sd0.07269130543508014, 32'sd0.04964895084938239, 32'sd-0.28499117851202543, 32'sd-0.0436077241540402, 32'sd-0.1849756571941903, 32'sd-0.12621909419110766, 32'sd0.006799675589396278, 32'sd-0.2169645305393021, 32'sd-0.1170516033454532, 32'sd0.13499837005748688, 32'sd-0.2163074899302213, 32'sd-0.17031350957737845, 32'sd-0.024159530108099014, 32'sd0.10831073702264124, 32'sd-0.20286890528379636, 32'sd0.010588920564385892, 32'sd0.036928974873133555, 32'sd0.08141937915279543, 32'sd0.04366382408431808, 32'sd-0.2135909525562721, 32'sd0.19762441211945017, 32'sd-0.09322078141012516, 32'sd0.18492919604191901, 32'sd0.04459618888823948, 32'sd-0.17603300601259703, 32'sd-0.11498264301023724, 32'sd0.053093962525602896, 32'sd0.09759126190550155, 32'sd0.2570383824669631, 32'sd-0.2016922876928038, 32'sd0.1374658328468221, 32'sd0.14077975051878858, 32'sd-0.04710370729045995, 32'sd0.21543618476501783, 32'sd-0.17974664345996882, 32'sd0.1032118134936366, 32'sd-0.14262270456494244, 32'sd0.13113642916725585, 32'sd-0.16597849985189125, 32'sd0.2398599054069721, 32'sd-0.04495842409988396, 32'sd0.0007016260409384573, 32'sd0.1737155851639222, 32'sd-0.2180062104784241, 32'sd-0.18140042374822582, 32'sd0.07151683477994424, 32'sd0.03645279098216084, 32'sd-0.09413745258403086, 32'sd0.11598578087719078, 32'sd0.0022560573291964836, 32'sd-0.235085345267184, 32'sd-0.08687384937909548, 32'sd-0.2973334888331643, 32'sd0.030232928509834105, 32'sd0.014294375418443285, 32'sd-0.09905670465888874, 32'sd0.2013382726200191, 32'sd-0.02434232747698675, 32'sd0.21700600836694967, 32'sd0.08438296294873597, 32'sd0.11377734623744787, 32'sd-0.09195777156454987, 32'sd-0.01885550167657027, 32'sd-0.05134167602438419, 32'sd0.11269699675847712, 32'sd0.04289162166962784, 32'sd-0.13347346022838052, 32'sd-0.11971149292378154, 32'sd-0.0030350341510345254},
        '{32'sd0.1113701453667729, 32'sd0.18941676444557962, 32'sd-0.17844724013483684, 32'sd-0.11693848650911542, 32'sd0.031189527591412296, 32'sd-0.08961383920781324, 32'sd-0.26620450956873054, 32'sd0.04798986419499786, 32'sd0.03168505954836458, 32'sd0.15514856674191163, 32'sd0.05990219964927756, 32'sd-0.12234386059111066, 32'sd0.2476924392969135, 32'sd0.07652204987983095, 32'sd0.16646326371621617, 32'sd-0.26867737074210885, 32'sd0.26567340090557934, 32'sd0.0032835398425488894, 32'sd0.012947809101297727, 32'sd0.01958632962895276, 32'sd-0.02036622127018347, 32'sd-0.14964264534289334, 32'sd0.0994791585484714, 32'sd-0.16460060119296843, 32'sd0.09605291844705277, 32'sd-0.1680223481907282, 32'sd0.13278968491260276, 32'sd-0.04264411198868085, 32'sd-0.08002290703822267, 32'sd0.20052076593330181, 32'sd0.1218183176922181, 32'sd-0.026075879548194708, 32'sd-0.15392656659262388, 32'sd-0.02214651292772515, 32'sd0.07236315726811424, 32'sd-0.2176186208870718, 32'sd0.19551616836805022, 32'sd0.07262637406439587, 32'sd0.15668994471123196, 32'sd-0.20705494292989077, 32'sd-0.15947574010876367, 32'sd-0.16058903078355244, 32'sd-0.1449081592818639, 32'sd0.23538586213711757, 32'sd-0.09880197575250994, 32'sd-0.14695188346030413, 32'sd0.20038095233564399, 32'sd0.06873220239673442, 32'sd-0.18975447196699663, 32'sd0.026602903767180948, 32'sd-0.13284776688778885, 32'sd0.07653966169166246, 32'sd0.2398003005878075, 32'sd-0.21254794700248686, 32'sd-0.2525212182814109, 32'sd-0.0953010631535735, 32'sd-0.07164626850976866, 32'sd0.11547227293423327, 32'sd-0.170656999178572, 32'sd-0.17055590145221447, 32'sd0.17953899182761263, 32'sd0.0969902752640618, 32'sd-0.09168215915123303, 32'sd0.10758962897736629, 32'sd-0.05675881330675213, 32'sd0.13394143504266978, 32'sd0.12065175570266498, 32'sd-0.17713671373356493, 32'sd-0.0324772229801441, 32'sd0.08131037019936328, 32'sd0.06297457480296417, 32'sd-0.04947581156752847, 32'sd0.009603496927010175, 32'sd0.19816855041730286, 32'sd0.11551844571573607, 32'sd0.17149591097371833, 32'sd-0.012113286732506823, 32'sd0.008046168057064028, 32'sd-0.15467442943660303, 32'sd-0.1590546229193791, 32'sd-0.08553143779445306, 32'sd-0.05098815202431051, 32'sd0.09168174003865562, 32'sd0.003909003778377015, 32'sd-0.04047176717850877, 32'sd-0.049081476314629724, 32'sd0.15830016286383175, 32'sd0.12210597447211448, 32'sd-0.1177357546884603, 32'sd-0.22079528810489243, 32'sd0.22419792145066306, 32'sd0.004816031849181646, 32'sd-0.08170098365486478, 32'sd-0.1756292261302256, 32'sd-0.19501701715864045, 32'sd0.029300472047024628, 32'sd-0.36063944481106547, 32'sd0.14455627613805885, 32'sd-0.1005297269393348, 32'sd0.13129015099004435, 32'sd0.156426498608931, 32'sd0.21793254369601145, 32'sd-0.036444655895004556, 32'sd-0.020299805936879686, 32'sd-0.21757552953140807, 32'sd0.06349282317414219, 32'sd0.07026465907037494, 32'sd-0.044627368714745326, 32'sd-0.03861303477816885, 32'sd0.04017709921439397, 32'sd-0.11808423465742217, 32'sd0.13481811002718952, 32'sd-0.1395812602611448, 32'sd0.0622334918857842, 32'sd-0.13519944664517744, 32'sd0.10988513286481648, 32'sd-0.059709220423090556, 32'sd-0.12614384759472097, 32'sd0.10240999331460589, 32'sd-0.1271442184529824, 32'sd0.06337650420983315, 32'sd-0.09831304312196729, 32'sd0.037045514572015506, 32'sd-0.08825058461648802, 32'sd-0.21811326716697998, 32'sd-0.018588960317767522, 32'sd0.09943816429237844, 32'sd0.11857812161264261},
        '{32'sd0.005320443301173771, 32'sd-0.2061205420608775, 32'sd0.06585234098937381, 32'sd-0.13825988198448455, 32'sd0.08853498281664607, 32'sd-0.007487675297579787, 32'sd0.23062362494157007, 32'sd-0.06470434414419224, 32'sd0.11901098894615676, 32'sd0.042586366327798275, 32'sd0.07046729385751321, 32'sd0.1843321677438639, 32'sd-0.17878987391377868, 32'sd0.1351253561540518, 32'sd-0.03643465518662514, 32'sd-0.16029401884481184, 32'sd0.15000973417970279, 32'sd0.15579300741777213, 32'sd-0.025417070085442785, 32'sd-0.14277238282299176, 32'sd0.02775640129329202, 32'sd-0.15030847158528052, 32'sd0.07405889176431202, 32'sd0.07677983570948173, 32'sd0.16531335564081073, 32'sd-0.060051778988022254, 32'sd0.04723081211919356, 32'sd0.14628002676113364, 32'sd-0.000885382372485997, 32'sd-0.006575804640102162, 32'sd0.08560780174628714, 32'sd0.018649422944944732, 32'sd-0.08500601701872167, 32'sd-0.1550278941231016, 32'sd-0.10427016971377594, 32'sd0.04004443356986279, 32'sd-0.13360102976452926, 32'sd0.13145836308846814, 32'sd-0.07299691691832927, 32'sd-0.0008271588788195307, 32'sd0.17167513347166555, 32'sd-0.18125488557369207, 32'sd0.04543647136628449, 32'sd0.17917046464325825, 32'sd-0.292383427200315, 32'sd0.1425317786660963, 32'sd0.08178766989472926, 32'sd0.0917224054868679, 32'sd0.01070350440147739, 32'sd-0.09740070005712191, 32'sd0.16123793972946782, 32'sd0.041468386104099246, 32'sd-0.18805447559154814, 32'sd0.12244941449528361, 32'sd0.024566809604923013, 32'sd0.170407698802525, 32'sd-0.11735135525827588, 32'sd0.204202751975778, 32'sd0.1579139353071361, 32'sd-0.06366893103615667, 32'sd-0.07249143601319274, 32'sd-0.2852040360058721, 32'sd-0.05908596180557615, 32'sd0.1658284332416117, 32'sd-0.09602483600193643, 32'sd0.054423349930256965, 32'sd0.17858054812630447, 32'sd0.2184943317437912, 32'sd-0.08072028647451408, 32'sd0.04866391171002818, 32'sd0.0963671839452084, 32'sd-0.038159499947829384, 32'sd-0.06707189387659984, 32'sd0.06463473623670216, 32'sd0.20877142554145062, 32'sd0.1871344123003396, 32'sd-0.17933179860599288, 32'sd-0.03676981980142796, 32'sd-0.11615207552658346, 32'sd-0.008443293959726962, 32'sd0.16932211927843124, 32'sd0.05239540214575486, 32'sd-0.2102380137370182, 32'sd0.06728022831775296, 32'sd-0.2122707103637739, 32'sd0.12710629570546889, 32'sd0.10170853699163707, 32'sd0.0065426332434593585, 32'sd-0.18369497058914305, 32'sd0.07785407222407545, 32'sd0.2113038080785981, 32'sd-0.021096864013040385, 32'sd0.12159353544441791, 32'sd-0.19792028611906617, 32'sd0.1892905661175911, 32'sd0.0583023960840518, 32'sd0.03440429615292557, 32'sd0.18810315492623178, 32'sd0.09035798427795348, 32'sd-0.017213717550863854, 32'sd0.00317801625537658, 32'sd0.20364558120398019, 32'sd-0.19350017786303317, 32'sd0.019513945249982536, 32'sd0.07076554855728567, 32'sd0.16111365374530726, 32'sd-0.034537544958395505, 32'sd-0.06095468972857607, 32'sd0.1022667851313789, 32'sd0.01596939397812447, 32'sd-0.04018118687702544, 32'sd0.09673263133818193, 32'sd0.24460570215459257, 32'sd-0.0734618008781218, 32'sd-0.04656472099303353, 32'sd0.09645993649517548, 32'sd-0.053230932740123325, 32'sd-0.1841523350410677, 32'sd0.2186961211836596, 32'sd-0.027698311194830516, 32'sd0.16450219274595415, 32'sd0.05797216992136884, 32'sd-0.123582939335422, 32'sd0.013837807416530654, 32'sd-0.0161270923949011, 32'sd0.07215935875274632, 32'sd-0.025534116424879332, 32'sd-0.19189894625220336}
    };

    localparam logic signed [31:0] layer1_biases [0:63] = '{
        32'sd0.07890242738825, 32'sd0.016901702800579798, 32'sd-0.15014795818333584, 32'sd-0.03773399763928362, 32'sd-0.02335163209332366, 32'sd-0.028904161017689552, 32'sd0.13915590369284203, 32'sd0.16934301555395667, 32'sd-0.02648637106865187, 32'sd0.06134790165228979, 32'sd-0.11911536129996808, 32'sd-0.19549658382751603, 32'sd0.10062707232392605, 32'sd-0.06396620846094381, 32'sd0.13870075843504764, 32'sd-0.029957591487481755, 32'sd-0.10505235882556203, 32'sd0.0008832333040850178, 32'sd-0.029594003406838376, 32'sd0.19934670057316342, 32'sd-0.030011266795953076, 32'sd-0.09143925328593736, 32'sd0.18832764124717935, 32'sd-0.03763855860867775, 32'sd-0.186975455181606, 32'sd0.07695183865415899, 32'sd0.1813521093062877, 32'sd-0.002081270001533263, 32'sd-0.07990881466096862, 32'sd-0.0797459505044078, 32'sd0.0022282339924661956, 32'sd-0.09873633652602486, 32'sd-0.1545077916434072, 32'sd0.05483396920838122, 32'sd0.148963750272084, 32'sd-0.09094519932995161, 32'sd0.06898241029298917, 32'sd0.19174849331554683, 32'sd0.22205209139680288, 32'sd-0.16287873244198078, 32'sd0.011230165681501038, 32'sd0.1836077462550824, 32'sd0.06553872060226211, 32'sd-0.157732309977709, 32'sd0.15740995015352255, 32'sd0.17158420434875002, 32'sd-0.2292678853771437, 32'sd0.04275906162240555, 32'sd0.2274245398521201, 32'sd0.042238603200310615, 32'sd-0.0004689291796547292, 32'sd0.150551428204761, 32'sd-0.12349043340015266, 32'sd0.07835389338504516, 32'sd0.07322602169538493, 32'sd-0.035051846662123756, 32'sd0.18427974147581375, 32'sd0.012053758082939353, 32'sd0.010283753506129487, 32'sd-0.09395530588501491, 32'sd0.13958006651041208, 32'sd0.06084110633277807, 32'sd0.22129072062303287, 32'sd-0.08347651283288059
    };

    //Layer 2: 64 inputs, 10 neurons
    localparam logic signed [31:0] layer2_weights [0:9][0:64] = '{
        '{32'sd0.19141445069845722, 32'sd-0.05473271130248055, 32'sd-0.0379756305276999, 32'sd0.34271360463802164, 32'sd-0.1354344950675868, 32'sd0.10277262326909924, 32'sd-0.49534343317103563, 32'sd0.2287555894399951, 32'sd0.3135453048358562, 32'sd0.23142019219926457, 32'sd-0.32255277426722956, 32'sd-0.03863944626627424, 32'sd-0.4636078876939725, 32'sd0.0978926772432343, 32'sd-0.1657613732003654, 32'sd-0.17482918990295324, 32'sd-0.34519691078173503, 32'sd-0.3841873355992827, 32'sd-0.37562192225328417, 32'sd-0.4082344392014307, 32'sd0.23858015077378442, 32'sd-0.13151075991534783, 32'sd0.1548179143838379, 32'sd0.21269142677264974, 32'sd0.08394754461393758, 32'sd-0.3443348842868656, 32'sd-0.03943947630827211, 32'sd-0.13526190937258717, 32'sd0.12392195581793976, 32'sd-0.3347147369028981, 32'sd-0.34604937675940467, 32'sd0.2253167039190944, 32'sd-0.3124462758679872, 32'sd-0.3419081998161168, 32'sd-0.42025728817482694, 32'sd-0.30094943749068065, 32'sd-0.21899470362317108, 32'sd-0.33745388472379434, 32'sd0.1557763260503133, 32'sd-0.23468662299715737, 32'sd0.11439711603557642, 32'sd0.23310281733200058, 32'sd0.12465101360209803, 32'sd0.07794379852240789, 32'sd-0.3717372596581085, 32'sd0.2123499259893269, 32'sd-0.2942434727956893, 32'sd-0.41409446945832495, 32'sd-0.1254864884484945, 32'sd0.315792258425798, 32'sd0.25417430396107715, 32'sd0.3589896388956954, 32'sd-0.3800612716866141, 32'sd0.0025484076712958864, 32'sd-0.1589676796503928, 32'sd0.2634774482167261, 32'sd0.3428968829618216, 32'sd0.2826894553681636, 32'sd-0.18322423985920058, 32'sd0.186023173192589, 32'sd0.34577349458862616, 32'sd-0.48618866762902396, 32'sd-0.37278595050161994, 32'sd0.03659408886858046},
        '{32'sd0.13945558979464406, 32'sd0.10431937664737424, 32'sd-0.19088106324472948, 32'sd0.25722108351487005, 32'sd0.23372339963781982, 32'sd0.0027850276619740266, 32'sd-0.05299942690962679, 32'sd-0.08490413447325017, 32'sd-0.051968829742950196, 32'sd-0.35903614305459436, 32'sd-0.33778213828141146, 32'sd0.12632504410482306, 32'sd-0.021398664403088886, 32'sd-0.41639023048486756, 32'sd-0.3337642219415796, 32'sd0.2932784979561823, 32'sd0.32414074700187423, 32'sd-0.3197853988638006, 32'sd-0.24282589790046435, 32'sd0.26828494635557504, 32'sd0.3725544103612544, 32'sd-0.27603045800354603, 32'sd0.010592968921293262, 32'sd0.31440785033583357, 32'sd0.3816828009961947, 32'sd0.048538649169251796, 32'sd-0.3311368985966095, 32'sd0.02246289794255768, 32'sd-0.337686516734316, 32'sd0.336436934632465, 32'sd-0.3941674023063687, 32'sd0.19511131909208126, 32'sd0.08201432259158353, 32'sd-0.14166089062400142, 32'sd-0.25760775109339723, 32'sd-0.5163756409437407, 32'sd-0.3248173271827846, 32'sd0.13285380287102724, 32'sd-0.38266274261346916, 32'sd-0.270955141019226, 32'sd0.14782047551194766, 32'sd-0.294438859879701, 32'sd0.31452149349539593, 32'sd-0.05720762926694285, 32'sd-0.1495003723136737, 32'sd-0.43035656530760247, 32'sd0.2263659980345605, 32'sd-0.1925615909731174, 32'sd-0.4825335205139854, 32'sd-0.09913319936750266, 32'sd-0.025782656859380425, 32'sd0.21527681723301703, 32'sd-0.08316039134630195, 32'sd-0.1924447179781557, 32'sd0.11372044025622698, 32'sd0.11996266775495969, 32'sd0.13210941065059134, 32'sd-0.2931408044279939, 32'sd0.35316440054184345, 32'sd0.06334662562928882, 32'sd-0.29175809417375864, 32'sd0.4090221019060916, 32'sd-0.27403218700853904, 32'sd-0.13041057926152402},
        '{32'sd0.030267494907296875, 32'sd-0.127042272610891, 32'sd0.36759403962537385, 32'sd0.19378023409781855, 32'sd0.15860272458626054, 32'sd-0.3508822745177931, 32'sd0.23437505977724918, 32'sd0.24133806503348967, 32'sd-0.08041043558703109, 32'sd-0.20512790283827906, 32'sd-0.22714541322507623, 32'sd0.28696339128292847, 32'sd-0.14284897581061035, 32'sd-0.006920672849142421, 32'sd0.09209085699508456, 32'sd0.042600035928536895, 32'sd-0.27586528316327996, 32'sd0.10277148636857136, 32'sd0.16345245548373477, 32'sd0.3075722525420259, 32'sd-0.12683137636204853, 32'sd-0.16625206815921417, 32'sd-0.17381293978913226, 32'sd-0.14073884908596382, 32'sd-0.16897515867386892, 32'sd-0.27774888480943327, 32'sd-0.009948452625822906, 32'sd-0.4671146229352994, 32'sd0.11629741652162942, 32'sd-0.16990364379714104, 32'sd0.02854619756248002, 32'sd0.19640945523819367, 32'sd-0.16249988097617418, 32'sd-0.2896764184824139, 32'sd-0.3145095706392847, 32'sd0.03084267648493712, 32'sd0.08572902394066598, 32'sd-0.16537855804510385, 32'sd-0.09000718837050659, 32'sd0.2154894272544899, 32'sd-0.3649967017697578, 32'sd0.0023769207761900157, 32'sd-0.323549064160835, 32'sd0.2684163165634101, 32'sd0.010542167507526823, 32'sd0.1302617061789021, 32'sd-0.16412432136440422, 32'sd0.3636326418591278, 32'sd0.23830579913538627, 32'sd-0.011510497094255093, 32'sd0.3689240269109286, 32'sd-0.008111690852714397, 32'sd0.05331777913279486, 32'sd0.33689019669488507, 32'sd-0.19393860676522656, 32'sd-0.31867237927737513, 32'sd-0.004459260460829312, 32'sd0.03749107213287588, 32'sd0.19246569546075287, 32'sd-0.089589962882438, 32'sd-0.35188985911116866, 32'sd-0.13322535764010363, 32'sd0.199549433020255, 32'sd-0.07123445220660417},
        '{32'sd0.05749502683837287, 32'sd0.026582039123984505, 32'sd0.20717426905435068, 32'sd0.11356654533671147, 32'sd-0.45382946680765585, 32'sd0.12695667109511447, 32'sd-0.3142981045251369, 32'sd0.2805469754301725, 32'sd0.139458771308345, 32'sd-0.08124945587606838, 32'sd0.09062284122651627, 32'sd-0.13291018007054595, 32'sd-0.3194554785628693, 32'sd0.03624516944426584, 32'sd-0.005174267947329018, 32'sd-0.29055262021918243, 32'sd0.28741456415992517, 32'sd0.15686960695493699, 32'sd0.31045513413689385, 32'sd-0.09067313137131248, 32'sd-0.357989651268917, 32'sd-0.20783580277040292, 32'sd-0.3857127702154846, 32'sd0.03388467986887699, 32'sd-0.06020204727677744, 32'sd0.33328558686388055, 32'sd-0.2552111230995789, 32'sd0.2183910050048773, 32'sd0.25394390943115935, 32'sd0.24959925549201972, 32'sd0.2963952414585705, 32'sd-0.31656076389751187, 32'sd-0.12284946019086884, 32'sd-0.24645289058909114, 32'sd0.28110397520949054, 32'sd0.18514410434507458, 32'sd-0.3753942421858096, 32'sd-0.008144136582259756, 32'sd0.025770170783660565, 32'sd-0.13108917161764433, 32'sd-0.1645325183309439, 32'sd0.32196012779396577, 32'sd0.02933471884118189, 32'sd0.20051265164515902, 32'sd-0.1715594440097634, 32'sd0.3341999869853428, 32'sd-0.3001773520307309, 32'sd-0.10126535074905757, 32'sd0.18235345310072335, 32'sd-0.12437864762947252, 32'sd-0.344490384124856, 32'sd0.11380379538261384, 32'sd-0.25415253941673777, 32'sd-0.1065822415161939, 32'sd0.03698461071763806, 32'sd0.15869670226974295, 32'sd-0.1995803896973124, 32'sd-0.39391169736807885, 32'sd-0.18173638397618835, 32'sd0.041465310424306005, 32'sd-0.24312812677389276, 32'sd0.36809918361142047, 32'sd-0.10535704463948836, 32'sd0.3267380646856233},
        '{32'sd-0.057496605198111624, 32'sd-0.06924997622177553, 32'sd-0.0679165068971247, 32'sd-0.5693254213455768, 32'sd0.2487737887428959, 32'sd-0.12709821211426944, 32'sd-0.4111833803800929, 32'sd-0.5102090010973817, 32'sd0.04302200287007302, 32'sd0.07960820038543394, 32'sd0.21020883175628022, 32'sd-0.12860428634236387, 32'sd0.3353586913522529, 32'sd-0.34278927536887116, 32'sd-0.442509659310754, 32'sd0.20277331431417348, 32'sd-0.27811678998039596, 32'sd0.04486137490309698, 32'sd0.15777471175879426, 32'sd-0.01103073197189138, 32'sd0.29137094884106146, 32'sd-0.12075931383207025, 32'sd-0.21049740935423922, 32'sd0.3620522969249711, 32'sd-0.06403741686652513, 32'sd-0.4473199306318343, 32'sd0.04235316377832709, 32'sd0.3292572115415764, 32'sd-0.2877199022548809, 32'sd0.168663267372474, 32'sd0.039975865340506546, 32'sd0.18646301828691142, 32'sd0.21260386980881507, 32'sd0.3288888330262427, 32'sd0.051902177949378264, 32'sd0.05744328374610806, 32'sd-0.02086178046659716, 32'sd0.01947447069342589, 32'sd0.3119507315286304, 32'sd-0.2107218123493312, 32'sd0.23351031521505, 32'sd-0.47575895494482145, 32'sd-0.06675694425577006, 32'sd0.1419564268296635, 32'sd-0.48598632418285365, 32'sd-0.18543512316729482, 32'sd-0.3747357265484507, 32'sd0.11699455161876027, 32'sd0.26174279372984566, 32'sd0.08969217664873692, 32'sd0.19529051259481214, 32'sd-0.4154020420086673, 32'sd0.03748322673222059, 32'sd0.27924994626280053, 32'sd-0.24289609777236645, 32'sd-0.41110637375204856, 32'sd-0.02724246611033031, 32'sd-0.14997255381503144, 32'sd-0.018439358103918217, 32'sd0.3536164774955274, 32'sd-0.06651257064439837, 32'sd-0.012875001860130759, 32'sd0.20357342397977546, 32'sd0.11962337685515749},
        '{32'sd-0.3852750984849929, 32'sd0.029852054115761466, 32'sd-0.0811079657691721, 32'sd-0.03279028905053023, 32'sd0.05077888589011638, 32'sd0.130197009921609, 32'sd0.24433737118503027, 32'sd0.12485224907285233, 32'sd-0.20489095707156182, 32'sd-0.04893169264697161, 32'sd0.1424610631033282, 32'sd0.05890609245804754, 32'sd0.16548610223118213, 32'sd0.3398480438611997, 32'sd-0.07959725819688182, 32'sd-0.3329913016031232, 32'sd-0.4023488058946217, 32'sd-0.0023430587448545633, 32'sd-0.39050530748668655, 32'sd-0.33321363818633526, 32'sd-0.012260770834893587, 32'sd0.2929262160361813, 32'sd0.0384682255533624, 32'sd0.22161613758516424, 32'sd0.027191910775293544, 32'sd0.22778857180714768, 32'sd-0.495489185816338, 32'sd-0.07896016694525528, 32'sd-0.07575176465193391, 32'sd-0.4573577549901302, 32'sd0.24310431933745552, 32'sd-0.2181358490976818, 32'sd0.1903109324517183, 32'sd0.075965074424552, 32'sd0.058676950660471565, 32'sd0.13484031409692693, 32'sd-0.08457903457820068, 32'sd0.37478230830437637, 32'sd-0.5628681000944369, 32'sd0.36005934390658495, 32'sd-0.03476605161013679, 32'sd-0.0685369793863901, 32'sd0.37711079583377904, 32'sd0.25113680165876684, 32'sd-0.09332757348844366, 32'sd0.07654572037554509, 32'sd0.1738625731407075, 32'sd-0.39935541354816945, 32'sd0.26093359926338094, 32'sd0.23361188994561025, 32'sd-0.4124823414924174, 32'sd0.10528472649494852, 32'sd-0.09481978811171755, 32'sd0.01037300630802922, 32'sd0.23630776507892345, 32'sd-0.18960914966779013, 32'sd-0.3953266643275367, 32'sd-0.21343044069411607, 32'sd0.24384007202898206, 32'sd-0.32152982135549946, 32'sd0.14916040038827186, 32'sd-0.2558438318423902, 32'sd0.2617818393356741, 32'sd-0.2672646826820461},
        '{32'sd-0.34155993020574954, 32'sd0.24818269496833167, 32'sd0.042580206590230686, 32'sd0.0361391088861395, 32'sd0.24855731458132346, 32'sd0.19215811360376978, 32'sd-0.0988792633128899, 32'sd-0.18467762778701194, 32'sd0.29825786816374633, 32'sd0.3666050292444358, 32'sd-0.24724152859068896, 32'sd0.0044043934698866655, 32'sd0.15521171897156316, 32'sd0.26856003881298707, 32'sd0.05511761379338089, 32'sd-0.021162158670727956, 32'sd-0.2056900775297141, 32'sd-0.07439638742374563, 32'sd-0.34834594506925304, 32'sd-0.03923159150189144, 32'sd-0.02766202781568702, 32'sd-0.31369521566416136, 32'sd0.11225575028209327, 32'sd0.1165888557112309, 32'sd0.44178355222974647, 32'sd-0.04736479518780336, 32'sd-0.303516587851339, 32'sd-0.010402889974586028, 32'sd0.30131648351100543, 32'sd0.2484123596189563, 32'sd0.14019030103063954, 32'sd-0.19721705925759478, 32'sd-0.26339979353217324, 32'sd0.24118869802732382, 32'sd-0.40962610365631685, 32'sd0.2944987208580412, 32'sd0.276443210618532, 32'sd-0.08993403068664793, 32'sd0.07148206532759646, 32'sd-0.3179429057423349, 32'sd-0.32907967400175875, 32'sd0.24220219663834983, 32'sd0.11189725592302426, 32'sd0.21364574465745922, 32'sd-0.3662602562920978, 32'sd-0.1893498784661194, 32'sd0.20822289436469746, 32'sd-0.14958015222334023, 32'sd-0.35553143750015004, 32'sd0.15974908209576988, 32'sd0.25282003948010434, 32'sd-0.23651267122010175, 32'sd0.175546563240566, 32'sd0.16756053573224747, 32'sd-0.2911347916151833, 32'sd-0.11455975893696092, 32'sd-0.3171369094380908, 32'sd0.30950519222476525, 32'sd-0.2787705981694796, 32'sd-0.28596429583408517, 32'sd-0.015254453762470048, 32'sd0.137047212016339, 32'sd0.041306757618595966, 32'sd-0.08476874813584076},
        '{32'sd-0.08236513754240248, 32'sd0.2630490879184157, 32'sd0.14826105493257696, 32'sd0.19619860166132586, 32'sd0.010261307582093801, 32'sd-0.38438683139965185, 32'sd0.2575568506174208, 32'sd-0.2774258190656574, 32'sd-0.34664062009377056, 32'sd0.04008961884762732, 32'sd0.3415228987713681, 32'sd0.0436417749324023, 32'sd-0.23007580145610323, 32'sd-0.26247817426039677, 32'sd-0.321036978245998, 32'sd0.20327133153223198, 32'sd0.2890588175076209, 32'sd-0.12502588565888337, 32'sd0.23115682982569216, 32'sd0.1603765120127169, 32'sd-0.0796525812927751, 32'sd-0.016594696498030394, 32'sd-0.3226980509883961, 32'sd0.15497497151694725, 32'sd-0.2857263506175931, 32'sd-0.09797150486065234, 32'sd-0.09360982138503643, 32'sd0.05799075060436488, 32'sd0.23177162393581144, 32'sd-0.31137456000856756, 32'sd-0.3320891753572984, 32'sd0.0292698182154449, 32'sd-0.14566095840770302, 32'sd0.1718350648952016, 32'sd0.06898412444940842, 32'sd-0.01728818852243991, 32'sd-0.06807728819982777, 32'sd-0.3162397789381797, 32'sd-0.0307019670704824, 32'sd0.3016669702972453, 32'sd0.2963413068196609, 32'sd-0.12575272638711132, 32'sd0.17251172525815286, 32'sd0.3763321069662733, 32'sd0.29038709650414746, 32'sd-0.08615926486835848, 32'sd0.10271196291140149, 32'sd-0.23835209102829608, 32'sd-0.22903718772431353, 32'sd-0.2735400309412271, 32'sd-0.2559005562831855, 32'sd0.02835245027623363, 32'sd0.24160910489187495, 32'sd-0.4235802012809427, 32'sd-0.26616066369808283, 32'sd-0.1882408814501285, 32'sd0.01572970784742376, 32'sd-0.1769978766148591, 32'sd-0.17840440888257963, 32'sd0.21529260460185876, 32'sd0.05291698535975401, 32'sd0.017946712692500193, 32'sd-0.12529749499532894, 32'sd0.1107675219950651},
        '{32'sd0.21023152700043557, 32'sd-0.03706268276813249, 32'sd-0.04484932904388398, 32'sd-0.39478009840940853, 32'sd0.35878454155042383, 32'sd-0.42631210889492516, 32'sd0.20609488528736997, 32'sd-0.41498284398868646, 32'sd0.28406448040165205, 32'sd0.31922001360301905, 32'sd-0.45513150437497296, 32'sd-0.2274397196423357, 32'sd0.35583355722577104, 32'sd0.11601860218868704, 32'sd0.11325226605573253, 32'sd-0.3440559155683922, 32'sd-0.2335769317141076, 32'sd-0.17989062120674662, 32'sd0.3181136251191669, 32'sd0.17981277979657093, 32'sd0.19660579431028186, 32'sd0.23925272869478761, 32'sd0.22077160378459176, 32'sd-0.44465239499768505, 32'sd-0.2905346030084494, 32'sd-0.13885118544748154, 32'sd0.035990227787062304, 32'sd-0.17096898451398698, 32'sd-0.08962281447563412, 32'sd-0.3326508952202071, 32'sd0.2032656349447625, 32'sd-0.4711353572904379, 32'sd-0.3605269091141561, 32'sd0.231407892296884, 32'sd0.06121663521530802, 32'sd-0.11429235177198986, 32'sd-0.17240773783828867, 32'sd0.05560098241057317, 32'sd0.27517078818948415, 32'sd0.013724946524734194, 32'sd0.2055129910333719, 32'sd0.3317953378021122, 32'sd0.16187226745126104, 32'sd-0.4767105044842239, 32'sd-0.036799749572820596, 32'sd-0.05728754537042738, 32'sd-0.2265463820380551, 32'sd0.34126067269008514, 32'sd0.04625572911346797, 32'sd0.191156282578504, 32'sd-0.22087666879254803, 32'sd-0.03932112635132785, 32'sd-0.10877547614480675, 32'sd0.18578763779530083, 32'sd-0.15739532653219376, 32'sd0.01648780127977026, 32'sd0.15937035868941082, 32'sd-0.10792610847974801, 32'sd-0.44710605266567705, 32'sd0.06550962730204313, 32'sd-0.0964930524099936, 32'sd-0.13377506286988305, 32'sd0.45402485403464965, 32'sd-0.31662180963558256},
        '{32'sd-0.09020235669269824, 32'sd-0.3706669389075602, 32'sd-0.46755335792367897, 32'sd0.29654037330212596, 32'sd0.226816244350971, 32'sd0.14230039140293507, 32'sd0.20623418932715587, 32'sd-0.093966901716003, 32'sd0.274764212912734, 32'sd-0.47617355540012685, 32'sd0.2407547125998175, 32'sd-0.3074792445361122, 32'sd0.29150149714191337, 32'sd0.21137403163848797, 32'sd0.25066016661735263, 32'sd-0.20390940785382916, 32'sd0.07579005997957555, 32'sd-0.07173888190406945, 32'sd-0.27987329258770827, 32'sd-0.18403260758155277, 32'sd-0.029053074988141896, 32'sd-0.13463769879280627, 32'sd-0.006332149024367528, 32'sd-0.3283531370379059, 32'sd-0.22105938058756797, 32'sd0.3642481189459236, 32'sd0.27417744348394785, 32'sd0.37001164980025664, 32'sd0.21317080088762924, 32'sd-0.24457568046948142, 32'sd0.08388404658358607, 32'sd0.06719195052146534, 32'sd0.05684943530065423, 32'sd0.28231801855935623, 32'sd0.19034178462202006, 32'sd-0.349092972547409, 32'sd0.308689082951335, 32'sd-0.20639350342627155, 32'sd0.2823775325745333, 32'sd0.13293954880908396, 32'sd0.13116769570280948, 32'sd-0.30896911222527446, 32'sd-0.22812605924885562, 32'sd-0.3992589786040839, 32'sd-0.1123972639283223, 32'sd-0.0012063606293848843, 32'sd-0.2399623955848701, 32'sd-0.3382889942910114, 32'sd0.0247459304580708, 32'sd0.3017857817425127, 32'sd-0.15784418235463993, 32'sd-0.1376853705607859, 32'sd-0.10416278329758137, 32'sd-0.04735056917061775, 32'sd0.21516230611311454, 32'sd0.004413864299878936, 32'sd0.030611261111414597, 32'sd-0.3495252664082127, 32'sd-0.044831116372621764, 32'sd-0.28195502319249327, 32'sd0.22695172492407276, 32'sd-0.07722028098113841, 32'sd-0.6281505119488039, 32'sd0.13640267406680773}
    };

    localparam logic signed [31:0] layer2_biases [0:9] = '{
        32'sd0.14905340143780746, 32'sd0.010366529004123087, 32'sd0.09709577964259249, 32'sd-0.25594789921617683, 32'sd-0.16395858763729224, 32'sd-0.0376090973127773, 32'sd-0.264875406613245, 32'sd-0.32752824517211326, 32'sd0.209751363949506, 32'sd-0.20854157121306932
    };


    //Intermediate outputs
    logic signed [31:0] layer0_out [0:127];
    logic signed [31:0] layer1_out [0:63];


    //Instantiate Layers
    //Layer 0
    layer #(
        .NEURONS(128),
        .PREV_LAYER_OUTPUTS(784)
    ) layer0 (
        .data_inputs(data_inputs),
        .weights(layer0_weights),
        .biases(layer0_biases),
        .data_outputs(layer0_out)
    );

    //Layer 1
    layer #(
        .NEURONS(64),
        .PREV_LAYER_OUTPUTS(128)
    ) layer1 (
        .data_inputs(layer0_out),
        .weights(layer1_weights),
        .biases(layer1_biases),
        .data_outputs(layer1_out)
    );

    //Layer 2
    layer #(
        .NEURONS(10),
        .PREV_LAYER_OUTPUTS(64)
    ) layer2 (
        .data_inputs(layer1_out),
        .weights(layer2_weights),
        .biases(layer2_biases),
        .data_outputs(data_outputs)
    );

endmodule
